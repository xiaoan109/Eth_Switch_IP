// removed module with interface ports: DcpFifo
