************************************************************************
* auCdl Netlist:
*
* Library Name:  SMIC_MEMORY
* Top Cell Name: S55NLLGDPH_X512Y8D16_BW
* Version:  V1.3
* View Name:     schematic
* Netlisted on:  Sat May 18 10:43:14 CST 2024
************************************************************************
*.BIPOLAR
*.RESI = 2000
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM


************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    S55NLLGDPH_X512Y8D16_BW_STWL_DEC
* View Name:    schematic
************************************************************************

.SUBCKT S55NLLGDPH_X512Y8D16_BW_STWL_DEC EMCLK STWL VDD VSS
M0 VSS 2 6 VSS N12LL L=6E-08 W=1E-06
M1 4 4 VSS VSS N12LL L=6E-08 W=4E-07
M2 9 8 EMCLK VSS N12LL L=6E-08 W=8E-07
M3 10 9 VSS VSS N12LL L=6E-08 W=3.5E-07
M4 VSS 9 10 VSS N12LL L=6E-08 W=3.5E-07
M5 11 10 VSS VSS N12LL L=6E-08 W=1.5E-06
M6 VSS 10 11 VSS N12LL L=6E-08 W=1.5E-06
M7 STWL 11 VSS VSS N12LL L=6E-08 W=2E-06
M8 VSS 11 STWL VSS N12LL L=6E-08 W=2E-06
M9 STWL 11 VDD VDD PHVT12LL L=6E-08 W=2.5E-06
M10 VDD 11 STWL VDD PHVT12LL L=6E-08 W=2.5E-06
M11 STWL 11 VDD VDD PHVT12LL L=6E-08 W=2.5E-06
M12 VDD 11 STWL VDD PHVT12LL L=6E-08 W=2.5E-06
M13 9 8 VDD VDD P12LL L=6E-08 W=4E-07
M14 8 4 VDD VDD P12LL L=6E-08 W=1E-06
M15 9 6 EMCLK VDD P12LL L=6E-08 W=4E-07
M16 VDD 2 2 VDD P12LL L=6E-08 W=4E-07
M17 10 9 VDD VDD P12LL L=6E-08 W=7E-07
M18 VDD 9 10 VDD P12LL L=6E-08 W=7E-07
M19 11 10 VDD VDD P12LL L=6E-08 W=1.5E-06
M20 VDD 10 11 VDD P12LL L=6E-08 W=1.5E-06
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    S55NLLGDPH_X512Y8D16_BW_BLSTRAP_B
* View Name:    schematic
************************************************************************

.SUBCKT S55NLLGDPH_X512Y8D16_BW_BLSTRAP_B BL BLX VDD VSS
MTA1 BLX VSS NET22 VSS DPNPGBHVT W=100.00N L=85.000N M=1
MTA0 BL VSS NET26 VSS DPNPGAHVT W=100.0N L=85.000N M=1
MTD1 NET31 VSS VSS VSS DPNPDHVT W=310.00N L=70.00N M=1
MTL1 NET33 VSS VDD VDD DPPLHVT W=85.000N L=70.00N M=1
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    S55NLLGDPH_X512Y8D16_BW_EDGECELL
* View Name:    schematic
************************************************************************

.SUBCKT S55NLLGDPH_X512Y8D16_BW_EDGECELL BA BB BXA BXB VDD VSS WLA
MTD0 VSS BCN BC VSS DPNPDHVT W=310.00N L=70.00N M=1
MM2 BCN BC VSS VSS DPNPDHVT W=310.00N L=70.00N M=1
MM1 BCN BC VDD VDD DPPLHVT W=85.000N L=70.00N M=1
MTL0 VDD BCN BC VDD DPPLHVT W=85.000N L=70.00N M=1
MTA1 BXA WLA BCN VSS DPNPGBHVT W=100.00N L=85.000N M=1
MN1 BC VSS BB VSS DPNPGBHVT W=100.00N L=85.000N M=1
MM0 BXB VSS BCN VSS DPNPGAHVT W=100.0N L=85.000N M=1
MTA0 BC WLA BA VSS DPNPGAHVT W=100.0N L=85.000N M=1
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    S55NLLGDPH_X512Y8D16_BW_EDGECELL8B
* View Name:    schematic
************************************************************************

.SUBCKT S55NLLGDPH_X512Y8D16_BW_EDGECELL8B BA0 BA7 BXA0 BXA7 VDD VSS WLA[7] WLA[6] WLA[5] WLA[4]
+WLA[3] WLA[2] WLA[1] WLA[0]
XI22 BA7 NET43 BXA7 NET42 VDD VSS WLA[7] S55NLLGDPH_X512Y8D16_BW_EDGECELL
XI19 NET52 NET85 NET51 NET84 VDD VSS WLA[4] S55NLLGDPH_X512Y8D16_BW_EDGECELL
XI18 NET52 NET57 NET51 NET56 VDD VSS WLA[3] S55NLLGDPH_X512Y8D16_BW_EDGECELL
XI16 NET73 NET64 NET72 NET63 VDD VSS WLA[1] S55NLLGDPH_X512Y8D16_BW_EDGECELL
XI17 NET73 NET57 NET72 NET56 VDD VSS WLA[2] S55NLLGDPH_X512Y8D16_BW_EDGECELL
XI21 NET80 NET43 NET79 NET42 VDD VSS WLA[6] S55NLLGDPH_X512Y8D16_BW_EDGECELL
XI20 NET80 NET85 NET79 NET84 VDD VSS WLA[5] S55NLLGDPH_X512Y8D16_BW_EDGECELL
XI15 BA0 NET64 BXA0 NET63 VDD VSS WLA[0] S55NLLGDPH_X512Y8D16_BW_EDGECELL
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    S55NLLGDPH_X512Y8D16_BW_EDGECELL66B_RED_LEFT
* View Name:    schematic
************************************************************************

.SUBCKT S55NLLGDPH_X512Y8D16_BW_EDGECELL66B_RED_LEFT RWL[0] RWL[1] VDD VSS WLA[63] WLA[62] WLA[61] WLA[60] WLA[59] WLA[58]
+WLA[57] WLA[56] WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48]
+WLA[47] WLA[46] WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38]
+WLA[37] WLA[36] WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28]
+WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18]
+WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8]
+WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0]
XI0 NET01 NET61 VDD VSS S55NLLGDPH_X512Y8D16_BW_BLSTRAP_B
XI1 NET01 NET31 NET61 NET91 VDD VSS RWL[0] S55NLLGDPH_X512Y8D16_BW_EDGECELL
XI2 NET02 NET31 NET62 NET91 VDD VSS RWL[1] S55NLLGDPH_X512Y8D16_BW_EDGECELL
XI3 NET02 NET32 NET62 NET92 VDD VSS WLA[7] WLA[6] WLA[5] WLA[4]
+WLA[3] WLA[2] WLA[1] WLA[0] S55NLLGDPH_X512Y8D16_BW_EDGECELL8B
XI4 NET03 NET32 NET63 NET92 VDD VSS WLA[15] WLA[14] WLA[13] WLA[12]
+WLA[11] WLA[10] WLA[9] WLA[8] S55NLLGDPH_X512Y8D16_BW_EDGECELL8B
XI5 NET03 NET33 NET63 NET93 VDD VSS WLA[23] WLA[22] WLA[21] WLA[20]
+WLA[19] WLA[18] WLA[17] WLA[16] S55NLLGDPH_X512Y8D16_BW_EDGECELL8B
XI6 NET04 NET33 NET64 NET93 VDD VSS WLA[31] WLA[30] WLA[29] WLA[28]
+WLA[27] WLA[26] WLA[25] WLA[24] S55NLLGDPH_X512Y8D16_BW_EDGECELL8B
XI7 NET04 NET34 NET64 NET94 VDD VSS WLA[39] WLA[38] WLA[37] WLA[36]
+WLA[35] WLA[34] WLA[33] WLA[32] S55NLLGDPH_X512Y8D16_BW_EDGECELL8B
XI8 NET05 NET34 NET65 NET94 VDD VSS WLA[47] WLA[46] WLA[45] WLA[44]
+WLA[43] WLA[42] WLA[41] WLA[40] S55NLLGDPH_X512Y8D16_BW_EDGECELL8B
XI9 NET05 NET35 NET65 NET95 VDD VSS WLA[55] WLA[54] WLA[53] WLA[52]
+WLA[51] WLA[50] WLA[49] WLA[48] S55NLLGDPH_X512Y8D16_BW_EDGECELL8B
XI10 NET06 NET35 NET66 NET95 VDD VSS WLA[63] WLA[62] WLA[61] WLA[60]
+WLA[59] WLA[58] WLA[57] WLA[56] S55NLLGDPH_X512Y8D16_BW_EDGECELL8B
XI11 NET06 NET66 VDD VSS S55NLLGDPH_X512Y8D16_BW_BLSTRAP_B
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    S55NLLGDPH_X512Y8D16_BW_BLSTRAP
* View Name:    schematic
************************************************************************

.SUBCKT S55NLLGDPH_X512Y8D16_BW_BLSTRAP BL BLX VDD VSS
MTA1 BL VSS NET22 VSS DPNPGBHVT W=100.00N L=85.000N M=1
MTA0 BLX VSS NET26 VSS DPNPGAHVT W=100.0N L=85.000N M=1
MTD1 NET31 VSS VSS VSS DPNPDHVT W=310.00N L=70.00N M=1
MTL1 NET33 VSS VDD VDD DPPLHVT W=85.000N L=70.00N M=1
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    S55NLLGDPH_X512Y8D16_BW_EDGECELL8A
* View Name:    schematic
************************************************************************

.SUBCKT S55NLLGDPH_X512Y8D16_BW_EDGECELL8A BB0 BB7 BXB0 BXB7 VDD VSS WLA[7] WLA[6] WLA[5] WLA[4]
+WLA[3] WLA[2] WLA[1] WLA[0]
XI19 NET52 NET43 NET51 NET42 VDD VSS WLA[4] S55NLLGDPH_X512Y8D16_BW_EDGECELL
XI20 NET52 NET64 NET51 NET63 VDD VSS WLA[5] S55NLLGDPH_X512Y8D16_BW_EDGECELL
XI22 NET59 BB7 NET58 BXB7 VDD VSS WLA[7] S55NLLGDPH_X512Y8D16_BW_EDGECELL
XI21 NET59 NET64 NET58 NET63 VDD VSS WLA[6] S55NLLGDPH_X512Y8D16_BW_EDGECELL
XI17 NET80 NET71 NET79 NET70 VDD VSS WLA[2] S55NLLGDPH_X512Y8D16_BW_EDGECELL
XI18 NET80 NET43 NET79 NET42 VDD VSS WLA[3] S55NLLGDPH_X512Y8D16_BW_EDGECELL
XI16 NET87 NET71 NET86 NET70 VDD VSS WLA[1] S55NLLGDPH_X512Y8D16_BW_EDGECELL
XI15 NET87 BB0 NET86 BXB0 VDD VSS WLA[0] S55NLLGDPH_X512Y8D16_BW_EDGECELL
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    S55NLLGDPH_X512Y8D16_BW_EDGECELL64A_LEFT
* View Name:    schematic
************************************************************************

.SUBCKT S55NLLGDPH_X512Y8D16_BW_EDGECELL64A_LEFT VDD VSS WLA[63] WLA[62] WLA[61] WLA[60] WLA[59] WLA[58] WLA[57] WLA[56]
+WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48] WLA[47] WLA[46]
+WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38] WLA[37] WLA[36]
+WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28] WLA[27] WLA[26]
+WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18] WLA[17] WLA[16]
+WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8] WLA[7] WLA[6]
+WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0]
XI0 NET01 NET61 VDD VSS S55NLLGDPH_X512Y8D16_BW_BLSTRAP
XI1 NET01 NET31 NET61 NET91 VDD VSS WLA[7] WLA[6] WLA[5] WLA[4]
+WLA[3] WLA[2] WLA[1] WLA[0] S55NLLGDPH_X512Y8D16_BW_EDGECELL8A
XI2 NET02 NET31 NET62 NET91 VDD VSS WLA[15] WLA[14] WLA[13] WLA[12]
+WLA[11] WLA[10] WLA[9] WLA[8] S55NLLGDPH_X512Y8D16_BW_EDGECELL8A
XI3 NET02 NET32 NET62 NET92 VDD VSS WLA[23] WLA[22] WLA[21] WLA[20]
+WLA[19] WLA[18] WLA[17] WLA[16] S55NLLGDPH_X512Y8D16_BW_EDGECELL8A
XI4 NET03 NET32 NET63 NET92 VDD VSS WLA[31] WLA[30] WLA[29] WLA[28]
+WLA[27] WLA[26] WLA[25] WLA[24] S55NLLGDPH_X512Y8D16_BW_EDGECELL8A
XI5 NET03 NET33 NET63 NET93 VDD VSS WLA[39] WLA[38] WLA[37] WLA[36]
+WLA[35] WLA[34] WLA[33] WLA[32] S55NLLGDPH_X512Y8D16_BW_EDGECELL8A
XI6 NET04 NET33 NET64 NET93 VDD VSS WLA[47] WLA[46] WLA[45] WLA[44]
+WLA[43] WLA[42] WLA[41] WLA[40] S55NLLGDPH_X512Y8D16_BW_EDGECELL8A
XI7 NET04 NET34 NET64 NET94 VDD VSS WLA[55] WLA[54] WLA[53] WLA[52]
+WLA[51] WLA[50] WLA[49] WLA[48] S55NLLGDPH_X512Y8D16_BW_EDGECELL8A
XI8 NET05 NET34 NET65 NET94 VDD VSS WLA[63] WLA[62] WLA[61] WLA[60]
+WLA[59] WLA[58] WLA[57] WLA[56] S55NLLGDPH_X512Y8D16_BW_EDGECELL8A
XI9 NET05 NET65 VDD VSS S55NLLGDPH_X512Y8D16_BW_BLSTRAP
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    S55NLLGDPH_X512Y8D16_BW_EDGECELL64B_LEFT
* View Name:    schematic
************************************************************************

.SUBCKT S55NLLGDPH_X512Y8D16_BW_EDGECELL64B_LEFT VDD VSS WLA[63] WLA[62] WLA[61] WLA[60] WLA[59] WLA[58] WLA[57] WLA[56]
+WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48] WLA[47] WLA[46]
+WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38] WLA[37] WLA[36]
+WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28] WLA[27] WLA[26]
+WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18] WLA[17] WLA[16]
+WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8] WLA[7] WLA[6]
+WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0]
XI0 NET01 NET61 VDD VSS S55NLLGDPH_X512Y8D16_BW_BLSTRAP_B
XI1 NET01 NET31 NET61 NET91 VDD VSS WLA[7] WLA[6] WLA[5] WLA[4]
+WLA[3] WLA[2] WLA[1] WLA[0] S55NLLGDPH_X512Y8D16_BW_EDGECELL8B
XI2 NET02 NET31 NET62 NET91 VDD VSS WLA[15] WLA[14] WLA[13] WLA[12]
+WLA[11] WLA[10] WLA[9] WLA[8] S55NLLGDPH_X512Y8D16_BW_EDGECELL8B
XI3 NET02 NET32 NET62 NET92 VDD VSS WLA[23] WLA[22] WLA[21] WLA[20]
+WLA[19] WLA[18] WLA[17] WLA[16] S55NLLGDPH_X512Y8D16_BW_EDGECELL8B
XI4 NET03 NET32 NET63 NET92 VDD VSS WLA[31] WLA[30] WLA[29] WLA[28]
+WLA[27] WLA[26] WLA[25] WLA[24] S55NLLGDPH_X512Y8D16_BW_EDGECELL8B
XI5 NET03 NET33 NET63 NET93 VDD VSS WLA[39] WLA[38] WLA[37] WLA[36]
+WLA[35] WLA[34] WLA[33] WLA[32] S55NLLGDPH_X512Y8D16_BW_EDGECELL8B
XI6 NET04 NET33 NET64 NET93 VDD VSS WLA[47] WLA[46] WLA[45] WLA[44]
+WLA[43] WLA[42] WLA[41] WLA[40] S55NLLGDPH_X512Y8D16_BW_EDGECELL8B
XI7 NET04 NET34 NET64 NET94 VDD VSS WLA[55] WLA[54] WLA[53] WLA[52]
+WLA[51] WLA[50] WLA[49] WLA[48] S55NLLGDPH_X512Y8D16_BW_EDGECELL8B
XI8 NET05 NET34 NET65 NET94 VDD VSS WLA[63] WLA[62] WLA[61] WLA[60]
+WLA[59] WLA[58] WLA[57] WLA[56] S55NLLGDPH_X512Y8D16_BW_EDGECELL8B
XI9 NET05 NET65 VDD VSS S55NLLGDPH_X512Y8D16_BW_BLSTRAP_B
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    S55NLLGDPH_X512Y8D16_BW_EDGECELL4A
* View Name:    schematic
************************************************************************

.SUBCKT S55NLLGDPH_X512Y8D16_BW_EDGECELL4A BB0 BB3 BXB0 BXB3 VDD VSS WLA[3] WLA[2] WLA[1] WLA[0]
XI22 NET80 BB3 NET58 BXB3 VDD VSS WLA[3] S55NLLGDPH_X512Y8D16_BW_EDGECELL
XI17 NET80 NET71 NET58 NET70 VDD VSS WLA[2] S55NLLGDPH_X512Y8D16_BW_EDGECELL
XI16 NET87 NET71 NET86 NET70 VDD VSS WLA[1] S55NLLGDPH_X512Y8D16_BW_EDGECELL
XI15 NET87 BB0 NET86 BXB0 VDD VSS WLA[0] S55NLLGDPH_X512Y8D16_BW_EDGECELL
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    S55NLLGDPH_X512Y8D16_BW_EDGECELL68A_TOP_LEFT
* View Name:    schematic
************************************************************************

.SUBCKT S55NLLGDPH_X512Y8D16_BW_EDGECELL68A_TOP_LEFT VDD VSS WLA[63] WLA[62] WLA[61] WLA[60] WLA[59] WLA[58] WLA[57] WLA[56]
+WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48] WLA[47] WLA[46]
+WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38] WLA[37] WLA[36]
+WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28] WLA[27] WLA[26]
+WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18] WLA[17] WLA[16]
+WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8] WLA[7] WLA[6]
+WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0]
XI0 NET01 NET61 VDD VSS S55NLLGDPH_X512Y8D16_BW_BLSTRAP
XI1 NET01 NET31 NET61 NET91 VDD VSS WLA[7] WLA[6] WLA[5] WLA[4]
+WLA[3] WLA[2] WLA[1] WLA[0] S55NLLGDPH_X512Y8D16_BW_EDGECELL8A
XI2 NET02 NET31 NET62 NET91 VDD VSS WLA[15] WLA[14] WLA[13] WLA[12]
+WLA[11] WLA[10] WLA[9] WLA[8] S55NLLGDPH_X512Y8D16_BW_EDGECELL8A
XI3 NET02 NET32 NET62 NET92 VDD VSS WLA[23] WLA[22] WLA[21] WLA[20]
+WLA[19] WLA[18] WLA[17] WLA[16] S55NLLGDPH_X512Y8D16_BW_EDGECELL8A
XI4 NET03 NET32 NET63 NET92 VDD VSS WLA[31] WLA[30] WLA[29] WLA[28]
+WLA[27] WLA[26] WLA[25] WLA[24] S55NLLGDPH_X512Y8D16_BW_EDGECELL8A
XI5 NET03 NET33 NET63 NET93 VDD VSS WLA[39] WLA[38] WLA[37] WLA[36]
+WLA[35] WLA[34] WLA[33] WLA[32] S55NLLGDPH_X512Y8D16_BW_EDGECELL8A
XI6 NET04 NET33 NET64 NET93 VDD VSS WLA[47] WLA[46] WLA[45] WLA[44]
+WLA[43] WLA[42] WLA[41] WLA[40] S55NLLGDPH_X512Y8D16_BW_EDGECELL8A
XI7 NET04 NET34 NET64 NET94 VDD VSS WLA[55] WLA[54] WLA[53] WLA[52]
+WLA[51] WLA[50] WLA[49] WLA[48] S55NLLGDPH_X512Y8D16_BW_EDGECELL8A
XI8 NET05 NET34 NET65 NET94 VDD VSS WLA[63] WLA[62] WLA[61] WLA[60]
+WLA[59] WLA[58] WLA[57] WLA[56] S55NLLGDPH_X512Y8D16_BW_EDGECELL8A
XI9 NET05 NET35 NET65 NET95 VDD VSS VSS VSS VSS VSS S55NLLGDPH_X512Y8D16_BW_EDGECELL4A
XI10 NET35 NET95 VDD VSS S55NLLGDPH_X512Y8D16_BW_BLSTRAP
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    S55NLLGDPH_X512Y8D16_BW_BITCELL_ST
* View Name:    schematic
************************************************************************

.SUBCKT S55NLLGDPH_X512Y8D16_BW_BITCELL_ST BA BB BXA BXB VDD VSS WLA
MTD0 VSS BCN BC VSS DPNPDHVT W=310.00N L=70.00N M=1
MM2 BCN BC VSS VSS DPNPDHVT W=310.00N L=70.00N M=1
MM1 BCN BC VDD VDD DPPLHVT W=85.000N L=70.00N M=1
MTL0 VDD BCN BC VDD DPPLHVT W=85.000N L=70.00N M=1
MTA1 BXA WLA BCN VSS DPNPGBHVT W=100.00N L=85.000N M=1
MN1 BC VSS BB VSS DPNPGBHVT W=100.00N L=85.000N M=1
MM0 BXB VSS BCN VSS DPNPGAHVT W=100.0N L=85.000N M=1
MTA0 BC WLA BA VSS DPNPGAHVT W=100.0N L=85.000N M=1
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    S55NLLGDPH_X512Y8D16_BW_BITCELL_ST8B
* View Name:    schematic
************************************************************************

.SUBCKT S55NLLGDPH_X512Y8D16_BW_BITCELL_ST8B BA0 BA7 BXA0 BXA7 DUM_BL VDD VSS WLA[7] WLA[6] WLA[5]
+WLA[4] WLA[3] WLA[2] WLA[1] WLA[0]
XI0 NET47 DUM_BL NET46 NET51 VDD VSS WLA[6] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST
XI1 BA7 DUM_BL BXA7 NET51 VDD VSS WLA[7] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST
XI2 NET47 DUM_BL NET46 NET58 VDD VSS WLA[5] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST
XI3 NET68 DUM_BL NET67 NET58 VDD VSS WLA[4] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST
XI4 NET68 DUM_BL NET67 NET72 VDD VSS WLA[3] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST
XI5 NET82 DUM_BL NET81 NET72 VDD VSS WLA[2] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST
XI6 NET82 DUM_BL NET81 NET86 VDD VSS WLA[1] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST
XI7 BA0 DUM_BL BXA0 NET86 VDD VSS WLA[0] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    S55NLLGDPH_X512Y8D16_BW_BITCELL_ST66B
* View Name:    schematic
************************************************************************

.SUBCKT S55NLLGDPH_X512Y8D16_BW_BITCELL_ST66B DUM_BL RWL[0] RWL[1] VDD VSS WLA[63] WLA[62] WLA[61] WLA[60] WLA[59]
+WLA[58] WLA[57] WLA[56] WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50] WLA[49]
+WLA[48] WLA[47] WLA[46] WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39]
+WLA[38] WLA[37] WLA[36] WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29]
+WLA[28] WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19]
+WLA[18] WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9]
+WLA[8] WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0]
XI0 NET01 NET61 VDD VSS S55NLLGDPH_X512Y8D16_BW_BLSTRAP_B
XI1 NET01 DUM_BL NET61 NET91 VDD VSS RWL[0] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST
XI2 NET02 DUM_BL NET62 NET91 VDD VSS RWL[1] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST
XI3 NET02 NET31 NET62 NET92 DUM_BL VDD VSS WLA[7] WLA[6] WLA[5]
+WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST8B
XI4 NET03 NET31 NET63 NET92 DUM_BL VDD VSS WLA[15] WLA[14] WLA[13]
+WLA[12] WLA[11] WLA[10] WLA[9] WLA[8] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST8B
XI5 NET03 NET32 NET63 NET93 DUM_BL VDD VSS WLA[23] WLA[22] WLA[21]
+WLA[20] WLA[19] WLA[18] WLA[17] WLA[16] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST8B
XI6 NET04 NET32 NET64 NET93 DUM_BL VDD VSS WLA[31] WLA[30] WLA[29]
+WLA[28] WLA[27] WLA[26] WLA[25] WLA[24] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST8B
XI7 NET04 NET33 NET64 NET94 DUM_BL VDD VSS WLA[39] WLA[38] WLA[37]
+WLA[36] WLA[35] WLA[34] WLA[33] WLA[32] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST8B
XI8 NET05 NET33 NET65 NET94 DUM_BL VDD VSS WLA[47] WLA[46] WLA[45]
+WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST8B
XI9 NET05 NET34 NET65 NET95 DUM_BL VDD VSS WLA[55] WLA[54] WLA[53]
+WLA[52] WLA[51] WLA[50] WLA[49] WLA[48] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST8B
XI10 NET06 NET34 NET66 NET95 DUM_BL VDD VSS WLA[63] WLA[62] WLA[61]
+WLA[60] WLA[59] WLA[58] WLA[57] WLA[56] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST8B
XI11 NET06 NET66 VDD VSS S55NLLGDPH_X512Y8D16_BW_BLSTRAP_B
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    S55NLLGDPH_X512Y8D16_BW_BITCELL_ST8A
* View Name:    schematic
************************************************************************

.SUBCKT S55NLLGDPH_X512Y8D16_BW_BITCELL_ST8A BXB0 BXB7 DUMBL VDD VSS WLA[7] WLA[6] WLA[5] WLA[4] WLA[3]
+WLA[2] WLA[1] WLA[0]
XI0 NET52 DUMBL NET51 BXB7 VDD VSS WLA[7] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST
XI1 NET52 DUMBL NET51 NET42 VDD VSS WLA[6] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST
XI2 NET59 DUMBL NET58 NET42 VDD VSS WLA[5] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST
XI3 NET59 DUMBL NET58 NET63 VDD VSS WLA[4] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST
XI4 NET73 DUMBL NET72 NET63 VDD VSS WLA[3] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST
XI5 NET73 DUMBL NET72 NET77 VDD VSS WLA[2] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST
XI6 NET87 DUMBL NET86 NET77 VDD VSS WLA[1] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST
XI7 NET87 DUMBL NET86 BXB0 VDD VSS WLA[0] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    S55NLLGDPH_X512Y8D16_BW_BITCELL_ST64A
* View Name:    schematic
************************************************************************

.SUBCKT S55NLLGDPH_X512Y8D16_BW_BITCELL_ST64A DUM_BL VDD VSS WLA[63] WLA[62] WLA[61] WLA[60] WLA[59] WLA[58] WLA[57]
+WLA[56] WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48] WLA[47]
+WLA[46] WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38] WLA[37]
+WLA[36] WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28] WLA[27]
+WLA[26] WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18] WLA[17]
+WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8] WLA[7]
+WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0]
XI0 DUM_BL NET025 VDD VSS S55NLLGDPH_X512Y8D16_BW_BLSTRAP
XI1 DUM_BL NET50 VDD VSS S55NLLGDPH_X512Y8D16_BW_BLSTRAP
XI2 NET32 NET37 DUM_BL VDD VSS WLA[23] WLA[22] WLA[21] WLA[20] WLA[19]
+WLA[18] WLA[17] WLA[16] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST8A
XI3 NET25 NET37 DUM_BL VDD VSS WLA[31] WLA[30] WLA[29] WLA[28] WLA[27]
+WLA[26] WLA[25] WLA[24] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST8A
XI4 NET051 NET044 DUM_BL VDD VSS WLA[55] WLA[54] WLA[53] WLA[52] WLA[51]
+WLA[50] WLA[49] WLA[48] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST8A
XI5 NET025 NET044 DUM_BL VDD VSS WLA[63] WLA[62] WLA[61] WLA[60] WLA[59]
+WLA[58] WLA[57] WLA[56] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST8A
XI6 NET051 NET038 DUM_BL VDD VSS WLA[47] WLA[46] WLA[45] WLA[44] WLA[43]
+WLA[42] WLA[41] WLA[40] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST8A
XI7 NET25 NET038 DUM_BL VDD VSS WLA[39] WLA[38] WLA[37] WLA[36] WLA[35]
+WLA[34] WLA[33] WLA[32] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST8A
XI8 NET32 NET43 DUM_BL VDD VSS WLA[15] WLA[14] WLA[13] WLA[12] WLA[11]
+WLA[10] WLA[9] WLA[8] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST8A
XI9 NET50 NET43 DUM_BL VDD VSS WLA[7] WLA[6] WLA[5] WLA[4] WLA[3]
+WLA[2] WLA[1] WLA[0] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST8A
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    S55NLLGDPH_X512Y8D16_BW_BITCELL_ST64B
* View Name:    schematic
************************************************************************

.SUBCKT S55NLLGDPH_X512Y8D16_BW_BITCELL_ST64B DUM_BL VDD VSS WLA[63] WLA[62] WLA[61] WLA[60] WLA[59] WLA[58] WLA[57]
+WLA[56] WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48] WLA[47]
+WLA[46] WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38] WLA[37]
+WLA[36] WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28] WLA[27]
+WLA[26] WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18] WLA[17]
+WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8] WLA[7]
+WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0]
XI0 NET69 NET66 VDD VSS S55NLLGDPH_X512Y8D16_BW_BLSTRAP_B
XI1 NET36 NET35 VDD VSS S55NLLGDPH_X512Y8D16_BW_BLSTRAP_B
XI2 NET059 NET049 NET056 NET052 DUM_BL VDD VSS WLA[55] WLA[54] WLA[53]
+WLA[52] WLA[51] WLA[50] WLA[49] WLA[48] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST8B
XI3 NET69 NET049 NET66 NET052 DUM_BL VDD VSS WLA[63] WLA[62] WLA[61]
+WLA[60] WLA[59] WLA[58] WLA[57] WLA[56] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST8B
XI4 NET36 NET41 NET35 NET44 DUM_BL VDD VSS WLA[7] WLA[6] WLA[5]
+WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST8B
XI5 NET51 NET41 NET48 NET44 DUM_BL VDD VSS WLA[15] WLA[14] WLA[13]
+WLA[12] WLA[11] WLA[10] WLA[9] WLA[8] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST8B
XI6 NET51 NET57 NET48 NET60 DUM_BL VDD VSS WLA[23] WLA[22] WLA[21]
+WLA[20] WLA[19] WLA[18] WLA[17] WLA[16] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST8B
XI7 NET0101 NET57 NET098 NET60 DUM_BL VDD VSS WLA[31] WLA[30] WLA[29]
+WLA[28] WLA[27] WLA[26] WLA[25] WLA[24] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST8B
XI8 NET059 NET065 NET056 NET068 DUM_BL VDD VSS WLA[47] WLA[46] WLA[45]
+WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST8B
XI9 NET0101 NET065 NET098 NET068 DUM_BL VDD VSS WLA[39] WLA[38] WLA[37]
+WLA[36] WLA[35] WLA[34] WLA[33] WLA[32] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST8B
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    S55NLLGDPH_X512Y8D16_BW_BITCELL_ST8B_TW
* View Name:    schematic
************************************************************************

.SUBCKT S55NLLGDPH_X512Y8D16_BW_BITCELL_ST8B_TW BA0 BA7 BXA0 BXA7 DUM_BL VDD VSS WLA[7] WLA[6] WLA[5]
+WLA[4] WLA[3] WLA[2] WLA[1] WLA[0]
XI0 BA7 NET45 BXA7 DUM_BL VDD VSS WLA[7] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST
XI1 NET54 NET45 NET53 DUM_BL VDD VSS WLA[6] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST
XI2 NET54 NET59 NET53 DUM_BL VDD VSS WLA[5] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST
XI3 NET68 NET59 NET67 DUM_BL VDD VSS WLA[4] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST
XI4 NET68 NET73 NET67 DUM_BL VDD VSS WLA[3] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST
XI5 NET82 NET73 NET81 DUM_BL VDD VSS WLA[2] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST
XI6 NET82 NET87 NET81 DUM_BL VDD VSS WLA[1] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST
XI7 BA0 NET87 BXA0 DUM_BL VDD VSS WLA[0] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    S55NLLGDPH_X512Y8D16_BW_BITCELL_ST64B_TW_LEFT
* View Name:    schematic
************************************************************************

.SUBCKT S55NLLGDPH_X512Y8D16_BW_BITCELL_ST64B_TW_LEFT DUM_BL VDD VSS WLA[63] WLA[62] WLA[61] WLA[60] WLA[59] WLA[58] WLA[57]
+WLA[56] WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48] WLA[47]
+WLA[46] WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38] WLA[37]
+WLA[36] WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28] WLA[27]
+WLA[26] WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18] WLA[17]
+WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8] WLA[7]
+WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0]
XI0 NET01 NET61 VDD VSS S55NLLGDPH_X512Y8D16_BW_BLSTRAP_B
XI1 NET01 NET31 NET61 NET91 DUM_BL VDD VSS WLA[7] WLA[6] WLA[5]
+WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST8B_TW
XI2 NET02 NET31 NET62 NET91 DUM_BL VDD VSS WLA[15] WLA[14] WLA[13]
+WLA[12] WLA[11] WLA[10] WLA[9] WLA[8] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST8B_TW
XI3 NET02 NET32 NET62 NET92 DUM_BL VDD VSS WLA[23] WLA[22] WLA[21]
+WLA[20] WLA[19] WLA[18] WLA[17] WLA[16] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST8B_TW
XI4 NET03 NET32 NET63 NET92 DUM_BL VDD VSS WLA[31] WLA[30] WLA[29]
+WLA[28] WLA[27] WLA[26] WLA[25] WLA[24] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST8B_TW
XI5 NET03 NET33 NET63 NET93 DUM_BL VDD VSS WLA[39] WLA[38] WLA[37]
+WLA[36] WLA[35] WLA[34] WLA[33] WLA[32] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST8B_TW
XI6 NET04 NET33 NET64 NET93 DUM_BL VDD VSS WLA[47] WLA[46] WLA[45]
+WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST8B_TW
XI7 NET04 NET34 NET64 NET94 DUM_BL VDD VSS WLA[55] WLA[54] WLA[53]
+WLA[52] WLA[51] WLA[50] WLA[49] WLA[48] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST8B_TW
XI8 NET05 NET34 NET65 NET94 DUM_BL VDD VSS WLA[63] WLA[62] WLA[61]
+WLA[60] WLA[59] WLA[58] WLA[57] WLA[56] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST8B_TW
XI9 NET05 NET65 VDD VSS S55NLLGDPH_X512Y8D16_BW_BLSTRAP_B
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    S55NLLGDPH_X512Y8D16_BW_BITCELL_ST8A_TW
* View Name:    schematic
************************************************************************

.SUBCKT S55NLLGDPH_X512Y8D16_BW_BITCELL_ST8A_TW BB0 BB7 DUMBL VDD VSS WLA[7] WLA[6] WLA[5] WLA[4] WLA[3]
+WLA[2] WLA[1] WLA[0]
XI0 NET52 NET43 NET51 DUMBL VDD VSS WLA[6] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST
XI1 NET52 BB7 NET51 DUMBL VDD VSS WLA[7] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST
XI2 NET59 NET43 NET58 DUMBL VDD VSS WLA[5] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST
XI3 NET59 NET64 NET58 DUMBL VDD VSS WLA[4] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST
XI4 NET73 NET64 NET72 DUMBL VDD VSS WLA[3] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST
XI5 NET73 NET78 NET72 DUMBL VDD VSS WLA[2] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST
XI6 NET87 NET78 NET86 DUMBL VDD VSS WLA[1] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST
XI7 NET87 BB0 NET86 DUMBL VDD VSS WLA[0] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    S55NLLGDPH_X512Y8D16_BW_BITCELL_ST64A_TW_LEFT
* View Name:    schematic
************************************************************************

.SUBCKT S55NLLGDPH_X512Y8D16_BW_BITCELL_ST64A_TW_LEFT DUM_BL VDD VSS WLA[63] WLA[62] WLA[61] WLA[60] WLA[59] WLA[58] WLA[57]
+WLA[56] WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48] WLA[47]
+WLA[46] WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38] WLA[37]
+WLA[36] WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28] WLA[27]
+WLA[26] WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18] WLA[17]
+WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8] WLA[7]
+WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0]
XI0 NET01 DUM_BL VDD VSS S55NLLGDPH_X512Y8D16_BW_BLSTRAP
XI1 NET01 NET31 DUM_BL VDD VSS WLA[7] WLA[6] WLA[5] WLA[4] WLA[3]
+WLA[2] WLA[1] WLA[0] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST8A_TW
XI2 NET02 NET31 DUM_BL VDD VSS WLA[15] WLA[14] WLA[13] WLA[12] WLA[11]
+WLA[10] WLA[9] WLA[8] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST8A_TW
XI3 NET02 NET32 DUM_BL VDD VSS WLA[23] WLA[22] WLA[21] WLA[20] WLA[19]
+WLA[18] WLA[17] WLA[16] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST8A_TW
XI4 NET03 NET32 DUM_BL VDD VSS WLA[31] WLA[30] WLA[29] WLA[28] WLA[27]
+WLA[26] WLA[25] WLA[24] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST8A_TW
XI5 NET03 NET33 DUM_BL VDD VSS WLA[39] WLA[38] WLA[37] WLA[36] WLA[35]
+WLA[34] WLA[33] WLA[32] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST8A_TW
XI6 NET04 NET33 DUM_BL VDD VSS WLA[47] WLA[46] WLA[45] WLA[44] WLA[43]
+WLA[42] WLA[41] WLA[40] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST8A_TW
XI7 NET04 NET34 DUM_BL VDD VSS WLA[55] WLA[54] WLA[53] WLA[52] WLA[51]
+WLA[50] WLA[49] WLA[48] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST8A_TW
XI8 NET05 NET34 DUM_BL VDD VSS WLA[63] WLA[62] WLA[61] WLA[60] WLA[59]
+WLA[58] WLA[57] WLA[56] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST8A_TW
XI9 NET05 DUM_BL VDD VSS S55NLLGDPH_X512Y8D16_BW_BLSTRAP
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    S55NLLGDPH_X512Y8D16_BW_BITCELL_ST4A_TW
* View Name:    schematic
************************************************************************

.SUBCKT S55NLLGDPH_X512Y8D16_BW_BITCELL_ST4A_TW BB0 BB3 BBX0 BBX3 VDD VSS WLA[3] WLA[2] WLA[1] WLA[0]
XI22 NET46 BB3 NET45 BBX3 VDD VSS WLA[3] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST
XI21 NET46 NET51 NET45 NET041 VDD VSS WLA[2] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST
XI20 NET60 NET51 NET59 NET041 VDD VSS WLA[1] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST
XI0 NET60 BB0 NET59 BBX0 VDD VSS WLA[0] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    S55NLLGDPH_X512Y8D16_BW_BITCELL_ST68A_TOP_TW_LEFT
* View Name:    schematic
************************************************************************

.SUBCKT S55NLLGDPH_X512Y8D16_BW_BITCELL_ST68A_TOP_TW_LEFT DUM_BL STWLA VDD VSS WLA[63] WLA[62] WLA[61] WLA[60] WLA[59] WLA[58]
+WLA[57] WLA[56] WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48]
+WLA[47] WLA[46] WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38]
+WLA[37] WLA[36] WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28]
+WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18]
+WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8]
+WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0]
XI0 NET01 DUM_BL VDD VSS S55NLLGDPH_X512Y8D16_BW_BLSTRAP
XI1 NET01 NET31 DUM_BL VDD VSS WLA[7] WLA[6] WLA[5] WLA[4] WLA[3]
+WLA[2] WLA[1] WLA[0] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST8A_TW
XI2 NET02 NET31 DUM_BL VDD VSS WLA[15] WLA[14] WLA[13] WLA[12] WLA[11]
+WLA[10] WLA[9] WLA[8] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST8A_TW
XI3 NET02 NET32 DUM_BL VDD VSS WLA[23] WLA[22] WLA[21] WLA[20] WLA[19]
+WLA[18] WLA[17] WLA[16] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST8A_TW
XI4 NET03 NET32 DUM_BL VDD VSS WLA[31] WLA[30] WLA[29] WLA[28] WLA[27]
+WLA[26] WLA[25] WLA[24] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST8A_TW
XI5 NET03 NET33 DUM_BL VDD VSS WLA[39] WLA[38] WLA[37] WLA[36] WLA[35]
+WLA[34] WLA[33] WLA[32] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST8A_TW
XI6 NET04 NET33 DUM_BL VDD VSS WLA[47] WLA[46] WLA[45] WLA[44] WLA[43]
+WLA[42] WLA[41] WLA[40] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST8A_TW
XI7 NET04 NET34 DUM_BL VDD VSS WLA[55] WLA[54] WLA[53] WLA[52] WLA[51]
+WLA[50] WLA[49] WLA[48] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST8A_TW
XI8 NET05 NET34 DUM_BL VDD VSS WLA[63] WLA[62] WLA[61] WLA[60] WLA[59]
+WLA[58] WLA[57] WLA[56] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST8A_TW
XI9 NET05 NET4 DUM_BL NET5 VDD VSS VSS STWLA STWLA VSS S55NLLGDPH_X512Y8D16_BW_BITCELL_ST4A_TW
XI10 NET4 NET5 VDD VSS S55NLLGDPH_X512Y8D16_BW_BLSTRAP
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    S55NLLGDPH_X512Y8D16_BW_BITCELL_HSDPH_HVT0974
* View Name:    schematic
************************************************************************

.SUBCKT S55NLLGDPH_X512Y8D16_BW_BITCELL_HSDPH_HVT0974 BA BB BXA BXB VDD VSS WLA WLB
MM4 BB WLB BC VSS DPNPGBHVT W=100.000N L=85.00N M=1
MM2 BXA WLA BCN VSS DPNPGBHVT W=100.000N L=85.00N M=1
MM0 BCN BC VSS VSS DPNPDHVT W=310.00N L=70.00N M=1
MM1 BC BCN VSS VSS DPNPDHVT W=310.00N L=70.00N M=1
MM3 BA WLA BC VSS DPNPGAHVT W=100.000N L=85.00N M=1
MM7 BXB WLB BCN VSS DPNPGAHVT W=100.000N L=85.00N M=1
MM5 BCN BC VDD VDD DPPLHVT W=85.000N L=70.00N M=1
MM6 BC BCN VDD VDD DPPLHVT W=85.000N L=70.00N M=1
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    S55NLLGDPH_X512Y8D16_BW_BITCELL2X2
* View Name:    schematic
************************************************************************

.SUBCKT S55NLLGDPH_X512Y8D16_BW_BITCELL2X2 BA[1] BA[0] BB[1] BB[0] BXA[1] BXA[0] BXB[1] BXB[0] VDD VSS
+WLA[0] WLA[1] WLB[0] WLB[1]
XI8 BA[0] BB[0] BXA[0] BXB[0] VDD VSS WLA[0] WLB[0] S55NLLGDPH_X512Y8D16_BW_BITCELL_HSDPH_HVT0974
XI11 BA[1] BB[1] BXA[1] BXB[1] VDD VSS WLA[1] WLB[1] S55NLLGDPH_X512Y8D16_BW_BITCELL_HSDPH_HVT0974
XI9 BA[0] BB[0] BXA[0] BXB[0] VDD VSS WLA[1] WLB[1] S55NLLGDPH_X512Y8D16_BW_BITCELL_HSDPH_HVT0974
XI10 BA[1] BB[1] BXA[1] BXB[1] VDD VSS WLA[0] WLB[0] S55NLLGDPH_X512Y8D16_BW_BITCELL_HSDPH_HVT0974
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    S55NLLGDPH_X512Y8D16_BW_BITCELL2X8_RD
* View Name:    schematic
************************************************************************

.SUBCKT S55NLLGDPH_X512Y8D16_BW_BITCELL2X8_RD BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[0] WLA[1] WLB[0] WLB[1]
XI11 BLA[3] BLA[2] BLB[3] BLB[2] BLXA[3] BLXA[2] BLXB[3] BLXB[2] VDD VSS 
+ WLA[0] WLA[1] WLB[0] WLB[1] S55NLLGDPH_X512Y8D16_BW_BITCELL2X2
XI12 BLA[5] BLA[4] BLB[5] BLB[4] BLXA[5] BLXA[4] BLXB[5] BLXB[4] VDD VSS 
+ WLA[0] WLA[1] WLB[0] WLB[1] S55NLLGDPH_X512Y8D16_BW_BITCELL2X2
XI13 BLA[7] BLA[6] BLB[7] BLB[6] BLXA[7] BLXA[6] BLXB[7] BLXB[6] VDD VSS 
+ WLA[0] WLA[1] WLB[0] WLB[1] S55NLLGDPH_X512Y8D16_BW_BITCELL2X2
XI0 BLA[1] BLA[0] BLB[1] BLB[0] BLXA[1] BLXA[0] BLXB[1] BLXB[0] VDD VSS WLA[0] 
+ WLA[1] WLB[0] WLB[1] S55NLLGDPH_X512Y8D16_BW_BITCELL2X2
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
* View Name:    schematic
************************************************************************

.SUBCKT S55NLLGDPH_X512Y8D16_BW_BITCELL2X8 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[1] WLA[0] WLB[1] WLB[0]
XI10 BLA[3] BLA[2] BLB[3] BLB[2] BLXA[3] BLXA[2] BLXB[3] BLXB[2] VDD VSS 
+ WLA[0] WLA[1] WLB[0] WLB[1] S55NLLGDPH_X512Y8D16_BW_BITCELL2X2
XI11 BLA[5] BLA[4] BLB[5] BLB[4] BLXA[5] BLXA[4] BLXB[5] BLXB[4] VDD VSS 
+ WLA[0] WLA[1] WLB[0] WLB[1] S55NLLGDPH_X512Y8D16_BW_BITCELL2X2
XI12 BLA[7] BLA[6] BLB[7] BLB[6] BLXA[7] BLXA[6] BLXB[7] BLXB[6] VDD VSS 
+ WLA[0] WLA[1] WLB[0] WLB[1] S55NLLGDPH_X512Y8D16_BW_BITCELL2X2
XI0 BLA[1] BLA[0] BLB[1] BLB[0] BLXA[1] BLXA[0] BLXB[1] BLXB[0] VDD VSS WLA[0] 
+ WLA[1] WLB[0] WLB[1] S55NLLGDPH_X512Y8D16_BW_BITCELL2X2
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    S55NLLGDPH_X512Y8D16_BW_BITCELL66X8B_RED
* View Name:    schematic
************************************************************************

.SUBCKT S55NLLGDPH_X512Y8D16_BW_BITCELL66X8B_RED BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] RWLA[0] RWLA[1] RWLB[0] RWLB[1] VDD VSS WLA[63] WLA[62]
+WLA[61] WLA[60] WLA[59] WLA[58] WLA[57] WLA[56] WLA[55] WLA[54] WLA[53] WLA[52]
+WLA[51] WLA[50] WLA[49] WLA[48] WLA[47] WLA[46] WLA[45] WLA[44] WLA[43] WLA[42]
+WLA[41] WLA[40] WLA[39] WLA[38] WLA[37] WLA[36] WLA[35] WLA[34] WLA[33] WLA[32]
+WLA[31] WLA[30] WLA[29] WLA[28] WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22]
+WLA[21] WLA[20] WLA[19] WLA[18] WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12]
+WLA[11] WLA[10] WLA[9] WLA[8] WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2]
+WLA[1] WLA[0] WLB[63] WLB[62] WLB[61] WLB[60] WLB[59] WLB[58] WLB[57] WLB[56]
+WLB[55] WLB[54] WLB[53] WLB[52] WLB[51] WLB[50] WLB[49] WLB[48] WLB[47] WLB[46]
+WLB[45] WLB[44] WLB[43] WLB[42] WLB[41] WLB[40] WLB[39] WLB[38] WLB[37] WLB[36]
+WLB[35] WLB[34] WLB[33] WLB[32] WLB[31] WLB[30] WLB[29] WLB[28] WLB[27] WLB[26]
+WLB[25] WLB[24] WLB[23] WLB[22] WLB[21] WLB[20] WLB[19] WLB[18] WLB[17] WLB[16]
+WLB[15] WLB[14] WLB[13] WLB[12] WLB[11] WLB[10] WLB[9] WLB[8] WLB[7] WLB[6]
+WLB[5] WLB[4] WLB[3] WLB[2] WLB[1] WLB[0]
XI0 BLA[0] BLXA[0] VDD VSS S55NLLGDPH_X512Y8D16_BW_BLSTRAP_B
XI1 BLA[0] BLXA[0] VDD VSS S55NLLGDPH_X512Y8D16_BW_BLSTRAP_B
XI2 BLA[1] BLXA[1] VDD VSS S55NLLGDPH_X512Y8D16_BW_BLSTRAP_B
XI3 BLA[1] BLXA[1] VDD VSS S55NLLGDPH_X512Y8D16_BW_BLSTRAP_B
XI4 BLA[2] BLXA[2] VDD VSS S55NLLGDPH_X512Y8D16_BW_BLSTRAP_B
XI5 BLA[2] BLXA[2] VDD VSS S55NLLGDPH_X512Y8D16_BW_BLSTRAP_B
XI6 BLA[3] BLXA[3] VDD VSS S55NLLGDPH_X512Y8D16_BW_BLSTRAP_B
XI7 BLA[3] BLXA[3] VDD VSS S55NLLGDPH_X512Y8D16_BW_BLSTRAP_B
XI8 BLA[4] BLXA[4] VDD VSS S55NLLGDPH_X512Y8D16_BW_BLSTRAP_B
XI9 BLA[4] BLXA[4] VDD VSS S55NLLGDPH_X512Y8D16_BW_BLSTRAP_B
XI10 BLA[5] BLXA[5] VDD VSS S55NLLGDPH_X512Y8D16_BW_BLSTRAP_B
XI11 BLA[5] BLXA[5] VDD VSS S55NLLGDPH_X512Y8D16_BW_BLSTRAP_B
XI12 BLA[6] BLXA[6] VDD VSS S55NLLGDPH_X512Y8D16_BW_BLSTRAP_B
XI13 BLA[6] BLXA[6] VDD VSS S55NLLGDPH_X512Y8D16_BW_BLSTRAP_B
XI14 BLA[7] BLXA[7] VDD VSS S55NLLGDPH_X512Y8D16_BW_BLSTRAP_B
XI15 BLA[7] BLXA[7] VDD VSS S55NLLGDPH_X512Y8D16_BW_BLSTRAP_B
XI16 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS RWLA[0] RWLA[1] RWLB[0] RWLB[1] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8_RD
XI17 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[1] WLA[0] WLB[1] WLB[0] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI18 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[3] WLA[2] WLB[3] WLB[2] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI19 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[5] WLA[4] WLB[5] WLB[4] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI20 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[7] WLA[6] WLB[7] WLB[6] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI21 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[9] WLA[8] WLB[9] WLB[8] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI22 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[11] WLA[10] WLB[11] WLB[10] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI23 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[13] WLA[12] WLB[13] WLB[12] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI24 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[15] WLA[14] WLB[15] WLB[14] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI25 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[17] WLA[16] WLB[17] WLB[16] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI26 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[19] WLA[18] WLB[19] WLB[18] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI27 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[21] WLA[20] WLB[21] WLB[20] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI28 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[23] WLA[22] WLB[23] WLB[22] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI29 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[25] WLA[24] WLB[25] WLB[24] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI30 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[27] WLA[26] WLB[27] WLB[26] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI31 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[29] WLA[28] WLB[29] WLB[28] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI32 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[31] WLA[30] WLB[31] WLB[30] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI33 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[33] WLA[32] WLB[33] WLB[32] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI34 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[35] WLA[34] WLB[35] WLB[34] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI35 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[37] WLA[36] WLB[37] WLB[36] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI36 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[39] WLA[38] WLB[39] WLB[38] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI37 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[41] WLA[40] WLB[41] WLB[40] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI38 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[43] WLA[42] WLB[43] WLB[42] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI39 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[45] WLA[44] WLB[45] WLB[44] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI40 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[47] WLA[46] WLB[47] WLB[46] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI41 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[49] WLA[48] WLB[49] WLB[48] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI42 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[51] WLA[50] WLB[51] WLB[50] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI43 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[53] WLA[52] WLB[53] WLB[52] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI44 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[55] WLA[54] WLB[55] WLB[54] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI45 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[57] WLA[56] WLB[57] WLB[56] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI46 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[59] WLA[58] WLB[59] WLB[58] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI47 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[61] WLA[60] WLB[61] WLB[60] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI48 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[63] WLA[62] WLB[63] WLB[62] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    S55NLLGDPH_X512Y8D16_BW_BITCELL64X8A
* View Name:    schematic
************************************************************************

.SUBCKT S55NLLGDPH_X512Y8D16_BW_BITCELL64X8A BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[63] WLA[62] WLA[61] WLA[60] WLA[59] WLA[58]
+WLA[57] WLA[56] WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48]
+WLA[47] WLA[46] WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38]
+WLA[37] WLA[36] WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28]
+WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18]
+WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8]
+WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] WLB[63] WLB[62]
+WLB[61] WLB[60] WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54] WLB[53] WLB[52]
+WLB[51] WLB[50] WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44] WLB[43] WLB[42]
+WLB[41] WLB[40] WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34] WLB[33] WLB[32]
+WLB[31] WLB[30] WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24] WLB[23] WLB[22]
+WLB[21] WLB[20] WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14] WLB[13] WLB[12]
+WLB[11] WLB[10] WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4] WLB[3] WLB[2]
+WLB[1] WLB[0]
XI0 BLB[0] BLXB[0] VDD VSS S55NLLGDPH_X512Y8D16_BW_BLSTRAP
XI1 BLB[0] BLXB[0] VDD VSS S55NLLGDPH_X512Y8D16_BW_BLSTRAP
XI2 BLB[1] BLXB[1] VDD VSS S55NLLGDPH_X512Y8D16_BW_BLSTRAP
XI3 BLB[1] BLXB[1] VDD VSS S55NLLGDPH_X512Y8D16_BW_BLSTRAP
XI4 BLB[2] BLXB[2] VDD VSS S55NLLGDPH_X512Y8D16_BW_BLSTRAP
XI5 BLB[2] BLXB[2] VDD VSS S55NLLGDPH_X512Y8D16_BW_BLSTRAP
XI6 BLB[3] BLXB[3] VDD VSS S55NLLGDPH_X512Y8D16_BW_BLSTRAP
XI7 BLB[3] BLXB[3] VDD VSS S55NLLGDPH_X512Y8D16_BW_BLSTRAP
XI8 BLB[4] BLXB[4] VDD VSS S55NLLGDPH_X512Y8D16_BW_BLSTRAP
XI9 BLB[4] BLXB[4] VDD VSS S55NLLGDPH_X512Y8D16_BW_BLSTRAP
XI10 BLB[5] BLXB[5] VDD VSS S55NLLGDPH_X512Y8D16_BW_BLSTRAP
XI11 BLB[5] BLXB[5] VDD VSS S55NLLGDPH_X512Y8D16_BW_BLSTRAP
XI12 BLB[6] BLXB[6] VDD VSS S55NLLGDPH_X512Y8D16_BW_BLSTRAP
XI13 BLB[6] BLXB[6] VDD VSS S55NLLGDPH_X512Y8D16_BW_BLSTRAP
XI14 BLB[7] BLXB[7] VDD VSS S55NLLGDPH_X512Y8D16_BW_BLSTRAP
XI15 BLB[7] BLXB[7] VDD VSS S55NLLGDPH_X512Y8D16_BW_BLSTRAP
XI16 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[1] WLA[0] WLB[1] WLB[0] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI17 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[3] WLA[2] WLB[3] WLB[2] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI18 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[5] WLA[4] WLB[5] WLB[4] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI19 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[7] WLA[6] WLB[7] WLB[6] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI20 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[9] WLA[8] WLB[9] WLB[8] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI21 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[11] WLA[10] WLB[11] WLB[10] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI22 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[13] WLA[12] WLB[13] WLB[12] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI23 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[15] WLA[14] WLB[15] WLB[14] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI24 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[17] WLA[16] WLB[17] WLB[16] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI25 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[19] WLA[18] WLB[19] WLB[18] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI26 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[21] WLA[20] WLB[21] WLB[20] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI27 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[23] WLA[22] WLB[23] WLB[22] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI28 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[25] WLA[24] WLB[25] WLB[24] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI29 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[27] WLA[26] WLB[27] WLB[26] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI30 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[29] WLA[28] WLB[29] WLB[28] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI31 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[31] WLA[30] WLB[31] WLB[30] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI32 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[33] WLA[32] WLB[33] WLB[32] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI33 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[35] WLA[34] WLB[35] WLB[34] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI34 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[37] WLA[36] WLB[37] WLB[36] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI35 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[39] WLA[38] WLB[39] WLB[38] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI36 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[41] WLA[40] WLB[41] WLB[40] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI37 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[43] WLA[42] WLB[43] WLB[42] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI38 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[45] WLA[44] WLB[45] WLB[44] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI39 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[47] WLA[46] WLB[47] WLB[46] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI40 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[49] WLA[48] WLB[49] WLB[48] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI41 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[51] WLA[50] WLB[51] WLB[50] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI42 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[53] WLA[52] WLB[53] WLB[52] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI43 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[55] WLA[54] WLB[55] WLB[54] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI44 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[57] WLA[56] WLB[57] WLB[56] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI45 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[59] WLA[58] WLB[59] WLB[58] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI46 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[61] WLA[60] WLB[61] WLB[60] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI47 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[63] WLA[62] WLB[63] WLB[62] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    S55NLLGDPH_X512Y8D16_BW_BITCELL64X8B
* View Name:    schematic
************************************************************************

.SUBCKT S55NLLGDPH_X512Y8D16_BW_BITCELL64X8B BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[63] WLA[62] WLA[61] WLA[60] WLA[59] WLA[58]
+WLA[57] WLA[56] WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48]
+WLA[47] WLA[46] WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38]
+WLA[37] WLA[36] WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28]
+WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18]
+WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8]
+WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] WLB[63] WLB[62]
+WLB[61] WLB[60] WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54] WLB[53] WLB[52]
+WLB[51] WLB[50] WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44] WLB[43] WLB[42]
+WLB[41] WLB[40] WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34] WLB[33] WLB[32]
+WLB[31] WLB[30] WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24] WLB[23] WLB[22]
+WLB[21] WLB[20] WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14] WLB[13] WLB[12]
+WLB[11] WLB[10] WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4] WLB[3] WLB[2]
+WLB[1] WLB[0]
XI0 BLA[0] BLXA[0] VDD VSS S55NLLGDPH_X512Y8D16_BW_BLSTRAP_B
XI1 BLA[0] BLXA[0] VDD VSS S55NLLGDPH_X512Y8D16_BW_BLSTRAP_B
XI2 BLA[1] BLXA[1] VDD VSS S55NLLGDPH_X512Y8D16_BW_BLSTRAP_B
XI3 BLA[1] BLXA[1] VDD VSS S55NLLGDPH_X512Y8D16_BW_BLSTRAP_B
XI4 BLA[2] BLXA[2] VDD VSS S55NLLGDPH_X512Y8D16_BW_BLSTRAP_B
XI5 BLA[2] BLXA[2] VDD VSS S55NLLGDPH_X512Y8D16_BW_BLSTRAP_B
XI6 BLA[3] BLXA[3] VDD VSS S55NLLGDPH_X512Y8D16_BW_BLSTRAP_B
XI7 BLA[3] BLXA[3] VDD VSS S55NLLGDPH_X512Y8D16_BW_BLSTRAP_B
XI8 BLA[4] BLXA[4] VDD VSS S55NLLGDPH_X512Y8D16_BW_BLSTRAP_B
XI9 BLA[4] BLXA[4] VDD VSS S55NLLGDPH_X512Y8D16_BW_BLSTRAP_B
XI10 BLA[5] BLXA[5] VDD VSS S55NLLGDPH_X512Y8D16_BW_BLSTRAP_B
XI11 BLA[5] BLXA[5] VDD VSS S55NLLGDPH_X512Y8D16_BW_BLSTRAP_B
XI12 BLA[6] BLXA[6] VDD VSS S55NLLGDPH_X512Y8D16_BW_BLSTRAP_B
XI13 BLA[6] BLXA[6] VDD VSS S55NLLGDPH_X512Y8D16_BW_BLSTRAP_B
XI14 BLA[7] BLXA[7] VDD VSS S55NLLGDPH_X512Y8D16_BW_BLSTRAP_B
XI15 BLA[7] BLXA[7] VDD VSS S55NLLGDPH_X512Y8D16_BW_BLSTRAP_B
XI16 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[1] WLA[0] WLB[1] WLB[0] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI17 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[3] WLA[2] WLB[3] WLB[2] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI18 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[5] WLA[4] WLB[5] WLB[4] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI19 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[7] WLA[6] WLB[7] WLB[6] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI20 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[9] WLA[8] WLB[9] WLB[8] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI21 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[11] WLA[10] WLB[11] WLB[10] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI22 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[13] WLA[12] WLB[13] WLB[12] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI23 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[15] WLA[14] WLB[15] WLB[14] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI24 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[17] WLA[16] WLB[17] WLB[16] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI25 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[19] WLA[18] WLB[19] WLB[18] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI26 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[21] WLA[20] WLB[21] WLB[20] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI27 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[23] WLA[22] WLB[23] WLB[22] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI28 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[25] WLA[24] WLB[25] WLB[24] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI29 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[27] WLA[26] WLB[27] WLB[26] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI30 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[29] WLA[28] WLB[29] WLB[28] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI31 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[31] WLA[30] WLB[31] WLB[30] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI32 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[33] WLA[32] WLB[33] WLB[32] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI33 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[35] WLA[34] WLB[35] WLB[34] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI34 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[37] WLA[36] WLB[37] WLB[36] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI35 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[39] WLA[38] WLB[39] WLB[38] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI36 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[41] WLA[40] WLB[41] WLB[40] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI37 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[43] WLA[42] WLB[43] WLB[42] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI38 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[45] WLA[44] WLB[45] WLB[44] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI39 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[47] WLA[46] WLB[47] WLB[46] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI40 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[49] WLA[48] WLB[49] WLB[48] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI41 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[51] WLA[50] WLB[51] WLB[50] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI42 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[53] WLA[52] WLB[53] WLB[52] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI43 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[55] WLA[54] WLB[55] WLB[54] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI44 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[57] WLA[56] WLB[57] WLB[56] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI45 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[59] WLA[58] WLB[59] WLB[58] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI46 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[61] WLA[60] WLB[61] WLB[60] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI47 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[63] WLA[62] WLB[63] WLB[62] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    S55NLLGDPH_X512Y8D16_BW_BITCELL2X2_STWL
* View Name:    schematic
************************************************************************

.SUBCKT S55NLLGDPH_X512Y8D16_BW_BITCELL2X2_STWL BB0 BB3 BXB0 BXB3 VDD VSS WLA[3] WLA[2] WLA[1] WLA[0]
+WLB[3] WLB[2] WLB[1] WLB[0]
XI8 NET72 BB0 NET71 BXB0 VDD VSS WLA[0] WLB[0] S55NLLGDPH_X512Y8D16_BW_BITCELL_HSDPH_HVT0974
XI11 NET64 BB3 NET63 BXB3 VDD VSS WLA[3] WLB[3] S55NLLGDPH_X512Y8D16_BW_BITCELL_HSDPH_HVT0974
XI9 NET72 NET78 NET71 NET77 VDD VSS WLA[1] WLB[1] S55NLLGDPH_X512Y8D16_BW_BITCELL_HSDPH_HVT0974
XI10 NET64 NET78 NET63 NET77 VDD VSS WLA[2] WLB[2] S55NLLGDPH_X512Y8D16_BW_BITCELL_HSDPH_HVT0974
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    S55NLLGDPH_X512Y8D16_BW_BITCELL68X8A_NOMID_TOP
* View Name:    schematic
************************************************************************

.SUBCKT S55NLLGDPH_X512Y8D16_BW_BITCELL68X8A_NOMID_TOP BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] RDWLA[3] RDWLA[2] RDWLA[1] RDWLA[0] RDWLB[3] RDWLB[2] RDWLB[1] RDWLB[0]
+VDD VSS WLA[63] WLA[62] WLA[61] WLA[60] WLA[59] WLA[58] WLA[57] WLA[56]
+WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48] WLA[47] WLA[46]
+WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38] WLA[37] WLA[36]
+WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28] WLA[27] WLA[26]
+WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18] WLA[17] WLA[16]
+WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8] WLA[7] WLA[6]
+WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] WLB[63] WLB[62] WLB[61] WLB[60]
+WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54] WLB[53] WLB[52] WLB[51] WLB[50]
+WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44] WLB[43] WLB[42] WLB[41] WLB[40]
+WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34] WLB[33] WLB[32] WLB[31] WLB[30]
+WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24] WLB[23] WLB[22] WLB[21] WLB[20]
+WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14] WLB[13] WLB[12] WLB[11] WLB[10]
+WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4] WLB[3] WLB[2] WLB[1] WLB[0]
XI0 BLB[0] NET033[8] BLXB[0] NET035[8] VDD VSS RDWLA[3] RDWLA[2] RDWLA[1] RDWLA[0]
+RDWLB[3] RDWLB[2] RDWLB[1] RDWLB[0] S55NLLGDPH_X512Y8D16_BW_BITCELL2X2_STWL
XI1 BLB[0] BLXB[0] VDD VSS S55NLLGDPH_X512Y8D16_BW_BLSTRAP
XI2 NET033[8] NET035[8] VDD VSS S55NLLGDPH_X512Y8D16_BW_BLSTRAP
XI3 BLB[1] NET033[7] BLXB[1] NET035[7] VDD VSS RDWLA[3] RDWLA[2] RDWLA[1] RDWLA[0]
+RDWLB[3] RDWLB[2] RDWLB[1] RDWLB[0] S55NLLGDPH_X512Y8D16_BW_BITCELL2X2_STWL
XI4 BLB[1] BLXB[1] VDD VSS S55NLLGDPH_X512Y8D16_BW_BLSTRAP
XI5 NET033[7] NET035[7] VDD VSS S55NLLGDPH_X512Y8D16_BW_BLSTRAP
XI6 BLB[2] NET033[6] BLXB[2] NET035[6] VDD VSS RDWLA[3] RDWLA[2] RDWLA[1] RDWLA[0]
+RDWLB[3] RDWLB[2] RDWLB[1] RDWLB[0] S55NLLGDPH_X512Y8D16_BW_BITCELL2X2_STWL
XI7 BLB[2] BLXB[2] VDD VSS S55NLLGDPH_X512Y8D16_BW_BLSTRAP
XI8 NET033[6] NET035[6] VDD VSS S55NLLGDPH_X512Y8D16_BW_BLSTRAP
XI9 BLB[3] NET033[5] BLXB[3] NET035[5] VDD VSS RDWLA[3] RDWLA[2] RDWLA[1] RDWLA[0]
+RDWLB[3] RDWLB[2] RDWLB[1] RDWLB[0] S55NLLGDPH_X512Y8D16_BW_BITCELL2X2_STWL
XI10 BLB[3] BLXB[3] VDD VSS S55NLLGDPH_X512Y8D16_BW_BLSTRAP
XI11 NET033[5] NET035[5] VDD VSS S55NLLGDPH_X512Y8D16_BW_BLSTRAP
XI12 BLB[4] NET033[4] BLXB[4] NET035[4] VDD VSS RDWLA[3] RDWLA[2] RDWLA[1] RDWLA[0]
+RDWLB[3] RDWLB[2] RDWLB[1] RDWLB[0] S55NLLGDPH_X512Y8D16_BW_BITCELL2X2_STWL
XI13 BLB[4] BLXB[4] VDD VSS S55NLLGDPH_X512Y8D16_BW_BLSTRAP
XI14 NET033[4] NET035[4] VDD VSS S55NLLGDPH_X512Y8D16_BW_BLSTRAP
XI15 BLB[5] NET033[3] BLXB[5] NET035[3] VDD VSS RDWLA[3] RDWLA[2] RDWLA[1] RDWLA[0]
+RDWLB[3] RDWLB[2] RDWLB[1] RDWLB[0] S55NLLGDPH_X512Y8D16_BW_BITCELL2X2_STWL
XI16 BLB[5] BLXB[5] VDD VSS S55NLLGDPH_X512Y8D16_BW_BLSTRAP
XI17 NET033[3] NET035[3] VDD VSS S55NLLGDPH_X512Y8D16_BW_BLSTRAP
XI18 BLB[6] NET033[2] BLXB[6] NET035[2] VDD VSS RDWLA[3] RDWLA[2] RDWLA[1] RDWLA[0]
+RDWLB[3] RDWLB[2] RDWLB[1] RDWLB[0] S55NLLGDPH_X512Y8D16_BW_BITCELL2X2_STWL
XI19 BLB[6] BLXB[6] VDD VSS S55NLLGDPH_X512Y8D16_BW_BLSTRAP
XI20 NET033[2] NET035[2] VDD VSS S55NLLGDPH_X512Y8D16_BW_BLSTRAP
XI21 BLB[7] NET033[1] BLXB[7] NET035[1] VDD VSS RDWLA[3] RDWLA[2] RDWLA[1] RDWLA[0]
+RDWLB[3] RDWLB[2] RDWLB[1] RDWLB[0] S55NLLGDPH_X512Y8D16_BW_BITCELL2X2_STWL
XI22 BLB[7] BLXB[7] VDD VSS S55NLLGDPH_X512Y8D16_BW_BLSTRAP
XI23 NET033[1] NET035[1] VDD VSS S55NLLGDPH_X512Y8D16_BW_BLSTRAP
XI24 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[1] WLA[0] WLB[1] WLB[0] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI25 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[3] WLA[2] WLB[3] WLB[2] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI26 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[5] WLA[4] WLB[5] WLB[4] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI27 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[7] WLA[6] WLB[7] WLB[6] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI28 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[9] WLA[8] WLB[9] WLB[8] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI29 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[11] WLA[10] WLB[11] WLB[10] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI30 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[13] WLA[12] WLB[13] WLB[12] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI31 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[15] WLA[14] WLB[15] WLB[14] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI32 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[17] WLA[16] WLB[17] WLB[16] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI33 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[19] WLA[18] WLB[19] WLB[18] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI34 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[21] WLA[20] WLB[21] WLB[20] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI35 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[23] WLA[22] WLB[23] WLB[22] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI36 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[25] WLA[24] WLB[25] WLB[24] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI37 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[27] WLA[26] WLB[27] WLB[26] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI38 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[29] WLA[28] WLB[29] WLB[28] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI39 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[31] WLA[30] WLB[31] WLB[30] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI40 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[33] WLA[32] WLB[33] WLB[32] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI41 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[35] WLA[34] WLB[35] WLB[34] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI42 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[37] WLA[36] WLB[37] WLB[36] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI43 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[39] WLA[38] WLB[39] WLB[38] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI44 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[41] WLA[40] WLB[41] WLB[40] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI45 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[43] WLA[42] WLB[43] WLB[42] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI46 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[45] WLA[44] WLB[45] WLB[44] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI47 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[47] WLA[46] WLB[47] WLB[46] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI48 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[49] WLA[48] WLB[49] WLB[48] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI49 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[51] WLA[50] WLB[51] WLB[50] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI50 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[53] WLA[52] WLB[53] WLB[52] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI51 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[55] WLA[54] WLB[55] WLB[54] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI52 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[57] WLA[56] WLB[57] WLB[56] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI53 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[59] WLA[58] WLB[59] WLB[58] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI54 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[61] WLA[60] WLB[61] WLB[60] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI55 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[63] WLA[62] WLB[63] WLB[62] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    S55NLLGDPH_X512Y8D16_BW_ARRAY512X8
* View Name:    schematic
************************************************************************

.SUBCKT S55NLLGDPH_X512Y8D16_BW_ARRAY512X8 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] RDWLA[3] RDWLA[2] RDWLA[1] RDWLA[0] RDWLB[3] RDWLB[2] RDWLB[1] RDWLB[0]
+RWLA[0] RWLA[1] RWLB[0] RWLB[1] VDD VSS WLA[511] WLA[510] WLA[509] WLA[508]
+WLA[507] WLA[506] WLA[505] WLA[504] WLA[503] WLA[502] WLA[501] WLA[500] WLA[499] WLA[498]
+WLA[497] WLA[496] WLA[495] WLA[494] WLA[493] WLA[492] WLA[491] WLA[490] WLA[489] WLA[488]
+WLA[487] WLA[486] WLA[485] WLA[484] WLA[483] WLA[482] WLA[481] WLA[480] WLA[479] WLA[478]
+WLA[477] WLA[476] WLA[475] WLA[474] WLA[473] WLA[472] WLA[471] WLA[470] WLA[469] WLA[468]
+WLA[467] WLA[466] WLA[465] WLA[464] WLA[463] WLA[462] WLA[461] WLA[460] WLA[459] WLA[458]
+WLA[457] WLA[456] WLA[455] WLA[454] WLA[453] WLA[452] WLA[451] WLA[450] WLA[449] WLA[448]
+WLA[447] WLA[446] WLA[445] WLA[444] WLA[443] WLA[442] WLA[441] WLA[440] WLA[439] WLA[438]
+WLA[437] WLA[436] WLA[435] WLA[434] WLA[433] WLA[432] WLA[431] WLA[430] WLA[429] WLA[428]
+WLA[427] WLA[426] WLA[425] WLA[424] WLA[423] WLA[422] WLA[421] WLA[420] WLA[419] WLA[418]
+WLA[417] WLA[416] WLA[415] WLA[414] WLA[413] WLA[412] WLA[411] WLA[410] WLA[409] WLA[408]
+WLA[407] WLA[406] WLA[405] WLA[404] WLA[403] WLA[402] WLA[401] WLA[400] WLA[399] WLA[398]
+WLA[397] WLA[396] WLA[395] WLA[394] WLA[393] WLA[392] WLA[391] WLA[390] WLA[389] WLA[388]
+WLA[387] WLA[386] WLA[385] WLA[384] WLA[383] WLA[382] WLA[381] WLA[380] WLA[379] WLA[378]
+WLA[377] WLA[376] WLA[375] WLA[374] WLA[373] WLA[372] WLA[371] WLA[370] WLA[369] WLA[368]
+WLA[367] WLA[366] WLA[365] WLA[364] WLA[363] WLA[362] WLA[361] WLA[360] WLA[359] WLA[358]
+WLA[357] WLA[356] WLA[355] WLA[354] WLA[353] WLA[352] WLA[351] WLA[350] WLA[349] WLA[348]
+WLA[347] WLA[346] WLA[345] WLA[344] WLA[343] WLA[342] WLA[341] WLA[340] WLA[339] WLA[338]
+WLA[337] WLA[336] WLA[335] WLA[334] WLA[333] WLA[332] WLA[331] WLA[330] WLA[329] WLA[328]
+WLA[327] WLA[326] WLA[325] WLA[324] WLA[323] WLA[322] WLA[321] WLA[320] WLA[319] WLA[318]
+WLA[317] WLA[316] WLA[315] WLA[314] WLA[313] WLA[312] WLA[311] WLA[310] WLA[309] WLA[308]
+WLA[307] WLA[306] WLA[305] WLA[304] WLA[303] WLA[302] WLA[301] WLA[300] WLA[299] WLA[298]
+WLA[297] WLA[296] WLA[295] WLA[294] WLA[293] WLA[292] WLA[291] WLA[290] WLA[289] WLA[288]
+WLA[287] WLA[286] WLA[285] WLA[284] WLA[283] WLA[282] WLA[281] WLA[280] WLA[279] WLA[278]
+WLA[277] WLA[276] WLA[275] WLA[274] WLA[273] WLA[272] WLA[271] WLA[270] WLA[269] WLA[268]
+WLA[267] WLA[266] WLA[265] WLA[264] WLA[263] WLA[262] WLA[261] WLA[260] WLA[259] WLA[258]
+WLA[257] WLA[256] WLA[255] WLA[254] WLA[253] WLA[252] WLA[251] WLA[250] WLA[249] WLA[248]
+WLA[247] WLA[246] WLA[245] WLA[244] WLA[243] WLA[242] WLA[241] WLA[240] WLA[239] WLA[238]
+WLA[237] WLA[236] WLA[235] WLA[234] WLA[233] WLA[232] WLA[231] WLA[230] WLA[229] WLA[228]
+WLA[227] WLA[226] WLA[225] WLA[224] WLA[223] WLA[222] WLA[221] WLA[220] WLA[219] WLA[218]
+WLA[217] WLA[216] WLA[215] WLA[214] WLA[213] WLA[212] WLA[211] WLA[210] WLA[209] WLA[208]
+WLA[207] WLA[206] WLA[205] WLA[204] WLA[203] WLA[202] WLA[201] WLA[200] WLA[199] WLA[198]
+WLA[197] WLA[196] WLA[195] WLA[194] WLA[193] WLA[192] WLA[191] WLA[190] WLA[189] WLA[188]
+WLA[187] WLA[186] WLA[185] WLA[184] WLA[183] WLA[182] WLA[181] WLA[180] WLA[179] WLA[178]
+WLA[177] WLA[176] WLA[175] WLA[174] WLA[173] WLA[172] WLA[171] WLA[170] WLA[169] WLA[168]
+WLA[167] WLA[166] WLA[165] WLA[164] WLA[163] WLA[162] WLA[161] WLA[160] WLA[159] WLA[158]
+WLA[157] WLA[156] WLA[155] WLA[154] WLA[153] WLA[152] WLA[151] WLA[150] WLA[149] WLA[148]
+WLA[147] WLA[146] WLA[145] WLA[144] WLA[143] WLA[142] WLA[141] WLA[140] WLA[139] WLA[138]
+WLA[137] WLA[136] WLA[135] WLA[134] WLA[133] WLA[132] WLA[131] WLA[130] WLA[129] WLA[128]
+WLA[127] WLA[126] WLA[125] WLA[124] WLA[123] WLA[122] WLA[121] WLA[120] WLA[119] WLA[118]
+WLA[117] WLA[116] WLA[115] WLA[114] WLA[113] WLA[112] WLA[111] WLA[110] WLA[109] WLA[108]
+WLA[107] WLA[106] WLA[105] WLA[104] WLA[103] WLA[102] WLA[101] WLA[100] WLA[99] WLA[98]
+WLA[97] WLA[96] WLA[95] WLA[94] WLA[93] WLA[92] WLA[91] WLA[90] WLA[89] WLA[88]
+WLA[87] WLA[86] WLA[85] WLA[84] WLA[83] WLA[82] WLA[81] WLA[80] WLA[79] WLA[78]
+WLA[77] WLA[76] WLA[75] WLA[74] WLA[73] WLA[72] WLA[71] WLA[70] WLA[69] WLA[68]
+WLA[67] WLA[66] WLA[65] WLA[64] WLA[63] WLA[62] WLA[61] WLA[60] WLA[59] WLA[58]
+WLA[57] WLA[56] WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48]
+WLA[47] WLA[46] WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38]
+WLA[37] WLA[36] WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28]
+WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18]
+WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8]
+WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] WLB[511] WLB[510]
+WLB[509] WLB[508] WLB[507] WLB[506] WLB[505] WLB[504] WLB[503] WLB[502] WLB[501] WLB[500]
+WLB[499] WLB[498] WLB[497] WLB[496] WLB[495] WLB[494] WLB[493] WLB[492] WLB[491] WLB[490]
+WLB[489] WLB[488] WLB[487] WLB[486] WLB[485] WLB[484] WLB[483] WLB[482] WLB[481] WLB[480]
+WLB[479] WLB[478] WLB[477] WLB[476] WLB[475] WLB[474] WLB[473] WLB[472] WLB[471] WLB[470]
+WLB[469] WLB[468] WLB[467] WLB[466] WLB[465] WLB[464] WLB[463] WLB[462] WLB[461] WLB[460]
+WLB[459] WLB[458] WLB[457] WLB[456] WLB[455] WLB[454] WLB[453] WLB[452] WLB[451] WLB[450]
+WLB[449] WLB[448] WLB[447] WLB[446] WLB[445] WLB[444] WLB[443] WLB[442] WLB[441] WLB[440]
+WLB[439] WLB[438] WLB[437] WLB[436] WLB[435] WLB[434] WLB[433] WLB[432] WLB[431] WLB[430]
+WLB[429] WLB[428] WLB[427] WLB[426] WLB[425] WLB[424] WLB[423] WLB[422] WLB[421] WLB[420]
+WLB[419] WLB[418] WLB[417] WLB[416] WLB[415] WLB[414] WLB[413] WLB[412] WLB[411] WLB[410]
+WLB[409] WLB[408] WLB[407] WLB[406] WLB[405] WLB[404] WLB[403] WLB[402] WLB[401] WLB[400]
+WLB[399] WLB[398] WLB[397] WLB[396] WLB[395] WLB[394] WLB[393] WLB[392] WLB[391] WLB[390]
+WLB[389] WLB[388] WLB[387] WLB[386] WLB[385] WLB[384] WLB[383] WLB[382] WLB[381] WLB[380]
+WLB[379] WLB[378] WLB[377] WLB[376] WLB[375] WLB[374] WLB[373] WLB[372] WLB[371] WLB[370]
+WLB[369] WLB[368] WLB[367] WLB[366] WLB[365] WLB[364] WLB[363] WLB[362] WLB[361] WLB[360]
+WLB[359] WLB[358] WLB[357] WLB[356] WLB[355] WLB[354] WLB[353] WLB[352] WLB[351] WLB[350]
+WLB[349] WLB[348] WLB[347] WLB[346] WLB[345] WLB[344] WLB[343] WLB[342] WLB[341] WLB[340]
+WLB[339] WLB[338] WLB[337] WLB[336] WLB[335] WLB[334] WLB[333] WLB[332] WLB[331] WLB[330]
+WLB[329] WLB[328] WLB[327] WLB[326] WLB[325] WLB[324] WLB[323] WLB[322] WLB[321] WLB[320]
+WLB[319] WLB[318] WLB[317] WLB[316] WLB[315] WLB[314] WLB[313] WLB[312] WLB[311] WLB[310]
+WLB[309] WLB[308] WLB[307] WLB[306] WLB[305] WLB[304] WLB[303] WLB[302] WLB[301] WLB[300]
+WLB[299] WLB[298] WLB[297] WLB[296] WLB[295] WLB[294] WLB[293] WLB[292] WLB[291] WLB[290]
+WLB[289] WLB[288] WLB[287] WLB[286] WLB[285] WLB[284] WLB[283] WLB[282] WLB[281] WLB[280]
+WLB[279] WLB[278] WLB[277] WLB[276] WLB[275] WLB[274] WLB[273] WLB[272] WLB[271] WLB[270]
+WLB[269] WLB[268] WLB[267] WLB[266] WLB[265] WLB[264] WLB[263] WLB[262] WLB[261] WLB[260]
+WLB[259] WLB[258] WLB[257] WLB[256] WLB[255] WLB[254] WLB[253] WLB[252] WLB[251] WLB[250]
+WLB[249] WLB[248] WLB[247] WLB[246] WLB[245] WLB[244] WLB[243] WLB[242] WLB[241] WLB[240]
+WLB[239] WLB[238] WLB[237] WLB[236] WLB[235] WLB[234] WLB[233] WLB[232] WLB[231] WLB[230]
+WLB[229] WLB[228] WLB[227] WLB[226] WLB[225] WLB[224] WLB[223] WLB[222] WLB[221] WLB[220]
+WLB[219] WLB[218] WLB[217] WLB[216] WLB[215] WLB[214] WLB[213] WLB[212] WLB[211] WLB[210]
+WLB[209] WLB[208] WLB[207] WLB[206] WLB[205] WLB[204] WLB[203] WLB[202] WLB[201] WLB[200]
+WLB[199] WLB[198] WLB[197] WLB[196] WLB[195] WLB[194] WLB[193] WLB[192] WLB[191] WLB[190]
+WLB[189] WLB[188] WLB[187] WLB[186] WLB[185] WLB[184] WLB[183] WLB[182] WLB[181] WLB[180]
+WLB[179] WLB[178] WLB[177] WLB[176] WLB[175] WLB[174] WLB[173] WLB[172] WLB[171] WLB[170]
+WLB[169] WLB[168] WLB[167] WLB[166] WLB[165] WLB[164] WLB[163] WLB[162] WLB[161] WLB[160]
+WLB[159] WLB[158] WLB[157] WLB[156] WLB[155] WLB[154] WLB[153] WLB[152] WLB[151] WLB[150]
+WLB[149] WLB[148] WLB[147] WLB[146] WLB[145] WLB[144] WLB[143] WLB[142] WLB[141] WLB[140]
+WLB[139] WLB[138] WLB[137] WLB[136] WLB[135] WLB[134] WLB[133] WLB[132] WLB[131] WLB[130]
+WLB[129] WLB[128] WLB[127] WLB[126] WLB[125] WLB[124] WLB[123] WLB[122] WLB[121] WLB[120]
+WLB[119] WLB[118] WLB[117] WLB[116] WLB[115] WLB[114] WLB[113] WLB[112] WLB[111] WLB[110]
+WLB[109] WLB[108] WLB[107] WLB[106] WLB[105] WLB[104] WLB[103] WLB[102] WLB[101] WLB[100]
+WLB[99] WLB[98] WLB[97] WLB[96] WLB[95] WLB[94] WLB[93] WLB[92] WLB[91] WLB[90]
+WLB[89] WLB[88] WLB[87] WLB[86] WLB[85] WLB[84] WLB[83] WLB[82] WLB[81] WLB[80]
+WLB[79] WLB[78] WLB[77] WLB[76] WLB[75] WLB[74] WLB[73] WLB[72] WLB[71] WLB[70]
+WLB[69] WLB[68] WLB[67] WLB[66] WLB[65] WLB[64] WLB[63] WLB[62] WLB[61] WLB[60]
+WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54] WLB[53] WLB[52] WLB[51] WLB[50]
+WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44] WLB[43] WLB[42] WLB[41] WLB[40]
+WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34] WLB[33] WLB[32] WLB[31] WLB[30]
+WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24] WLB[23] WLB[22] WLB[21] WLB[20]
+WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14] WLB[13] WLB[12] WLB[11] WLB[10]
+WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4] WLB[3] WLB[2] WLB[1] WLB[0]
XI0 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] RWLA[0] RWLA[1] RWLB[0] RWLB[1] VDD VSS WLA[63] WLA[62]
+WLA[61] WLA[60] WLA[59] WLA[58] WLA[57] WLA[56] WLA[55] WLA[54] WLA[53] WLA[52]
+WLA[51] WLA[50] WLA[49] WLA[48] WLA[47] WLA[46] WLA[45] WLA[44] WLA[43] WLA[42]
+WLA[41] WLA[40] WLA[39] WLA[38] WLA[37] WLA[36] WLA[35] WLA[34] WLA[33] WLA[32]
+WLA[31] WLA[30] WLA[29] WLA[28] WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22]
+WLA[21] WLA[20] WLA[19] WLA[18] WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12]
+WLA[11] WLA[10] WLA[9] WLA[8] WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2]
+WLA[1] WLA[0] WLB[63] WLB[62] WLB[61] WLB[60] WLB[59] WLB[58] WLB[57] WLB[56]
+WLB[55] WLB[54] WLB[53] WLB[52] WLB[51] WLB[50] WLB[49] WLB[48] WLB[47] WLB[46]
+WLB[45] WLB[44] WLB[43] WLB[42] WLB[41] WLB[40] WLB[39] WLB[38] WLB[37] WLB[36]
+WLB[35] WLB[34] WLB[33] WLB[32] WLB[31] WLB[30] WLB[29] WLB[28] WLB[27] WLB[26]
+WLB[25] WLB[24] WLB[23] WLB[22] WLB[21] WLB[20] WLB[19] WLB[18] WLB[17] WLB[16]
+WLB[15] WLB[14] WLB[13] WLB[12] WLB[11] WLB[10] WLB[9] WLB[8] WLB[7] WLB[6]
+WLB[5] WLB[4] WLB[3] WLB[2] WLB[1] WLB[0] S55NLLGDPH_X512Y8D16_BW_BITCELL66X8B_RED
XI1 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[127] WLA[126] WLA[125] WLA[124] WLA[123] WLA[122]
+WLA[121] WLA[120] WLA[119] WLA[118] WLA[117] WLA[116] WLA[115] WLA[114] WLA[113] WLA[112]
+WLA[111] WLA[110] WLA[109] WLA[108] WLA[107] WLA[106] WLA[105] WLA[104] WLA[103] WLA[102]
+WLA[101] WLA[100] WLA[99] WLA[98] WLA[97] WLA[96] WLA[95] WLA[94] WLA[93] WLA[92]
+WLA[91] WLA[90] WLA[89] WLA[88] WLA[87] WLA[86] WLA[85] WLA[84] WLA[83] WLA[82]
+WLA[81] WLA[80] WLA[79] WLA[78] WLA[77] WLA[76] WLA[75] WLA[74] WLA[73] WLA[72]
+WLA[71] WLA[70] WLA[69] WLA[68] WLA[67] WLA[66] WLA[65] WLA[64] WLB[127] WLB[126]
+WLB[125] WLB[124] WLB[123] WLB[122] WLB[121] WLB[120] WLB[119] WLB[118] WLB[117] WLB[116]
+WLB[115] WLB[114] WLB[113] WLB[112] WLB[111] WLB[110] WLB[109] WLB[108] WLB[107] WLB[106]
+WLB[105] WLB[104] WLB[103] WLB[102] WLB[101] WLB[100] WLB[99] WLB[98] WLB[97] WLB[96]
+WLB[95] WLB[94] WLB[93] WLB[92] WLB[91] WLB[90] WLB[89] WLB[88] WLB[87] WLB[86]
+WLB[85] WLB[84] WLB[83] WLB[82] WLB[81] WLB[80] WLB[79] WLB[78] WLB[77] WLB[76]
+WLB[75] WLB[74] WLB[73] WLB[72] WLB[71] WLB[70] WLB[69] WLB[68] WLB[67] WLB[66]
+WLB[65] WLB[64] S55NLLGDPH_X512Y8D16_BW_BITCELL64X8A
XI2 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[191] WLA[190] WLA[189] WLA[188] WLA[187] WLA[186]
+WLA[185] WLA[184] WLA[183] WLA[182] WLA[181] WLA[180] WLA[179] WLA[178] WLA[177] WLA[176]
+WLA[175] WLA[174] WLA[173] WLA[172] WLA[171] WLA[170] WLA[169] WLA[168] WLA[167] WLA[166]
+WLA[165] WLA[164] WLA[163] WLA[162] WLA[161] WLA[160] WLA[159] WLA[158] WLA[157] WLA[156]
+WLA[155] WLA[154] WLA[153] WLA[152] WLA[151] WLA[150] WLA[149] WLA[148] WLA[147] WLA[146]
+WLA[145] WLA[144] WLA[143] WLA[142] WLA[141] WLA[140] WLA[139] WLA[138] WLA[137] WLA[136]
+WLA[135] WLA[134] WLA[133] WLA[132] WLA[131] WLA[130] WLA[129] WLA[128] WLB[191] WLB[190]
+WLB[189] WLB[188] WLB[187] WLB[186] WLB[185] WLB[184] WLB[183] WLB[182] WLB[181] WLB[180]
+WLB[179] WLB[178] WLB[177] WLB[176] WLB[175] WLB[174] WLB[173] WLB[172] WLB[171] WLB[170]
+WLB[169] WLB[168] WLB[167] WLB[166] WLB[165] WLB[164] WLB[163] WLB[162] WLB[161] WLB[160]
+WLB[159] WLB[158] WLB[157] WLB[156] WLB[155] WLB[154] WLB[153] WLB[152] WLB[151] WLB[150]
+WLB[149] WLB[148] WLB[147] WLB[146] WLB[145] WLB[144] WLB[143] WLB[142] WLB[141] WLB[140]
+WLB[139] WLB[138] WLB[137] WLB[136] WLB[135] WLB[134] WLB[133] WLB[132] WLB[131] WLB[130]
+WLB[129] WLB[128] S55NLLGDPH_X512Y8D16_BW_BITCELL64X8B
XI3 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[255] WLA[254] WLA[253] WLA[252] WLA[251] WLA[250]
+WLA[249] WLA[248] WLA[247] WLA[246] WLA[245] WLA[244] WLA[243] WLA[242] WLA[241] WLA[240]
+WLA[239] WLA[238] WLA[237] WLA[236] WLA[235] WLA[234] WLA[233] WLA[232] WLA[231] WLA[230]
+WLA[229] WLA[228] WLA[227] WLA[226] WLA[225] WLA[224] WLA[223] WLA[222] WLA[221] WLA[220]
+WLA[219] WLA[218] WLA[217] WLA[216] WLA[215] WLA[214] WLA[213] WLA[212] WLA[211] WLA[210]
+WLA[209] WLA[208] WLA[207] WLA[206] WLA[205] WLA[204] WLA[203] WLA[202] WLA[201] WLA[200]
+WLA[199] WLA[198] WLA[197] WLA[196] WLA[195] WLA[194] WLA[193] WLA[192] WLB[255] WLB[254]
+WLB[253] WLB[252] WLB[251] WLB[250] WLB[249] WLB[248] WLB[247] WLB[246] WLB[245] WLB[244]
+WLB[243] WLB[242] WLB[241] WLB[240] WLB[239] WLB[238] WLB[237] WLB[236] WLB[235] WLB[234]
+WLB[233] WLB[232] WLB[231] WLB[230] WLB[229] WLB[228] WLB[227] WLB[226] WLB[225] WLB[224]
+WLB[223] WLB[222] WLB[221] WLB[220] WLB[219] WLB[218] WLB[217] WLB[216] WLB[215] WLB[214]
+WLB[213] WLB[212] WLB[211] WLB[210] WLB[209] WLB[208] WLB[207] WLB[206] WLB[205] WLB[204]
+WLB[203] WLB[202] WLB[201] WLB[200] WLB[199] WLB[198] WLB[197] WLB[196] WLB[195] WLB[194]
+WLB[193] WLB[192] S55NLLGDPH_X512Y8D16_BW_BITCELL64X8A
XI4 BLXA[7] BLXA[6] BLXA[5] BLXA[4] BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6]
+BLXB[5] BLXB[4] BLXB[3] BLXB[2] BLXB[1] BLXB[0] BLA[7] BLA[6] BLA[5] BLA[4]
+BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6] BLB[5] BLB[4] BLB[3] BLB[2]
+BLB[1] BLB[0] VDD VSS WLA[319] WLA[318] WLA[317] WLA[316] WLA[315] WLA[314]
+WLA[313] WLA[312] WLA[311] WLA[310] WLA[309] WLA[308] WLA[307] WLA[306] WLA[305] WLA[304]
+WLA[303] WLA[302] WLA[301] WLA[300] WLA[299] WLA[298] WLA[297] WLA[296] WLA[295] WLA[294]
+WLA[293] WLA[292] WLA[291] WLA[290] WLA[289] WLA[288] WLA[287] WLA[286] WLA[285] WLA[284]
+WLA[283] WLA[282] WLA[281] WLA[280] WLA[279] WLA[278] WLA[277] WLA[276] WLA[275] WLA[274]
+WLA[273] WLA[272] WLA[271] WLA[270] WLA[269] WLA[268] WLA[267] WLA[266] WLA[265] WLA[264]
+WLA[263] WLA[262] WLA[261] WLA[260] WLA[259] WLA[258] WLA[257] WLA[256] WLB[319] WLB[318]
+WLB[317] WLB[316] WLB[315] WLB[314] WLB[313] WLB[312] WLB[311] WLB[310] WLB[309] WLB[308]
+WLB[307] WLB[306] WLB[305] WLB[304] WLB[303] WLB[302] WLB[301] WLB[300] WLB[299] WLB[298]
+WLB[297] WLB[296] WLB[295] WLB[294] WLB[293] WLB[292] WLB[291] WLB[290] WLB[289] WLB[288]
+WLB[287] WLB[286] WLB[285] WLB[284] WLB[283] WLB[282] WLB[281] WLB[280] WLB[279] WLB[278]
+WLB[277] WLB[276] WLB[275] WLB[274] WLB[273] WLB[272] WLB[271] WLB[270] WLB[269] WLB[268]
+WLB[267] WLB[266] WLB[265] WLB[264] WLB[263] WLB[262] WLB[261] WLB[260] WLB[259] WLB[258]
+WLB[257] WLB[256] S55NLLGDPH_X512Y8D16_BW_BITCELL64X8B
XI5 BLXA[7] BLXA[6] BLXA[5] BLXA[4] BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6]
+BLXB[5] BLXB[4] BLXB[3] BLXB[2] BLXB[1] BLXB[0] BLA[7] BLA[6] BLA[5] BLA[4]
+BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6] BLB[5] BLB[4] BLB[3] BLB[2]
+BLB[1] BLB[0] VDD VSS WLA[383] WLA[382] WLA[381] WLA[380] WLA[379] WLA[378]
+WLA[377] WLA[376] WLA[375] WLA[374] WLA[373] WLA[372] WLA[371] WLA[370] WLA[369] WLA[368]
+WLA[367] WLA[366] WLA[365] WLA[364] WLA[363] WLA[362] WLA[361] WLA[360] WLA[359] WLA[358]
+WLA[357] WLA[356] WLA[355] WLA[354] WLA[353] WLA[352] WLA[351] WLA[350] WLA[349] WLA[348]
+WLA[347] WLA[346] WLA[345] WLA[344] WLA[343] WLA[342] WLA[341] WLA[340] WLA[339] WLA[338]
+WLA[337] WLA[336] WLA[335] WLA[334] WLA[333] WLA[332] WLA[331] WLA[330] WLA[329] WLA[328]
+WLA[327] WLA[326] WLA[325] WLA[324] WLA[323] WLA[322] WLA[321] WLA[320] WLB[383] WLB[382]
+WLB[381] WLB[380] WLB[379] WLB[378] WLB[377] WLB[376] WLB[375] WLB[374] WLB[373] WLB[372]
+WLB[371] WLB[370] WLB[369] WLB[368] WLB[367] WLB[366] WLB[365] WLB[364] WLB[363] WLB[362]
+WLB[361] WLB[360] WLB[359] WLB[358] WLB[357] WLB[356] WLB[355] WLB[354] WLB[353] WLB[352]
+WLB[351] WLB[350] WLB[349] WLB[348] WLB[347] WLB[346] WLB[345] WLB[344] WLB[343] WLB[342]
+WLB[341] WLB[340] WLB[339] WLB[338] WLB[337] WLB[336] WLB[335] WLB[334] WLB[333] WLB[332]
+WLB[331] WLB[330] WLB[329] WLB[328] WLB[327] WLB[326] WLB[325] WLB[324] WLB[323] WLB[322]
+WLB[321] WLB[320] S55NLLGDPH_X512Y8D16_BW_BITCELL64X8A
XI6 BLXA[7] BLXA[6] BLXA[5] BLXA[4] BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6]
+BLXB[5] BLXB[4] BLXB[3] BLXB[2] BLXB[1] BLXB[0] BLA[7] BLA[6] BLA[5] BLA[4]
+BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6] BLB[5] BLB[4] BLB[3] BLB[2]
+BLB[1] BLB[0] VDD VSS WLA[447] WLA[446] WLA[445] WLA[444] WLA[443] WLA[442]
+WLA[441] WLA[440] WLA[439] WLA[438] WLA[437] WLA[436] WLA[435] WLA[434] WLA[433] WLA[432]
+WLA[431] WLA[430] WLA[429] WLA[428] WLA[427] WLA[426] WLA[425] WLA[424] WLA[423] WLA[422]
+WLA[421] WLA[420] WLA[419] WLA[418] WLA[417] WLA[416] WLA[415] WLA[414] WLA[413] WLA[412]
+WLA[411] WLA[410] WLA[409] WLA[408] WLA[407] WLA[406] WLA[405] WLA[404] WLA[403] WLA[402]
+WLA[401] WLA[400] WLA[399] WLA[398] WLA[397] WLA[396] WLA[395] WLA[394] WLA[393] WLA[392]
+WLA[391] WLA[390] WLA[389] WLA[388] WLA[387] WLA[386] WLA[385] WLA[384] WLB[447] WLB[446]
+WLB[445] WLB[444] WLB[443] WLB[442] WLB[441] WLB[440] WLB[439] WLB[438] WLB[437] WLB[436]
+WLB[435] WLB[434] WLB[433] WLB[432] WLB[431] WLB[430] WLB[429] WLB[428] WLB[427] WLB[426]
+WLB[425] WLB[424] WLB[423] WLB[422] WLB[421] WLB[420] WLB[419] WLB[418] WLB[417] WLB[416]
+WLB[415] WLB[414] WLB[413] WLB[412] WLB[411] WLB[410] WLB[409] WLB[408] WLB[407] WLB[406]
+WLB[405] WLB[404] WLB[403] WLB[402] WLB[401] WLB[400] WLB[399] WLB[398] WLB[397] WLB[396]
+WLB[395] WLB[394] WLB[393] WLB[392] WLB[391] WLB[390] WLB[389] WLB[388] WLB[387] WLB[386]
+WLB[385] WLB[384] S55NLLGDPH_X512Y8D16_BW_BITCELL64X8B
XI7 BLXA[7] BLXA[6] BLXA[5] BLXA[4] BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6]
+BLXB[5] BLXB[4] BLXB[3] BLXB[2] BLXB[1] BLXB[0] BLA[7] BLA[6] BLA[5] BLA[4]
+BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6] BLB[5] BLB[4] BLB[3] BLB[2]
+BLB[1] BLB[0] RDWLA[3] RDWLA[2] RDWLA[1] RDWLA[0] RDWLB[3] RDWLB[2] RDWLB[1] RDWLB[0]
+VDD VSS WLA[511] WLA[510] WLA[509] WLA[508] WLA[507] WLA[506] WLA[505] WLA[504]
+WLA[503] WLA[502] WLA[501] WLA[500] WLA[499] WLA[498] WLA[497] WLA[496] WLA[495] WLA[494]
+WLA[493] WLA[492] WLA[491] WLA[490] WLA[489] WLA[488] WLA[487] WLA[486] WLA[485] WLA[484]
+WLA[483] WLA[482] WLA[481] WLA[480] WLA[479] WLA[478] WLA[477] WLA[476] WLA[475] WLA[474]
+WLA[473] WLA[472] WLA[471] WLA[470] WLA[469] WLA[468] WLA[467] WLA[466] WLA[465] WLA[464]
+WLA[463] WLA[462] WLA[461] WLA[460] WLA[459] WLA[458] WLA[457] WLA[456] WLA[455] WLA[454]
+WLA[453] WLA[452] WLA[451] WLA[450] WLA[449] WLA[448] WLB[511] WLB[510] WLB[509] WLB[508]
+WLB[507] WLB[506] WLB[505] WLB[504] WLB[503] WLB[502] WLB[501] WLB[500] WLB[499] WLB[498]
+WLB[497] WLB[496] WLB[495] WLB[494] WLB[493] WLB[492] WLB[491] WLB[490] WLB[489] WLB[488]
+WLB[487] WLB[486] WLB[485] WLB[484] WLB[483] WLB[482] WLB[481] WLB[480] WLB[479] WLB[478]
+WLB[477] WLB[476] WLB[475] WLB[474] WLB[473] WLB[472] WLB[471] WLB[470] WLB[469] WLB[468]
+WLB[467] WLB[466] WLB[465] WLB[464] WLB[463] WLB[462] WLB[461] WLB[460] WLB[459] WLB[458]
+WLB[457] WLB[456] WLB[455] WLB[454] WLB[453] WLB[452] WLB[451] WLB[450] WLB[449] WLB[448] S55NLLGDPH_X512Y8D16_BW_BITCELL68X8A_NOMID_TOP
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    S55NLLGDPH_X512Y8D16_BW_YMX8SAWRA_B_BW
* View Name:    schematic
************************************************************************

.SUBCKT S55NLLGDPH_X512Y8D16_BW_YMX8SAWRA_B_BW BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] BWENA BWENB CLKA CLKB CLKXA CLKXB DATAA DATAB
+DOUTA DOUTB SACK1A SACK1B SACK4A SACK4B VDD VSS WEA WEB
+YXA[7] YXA[6] YXA[5] YXA[4] YXA[3] YXA[2] YXA[1] YXA[0] YXB[7] YXB[6]
+YXB[5] YXB[4] YXB[3] YXB[2] YXB[1] YXB[0]
M0 101 51 VSS VSS N12LL L=6E-08 W=1.2E-06
M1 VSS 109 108 VSS N12LL L=6E-08 W=1.5E-06
M2 104 101 VSS VSS N12LL L=6E-08 W=1.5E-06
M3 319 SACK4A 102 VSS N12LL L=6E-08 W=4E-07
M4 VSS SACK4A 103 VSS N12LL L=6E-08 W=4E-07
M5 104 3 BLXA[0] VSS N12LL L=6E-08 W=1.5E-06
M6 105 YXA[0] VSS VSS N12LL L=6E-08 W=4E-07
M7 VSS SACK1A 319 VSS N12LL L=6E-08 W=4E-07
M8 106 103 VSS VSS N12LL L=6E-08 W=8E-07
M9 BLA[0] 4 104 VSS N12LL L=6E-08 W=1.5E-06
M10 VSS 105 51 VSS N12LL L=6E-08 W=1.2E-06
M11 54 102 VSS VSS N12LL L=6E-08 W=5E-07
M12 58 107 VSS VSS N12LL L=6E-08 W=1.2E-06
M13 113 56 61 VSS N12LL L=1E-07 W=1.5E-06
M14 108 4 BLA[1] VSS N12LL L=6E-08 W=1.5E-06
M15 326 106 VSS VSS N12LL L=6E-08 W=1E-06
M16 113 116 326 VSS N12LL L=6E-08 W=1E-06
M17 VSS YXA[1] 107 VSS N12LL L=6E-08 W=4E-07
M18 61 56 113 VSS N12LL L=1E-07 W=1.5E-06
M19 BLXA[1] 3 108 VSS N12LL L=6E-08 W=1.5E-06
M20 327 56 110 VSS N12LL L=6E-08 W=1E-06
M21 VSS 110 DOUTA VSS N12LL L=6E-08 W=7.5E-07
M22 VSS 112 327 VSS N12LL L=6E-08 W=1E-06
M23 VSS 58 109 VSS N12LL L=6E-08 W=1.2E-06
M24 DOUTA 110 VSS VSS N12LL L=6E-08 W=7.5E-07
M25 334 110 VSS VSS N12LL L=6E-08 W=1E-06
M26 111 59 VSS VSS N12LL L=6E-08 W=1.2E-06
M27 118 120 VSS VSS N12LL L=6E-08 W=1.5E-06
M28 VSS 111 114 VSS N12LL L=6E-08 W=1.5E-06
M29 112 61 334 VSS N12LL L=6E-08 W=1E-06
M30 113 61 56 VSS N12LL L=1E-07 W=1.5E-06
M31 114 5 BLB[1] VSS N12LL L=6E-08 W=1.5E-06
M32 115 YXB[1] VSS VSS N12LL L=6E-08 W=4E-07
M33 BLXB[1] 6 114 VSS N12LL L=6E-08 W=1.5E-06
M34 56 61 113 VSS N12LL L=1E-07 W=1.5E-06
M35 VSS 115 59 VSS N12LL L=6E-08 W=1.2E-06
M36 63 117 VSS VSS N12LL L=6E-08 W=1.2E-06
M37 118 6 BLXB[0] VSS N12LL L=6E-08 W=1.5E-06
M38 VSS 119 116 VSS N12LL L=6E-08 W=5E-07
M39 VSS YXB[0] 117 VSS N12LL L=6E-08 W=4E-07
M40 BLB[0] 5 118 VSS N12LL L=6E-08 W=1.5E-06
M41 119 SACK1A VSS VSS N12LL L=6E-08 W=4E-07
M42 VSS 63 120 VSS N12LL L=6E-08 W=1.2E-06
M43 121 64 VSS VSS N12LL L=6E-08 W=1.2E-06
M44 VSS 132 131 VSS N12LL L=6E-08 W=1.5E-06
M45 123 121 VSS VSS N12LL L=6E-08 W=1.5E-06
M46 123 5 BLB[2] VSS N12LL L=6E-08 W=1.5E-06
M47 127 CLKXA 66 VSS N12LL L=6E-08 W=7E-07
M48 124 YXB[2] VSS VSS N12LL L=6E-08 W=4E-07
M49 VSS 144 122 VSS N12LL L=6E-08 W=4E-07
M50 348 122 VSS VSS N12LL L=6E-08 W=1E-06
M51 BLXB[2] 6 123 VSS N12LL L=6E-08 W=1.5E-06
M52 VSS 144 127 VSS N12LL L=6E-07 W=1.2E-07
M53 130 137 348 VSS N12LL L=6E-08 W=1E-06
M54 VSS 124 64 VSS N12LL L=6E-08 W=1.2E-06
M55 137 146 VSS VSS N12LL L=6E-08 W=5E-07
M56 70 129 VSS VSS N12LL L=6E-08 W=1.2E-06
M57 131 6 BLXB[3] VSS N12LL L=6E-08 W=1.5E-06
M58 VSS DATAA 126 VSS N12LL L=6E-08 W=4E-07
M59 128 126 VSS VSS N12LL L=3E-07 W=4E-07
M60 VSS 128 125 VSS N12LL L=2E-07 W=4E-07
M61 66 125 VSS VSS N12LL L=6E-08 W=3.5E-07
M62 VSS 125 66 VSS N12LL L=6E-08 W=3.5E-07
M63 VSS VSS DATAA VSS N12LL L=6E-08 W=2E-07
M64 VSS YXB[3] 129 VSS N12LL L=6E-08 W=4E-07
M65 BLB[3] 5 131 VSS N12LL L=6E-08 W=1.5E-06
M66 3 130 VSS VSS N12LL L=6E-08 W=1E-06
M67 144 127 VSS VSS N12LL L=6E-08 W=5E-07
M68 VSS 130 3 VSS N12LL L=6E-08 W=1E-06
M69 VSS 70 132 VSS N12LL L=6E-08 W=1.2E-06
M70 4 141 VSS VSS N12LL L=6E-08 W=1E-06
M71 133 71 VSS VSS N12LL L=6E-08 W=1.2E-06
M72 145 147 VSS VSS N12LL L=6E-08 W=1.5E-06
M73 VSS 133 134 VSS N12LL L=6E-08 W=1.5E-06
M74 VSS 138 143 VSS N12LL L=6E-08 W=4E-07
M75 VSS VSS BWENA VSS N12LL L=6E-08 W=2E-07
M76 VSS BWENA 136 VSS N12LL L=6E-08 W=4E-07
M77 140 136 VSS VSS N12LL L=3E-07 W=4E-07
M78 VSS 140 139 VSS N12LL L=2E-07 W=4E-07
M79 73 139 VSS VSS N12LL L=6E-08 W=3.5E-07
M80 VSS 139 73 VSS N12LL L=6E-08 W=3.5E-07
M81 VSS 141 4 VSS N12LL L=6E-08 W=1E-06
M82 134 3 BLXA[3] VSS N12LL L=6E-08 W=1.5E-06
M83 135 YXA[3] VSS VSS N12LL L=6E-08 W=4E-07
M84 138 143 VSS VSS N12LL L=6E-07 W=1.2E-07
M85 BLA[3] 4 134 VSS N12LL L=6E-08 W=1.5E-06
M86 VSS 135 71 VSS N12LL L=6E-08 W=1.2E-06
M87 75 142 VSS VSS N12LL L=6E-08 W=1.2E-06
M88 367 137 141 VSS N12LL L=6E-08 W=1E-06
M89 145 4 BLA[2] VSS N12LL L=6E-08 W=1.5E-06
M90 VSS 144 367 VSS N12LL L=6E-08 W=1E-06
M91 VSS YXA[2] 142 VSS N12LL L=6E-08 W=4E-07
M92 73 CLKXA 138 VSS N12LL L=6E-08 W=7E-07
M93 BLXA[2] 3 145 VSS N12LL L=6E-08 W=1.5E-06
M94 368 143 146 VSS N12LL L=6E-08 W=4E-07
M95 VSS WEA 368 VSS N12LL L=6E-08 W=4E-07
M96 VSS 75 147 VSS N12LL L=6E-08 W=1.2E-06
M97 375 WEB VSS VSS N12LL L=6E-08 W=4E-07
M98 148 76 VSS VSS N12LL L=6E-08 W=1.2E-06
M99 VSS 160 158 VSS N12LL L=6E-08 W=1.5E-06
M100 149 148 VSS VSS N12LL L=6E-08 W=1.5E-06
M101 150 159 375 VSS N12LL L=6E-08 W=4E-07
M102 149 3 BLXA[4] VSS N12LL L=6E-08 W=1.5E-06
M103 154 CLKXB 77 VSS N12LL L=6E-08 W=7E-07
M104 151 YXA[4] VSS VSS N12LL L=6E-08 W=4E-07
M105 376 172 VSS VSS N12LL L=6E-08 W=1E-06
M106 BLA[4] 4 149 VSS N12LL L=6E-08 W=1.5E-06
M107 VSS 159 154 VSS N12LL L=6E-07 W=1.2E-07
M108 157 165 376 VSS N12LL L=6E-08 W=1E-06
M109 VSS 151 76 VSS N12LL L=6E-08 W=1.2E-06
M110 82 156 VSS VSS N12LL L=6E-08 W=1.2E-06
M111 158 4 BLA[5] VSS N12LL L=6E-08 W=1.5E-06
M112 VSS BWENB 153 VSS N12LL L=6E-08 W=4E-07
M113 155 153 VSS VSS N12LL L=3E-07 W=4E-07
M114 VSS 155 152 VSS N12LL L=2E-07 W=4E-07
M115 77 152 VSS VSS N12LL L=6E-08 W=3.5E-07
M116 VSS 152 77 VSS N12LL L=6E-08 W=3.5E-07
M117 VSS VSS BWENB VSS N12LL L=6E-08 W=2E-07
M118 VSS YXA[5] 156 VSS N12LL L=6E-08 W=4E-07
M119 BLXA[5] 3 158 VSS N12LL L=6E-08 W=1.5E-06
M120 5 157 VSS VSS N12LL L=6E-08 W=1E-06
M121 159 154 VSS VSS N12LL L=6E-08 W=4E-07
M122 VSS 157 5 VSS N12LL L=6E-08 W=1E-06
M123 VSS 82 160 VSS N12LL L=6E-08 W=1.2E-06
M124 6 169 VSS VSS N12LL L=6E-08 W=1E-06
M125 161 83 VSS VSS N12LL L=6E-08 W=1.2E-06
M126 171 174 VSS VSS N12LL L=6E-08 W=1.5E-06
M127 VSS 161 162 VSS N12LL L=6E-08 W=1.5E-06
M128 VSS 166 172 VSS N12LL L=6E-08 W=5E-07
M129 VSS VSS DATAB VSS N12LL L=6E-08 W=2E-07
M130 VSS DATAB 164 VSS N12LL L=6E-08 W=4E-07
M131 168 164 VSS VSS N12LL L=3E-07 W=4E-07
M132 VSS 168 167 VSS N12LL L=2E-07 W=4E-07
M133 86 167 VSS VSS N12LL L=6E-08 W=3.5E-07
M134 VSS 167 86 VSS N12LL L=6E-08 W=3.5E-07
M135 VSS 169 6 VSS N12LL L=6E-08 W=1E-06
M136 162 5 BLB[5] VSS N12LL L=6E-08 W=1.5E-06
M137 163 YXB[5] VSS VSS N12LL L=6E-08 W=4E-07
M138 166 172 VSS VSS N12LL L=6E-07 W=1.2E-07
M139 BLXB[5] 6 162 VSS N12LL L=6E-08 W=1.5E-06
M140 VSS 163 83 VSS N12LL L=6E-08 W=1.2E-06
M141 VSS 150 165 VSS N12LL L=6E-08 W=5E-07
M142 87 170 VSS VSS N12LL L=6E-08 W=1.2E-06
M143 395 165 169 VSS N12LL L=6E-08 W=1E-06
M144 171 6 BLXB[4] VSS N12LL L=6E-08 W=1.5E-06
M145 173 172 VSS VSS N12LL L=6E-08 W=4E-07
M146 VSS 173 395 VSS N12LL L=6E-08 W=1E-06
M147 VSS YXB[4] 170 VSS N12LL L=6E-08 W=4E-07
M148 86 CLKXB 166 VSS N12LL L=6E-08 W=7E-07
M149 BLB[4] 5 171 VSS N12LL L=6E-08 W=1.5E-06
M150 VSS 87 174 VSS N12LL L=6E-08 W=1.2E-06
M151 175 88 VSS VSS N12LL L=6E-08 W=1.2E-06
M152 VSS 182 181 VSS N12LL L=6E-08 W=1.5E-06
M153 177 175 VSS VSS N12LL L=6E-08 W=1.5E-06
M154 VSS SACK1B 176 VSS N12LL L=6E-08 W=4E-07
M155 177 5 BLB[6] VSS N12LL L=6E-08 W=1.5E-06
M156 178 YXB[6] VSS VSS N12LL L=6E-08 W=4E-07
M157 179 176 VSS VSS N12LL L=6E-08 W=5E-07
M158 BLXB[6] 6 177 VSS N12LL L=6E-08 W=1.5E-06
M159 VSS 178 88 VSS N12LL L=6E-08 W=1.2E-06
M160 94 180 VSS VSS N12LL L=6E-08 W=1.2E-06
M161 186 92 96 VSS N12LL L=1E-07 W=1.5E-06
M162 181 6 BLXB[7] VSS N12LL L=6E-08 W=1.5E-06
M163 409 189 VSS VSS N12LL L=6E-08 W=1E-06
M164 186 179 409 VSS N12LL L=6E-08 W=1E-06
M165 VSS YXB[7] 180 VSS N12LL L=6E-08 W=4E-07
M166 96 92 186 VSS N12LL L=1E-07 W=1.5E-06
M167 BLB[7] 5 181 VSS N12LL L=6E-08 W=1.5E-06
M168 410 92 183 VSS N12LL L=6E-08 W=1E-06
M169 VSS 185 DOUTB VSS N12LL L=6E-08 W=7.5E-07
M170 VSS 185 410 VSS N12LL L=6E-08 W=1E-06
M171 VSS 94 182 VSS N12LL L=6E-08 W=1.2E-06
M172 DOUTB 185 VSS VSS N12LL L=6E-08 W=7.5E-07
M173 417 183 VSS VSS N12LL L=6E-08 W=1E-06
M174 184 95 VSS VSS N12LL L=6E-08 W=1.2E-06
M175 191 194 VSS VSS N12LL L=6E-08 W=1.5E-06
M176 VSS 184 187 VSS N12LL L=6E-08 W=1.5E-06
M177 185 96 417 VSS N12LL L=6E-08 W=1E-06
M178 186 96 92 VSS N12LL L=1E-07 W=1.5E-06
M179 187 3 BLXA[7] VSS N12LL L=6E-08 W=1.5E-06
M180 188 YXA[7] VSS VSS N12LL L=6E-08 W=4E-07
M181 BLA[7] 4 187 VSS N12LL L=6E-08 W=1.5E-06
M182 92 96 186 VSS N12LL L=1E-07 W=1.5E-06
M183 VSS 188 95 VSS N12LL L=6E-08 W=1.2E-06
M184 VSS 193 97 VSS N12LL L=6E-08 W=5E-07
M185 100 190 VSS VSS N12LL L=6E-08 W=1.2E-06
M186 191 4 BLA[6] VSS N12LL L=6E-08 W=1.5E-06
M187 VSS 192 189 VSS N12LL L=6E-08 W=8E-07
M188 424 SACK1B VSS VSS N12LL L=6E-08 W=4E-07
M189 VSS YXA[6] 190 VSS N12LL L=6E-08 W=4E-07
M190 BLXA[6] 3 191 VSS N12LL L=6E-08 W=1.5E-06
M191 192 SACK4B VSS VSS N12LL L=6E-08 W=4E-07
M192 193 SACK4B 424 VSS N12LL L=6E-08 W=4E-07
M193 VSS 100 194 VSS N12LL L=6E-08 W=1.2E-06
M194 BLXA[0] 101 VDD VDD P12LL L=6E-08 W=2E-06
M195 101 51 VDD VDD P12LL L=6E-08 W=1.2E-06
M196 102 SACK4A VDD VDD P12LL L=6E-08 W=4E-07
M197 VDD SACK4A 103 VDD P12LL L=6E-08 W=8E-07
M198 BLA[0] 101 BLXA[0] VDD P12LL L=6E-08 W=2E-06
M199 105 YXA[0] VDD VDD P12LL L=6E-08 W=4E-07
M200 BLXA[0] 51 32 VDD P12LL L=6E-08 W=3E-07
M201 BLA[0] 51 50 VDD P12LL L=6E-08 W=3E-07
M202 VDD SACK1A 102 VDD P12LL L=6E-08 W=4E-07
M203 106 103 VDD VDD P12LL L=6E-08 W=1.6E-06
M204 VDD 101 BLA[0] VDD P12LL L=6E-08 W=2E-06
M205 32 51 BLXA[0] VDD P12LL L=6E-08 W=3E-07
M206 50 51 BLA[0] VDD P12LL L=6E-08 W=3E-07
M207 VDD 105 51 VDD P12LL L=6E-08 W=1.2E-06
M208 54 102 VDD VDD P12LL L=6E-08 W=1E-06
M209 56 54 50 VDD P12LL L=6E-08 W=7E-07
M210 50 54 56 VDD P12LL L=6E-08 W=7E-07
M211 BLXA[1] 58 32 VDD P12LL L=6E-08 W=3E-07
M212 BLA[1] 58 50 VDD P12LL L=6E-08 W=3E-07
M213 58 107 VDD VDD P12LL L=6E-08 W=1.2E-06
M214 VDD 56 61 VDD P12LL L=1E-07 W=4E-07
M215 VDD 106 50 VDD P12LL L=6E-08 W=5E-07
M216 50 106 VDD VDD P12LL L=6E-08 W=5E-07
M217 32 106 50 VDD P12LL L=6E-08 W=5E-07
M218 BLA[1] 109 VDD VDD P12LL L=6E-08 W=2E-06
M219 32 58 BLXA[1] VDD P12LL L=6E-08 W=3E-07
M220 50 58 BLA[1] VDD P12LL L=6E-08 W=3E-07
M221 61 56 VDD VDD P12LL L=1E-07 W=4E-07
M222 VDD YXA[1] 107 VDD P12LL L=6E-08 W=4E-07
M223 110 56 VDD VDD P12LL L=6E-08 W=1E-06
M224 BLXA[1] 109 BLA[1] VDD P12LL L=6E-08 W=2E-06
M225 VDD 110 DOUTA VDD P12LL L=6E-08 W=1.5E-06
M226 VDD 112 110 VDD P12LL L=6E-08 W=1E-06
M227 VDD 58 109 VDD P12LL L=6E-08 W=1.2E-06
M228 VDD 109 BLXA[1] VDD P12LL L=6E-08 W=2E-06
M229 BLB[1] 111 VDD VDD P12LL L=6E-08 W=2E-06
M230 DOUTA 110 VDD VDD P12LL L=6E-08 W=1.5E-06
M231 112 110 VDD VDD P12LL L=6E-08 W=1E-06
M232 111 59 VDD VDD P12LL L=6E-08 W=1.2E-06
M233 61 54 32 VDD P12LL L=6E-08 W=7E-07
M234 32 54 61 VDD P12LL L=6E-08 W=7E-07
M235 VDD 106 32 VDD P12LL L=6E-08 W=5E-07
M236 32 106 VDD VDD P12LL L=6E-08 W=5E-07
M237 50 106 32 VDD P12LL L=6E-08 W=5E-07
M238 BLXB[1] 111 BLB[1] VDD P12LL L=6E-08 W=2E-06
M239 VDD 61 112 VDD P12LL L=6E-08 W=1E-06
M240 VDD 61 56 VDD P12LL L=1E-07 W=4E-07
M241 115 YXB[1] VDD VDD P12LL L=6E-08 W=4E-07
M242 BLB[1] 59 46 VDD P12LL L=6E-08 W=3E-07
M243 BLXB[1] 59 48 VDD P12LL L=6E-08 W=3E-07
M244 VDD 111 BLXB[1] VDD P12LL L=6E-08 W=2E-06
M245 56 61 VDD VDD P12LL L=1E-07 W=4E-07
M246 46 59 BLB[1] VDD P12LL L=6E-08 W=3E-07
M247 48 59 BLXB[1] VDD P12LL L=6E-08 W=3E-07
M248 VDD 115 59 VDD P12LL L=6E-08 W=1.2E-06
M249 BLB[0] 63 46 VDD P12LL L=6E-08 W=3E-07
M250 BLXB[0] 63 48 VDD P12LL L=6E-08 W=3E-07
M251 63 117 VDD VDD P12LL L=6E-08 W=1.2E-06
M252 BLXB[0] 120 VDD VDD P12LL L=6E-08 W=2E-06
M253 VDD 119 116 VDD P12LL L=6E-08 W=1E-06
M254 46 63 BLB[0] VDD P12LL L=6E-08 W=3E-07
M255 48 63 BLXB[0] VDD P12LL L=6E-08 W=3E-07
M256 VDD YXB[0] 117 VDD P12LL L=6E-08 W=4E-07
M257 BLB[0] 120 BLXB[0] VDD P12LL L=6E-08 W=2E-06
M258 119 SACK1A VDD VDD P12LL L=6E-08 W=4E-07
M259 VDD 63 120 VDD P12LL L=6E-08 W=1.2E-06
M260 VDD 120 BLB[0] VDD P12LL L=6E-08 W=2E-06
M261 BLB[2] 121 VDD VDD P12LL L=6E-08 W=2E-06
M262 121 64 VDD VDD P12LL L=6E-08 W=1.2E-06
M263 VDD VDD DATAA VDD P12LL L=6E-08 W=2E-07
M264 VDD DATAA 126 VDD P12LL L=6E-08 W=4E-07
M265 128 126 VDD VDD P12LL L=3E-07 W=4E-07
M266 VDD 128 125 VDD P12LL L=2E-07 W=4E-07
M267 66 125 VDD VDD P12LL L=6E-08 W=3.5E-07
M268 VDD 125 66 VDD P12LL L=6E-08 W=3.5E-07
M269 BLXB[2] 121 BLB[2] VDD P12LL L=6E-08 W=2E-06
M270 124 YXB[2] VDD VDD P12LL L=6E-08 W=4E-07
M271 VDD 144 122 VDD P12LL L=6E-08 W=4E-07
M272 130 122 VDD VDD P12LL L=6E-08 W=8E-07
M273 BLB[2] 64 46 VDD P12LL L=6E-08 W=3E-07
M274 BLXB[2] 64 48 VDD P12LL L=6E-08 W=3E-07
M275 VDD 121 BLXB[2] VDD P12LL L=6E-08 W=2E-06
M276 127 CLKA 66 VDD P12LL L=6E-08 W=7E-07
M277 VDD 137 130 VDD P12LL L=6E-08 W=8E-07
M278 46 64 BLB[2] VDD P12LL L=6E-08 W=3E-07
M279 48 64 BLXB[2] VDD P12LL L=6E-08 W=3E-07
M280 VDD 124 64 VDD P12LL L=6E-08 W=1.2E-06
M281 137 146 VDD VDD P12LL L=6E-08 W=1E-06
M282 VDD 144 127 VDD P12LL L=3E-07 W=1.2E-07
M283 BLB[3] 70 46 VDD P12LL L=6E-08 W=3E-07
M284 BLXB[3] 70 48 VDD P12LL L=6E-08 W=3E-07
M285 70 129 VDD VDD P12LL L=6E-08 W=1.2E-06
M286 BLXB[3] 132 VDD VDD P12LL L=6E-08 W=2E-06
M287 46 70 BLB[3] VDD P12LL L=6E-08 W=3E-07
M288 48 70 BLXB[3] VDD P12LL L=6E-08 W=3E-07
M289 VDD YXB[3] 129 VDD P12LL L=6E-08 W=4E-07
M290 3 130 VDD VDD P12LL L=6E-08 W=2E-06
M291 BLB[3] 132 BLXB[3] VDD P12LL L=6E-08 W=2E-06
M292 144 127 VDD VDD P12LL L=6E-08 W=8E-07
M293 VDD 130 3 VDD P12LL L=6E-08 W=2E-06
M294 VDD 70 132 VDD P12LL L=6E-08 W=1.2E-06
M295 VDD 132 BLB[3] VDD P12LL L=6E-08 W=2E-06
M296 BLXA[3] 133 VDD VDD P12LL L=6E-08 W=2E-06
M297 4 141 VDD VDD P12LL L=6E-08 W=2E-06
M298 133 71 VDD VDD P12LL L=6E-08 W=1.2E-06
M299 VDD 138 143 VDD P12LL L=6E-08 W=4E-07
M300 BLA[3] 133 BLXA[3] VDD P12LL L=6E-08 W=2E-06
M301 VDD 141 4 VDD P12LL L=6E-08 W=2E-06
M302 135 YXA[3] VDD VDD P12LL L=6E-08 W=4E-07
M303 BLXA[3] 71 32 VDD P12LL L=6E-08 W=3E-07
M304 BLA[3] 71 50 VDD P12LL L=6E-08 W=3E-07
M305 138 143 VDD VDD P12LL L=3E-07 W=1.2E-07
M306 VDD 133 BLA[3] VDD P12LL L=6E-08 W=2E-06
M307 32 71 BLXA[3] VDD P12LL L=6E-08 W=3E-07
M308 50 71 BLA[3] VDD P12LL L=6E-08 W=3E-07
M309 VDD 135 71 VDD P12LL L=6E-08 W=1.2E-06
M310 BLXA[2] 75 32 VDD P12LL L=6E-08 W=3E-07
M311 BLA[2] 75 50 VDD P12LL L=6E-08 W=3E-07
M312 75 142 VDD VDD P12LL L=6E-08 W=1.2E-06
M313 141 137 VDD VDD P12LL L=6E-08 W=8E-07
M314 73 CLKA 138 VDD P12LL L=6E-08 W=7E-07
M315 VDD BWENA 136 VDD P12LL L=6E-08 W=4E-07
M316 140 136 VDD VDD P12LL L=3E-07 W=4E-07
M317 VDD 140 139 VDD P12LL L=2E-07 W=4E-07
M318 73 139 VDD VDD P12LL L=6E-08 W=3.5E-07
M319 VDD 139 73 VDD P12LL L=6E-08 W=3.5E-07
M320 BLA[2] 147 VDD VDD P12LL L=6E-08 W=2E-06
M321 VDD 143 146 VDD P12LL L=6E-08 W=4E-07
M322 32 75 BLXA[2] VDD P12LL L=6E-08 W=3E-07
M323 50 75 BLA[2] VDD P12LL L=6E-08 W=3E-07
M324 VDD 144 141 VDD P12LL L=6E-08 W=8E-07
M325 VDD VDD BWENA VDD P12LL L=6E-08 W=2E-07
M326 VDD YXA[2] 142 VDD P12LL L=6E-08 W=4E-07
M327 BLXA[2] 147 BLA[2] VDD P12LL L=6E-08 W=2E-06
M328 146 WEA VDD VDD P12LL L=6E-08 W=4E-07
M329 VDD 75 147 VDD P12LL L=6E-08 W=1.2E-06
M330 VDD 147 BLXA[2] VDD P12LL L=6E-08 W=2E-06
M331 BLXA[4] 148 VDD VDD P12LL L=6E-08 W=2E-06
M332 148 76 VDD VDD P12LL L=6E-08 W=1.2E-06
M333 VDD WEB 150 VDD P12LL L=6E-08 W=4E-07
M334 VDD VDD BWENB VDD P12LL L=6E-08 W=2E-07
M335 VDD BWENB 153 VDD P12LL L=6E-08 W=4E-07
M336 155 153 VDD VDD P12LL L=3E-07 W=4E-07
M337 VDD 155 152 VDD P12LL L=2E-07 W=4E-07
M338 77 152 VDD VDD P12LL L=6E-08 W=3.5E-07
M339 VDD 152 77 VDD P12LL L=6E-08 W=3.5E-07
M340 BLA[4] 148 BLXA[4] VDD P12LL L=6E-08 W=2E-06
M341 151 YXA[4] VDD VDD P12LL L=6E-08 W=4E-07
M342 157 172 VDD VDD P12LL L=6E-08 W=8E-07
M343 BLXA[4] 76 32 VDD P12LL L=6E-08 W=3E-07
M344 BLA[4] 76 50 VDD P12LL L=6E-08 W=3E-07
M345 150 159 VDD VDD P12LL L=6E-08 W=4E-07
M346 VDD 148 BLA[4] VDD P12LL L=6E-08 W=2E-06
M347 154 CLKB 77 VDD P12LL L=6E-08 W=7E-07
M348 VDD 165 157 VDD P12LL L=6E-08 W=8E-07
M349 32 76 BLXA[4] VDD P12LL L=6E-08 W=3E-07
M350 50 76 BLA[4] VDD P12LL L=6E-08 W=3E-07
M351 VDD 151 76 VDD P12LL L=6E-08 W=1.2E-06
M352 VDD 159 154 VDD P12LL L=3E-07 W=1.2E-07
M353 BLXA[5] 82 32 VDD P12LL L=6E-08 W=3E-07
M354 BLA[5] 82 50 VDD P12LL L=6E-08 W=3E-07
M355 82 156 VDD VDD P12LL L=6E-08 W=1.2E-06
M356 BLA[5] 160 VDD VDD P12LL L=6E-08 W=2E-06
M357 32 82 BLXA[5] VDD P12LL L=6E-08 W=3E-07
M358 50 82 BLA[5] VDD P12LL L=6E-08 W=3E-07
M359 VDD YXA[5] 156 VDD P12LL L=6E-08 W=4E-07
M360 5 157 VDD VDD P12LL L=6E-08 W=2E-06
M361 BLXA[5] 160 BLA[5] VDD P12LL L=6E-08 W=2E-06
M362 159 154 VDD VDD P12LL L=6E-08 W=4E-07
M363 VDD 157 5 VDD P12LL L=6E-08 W=2E-06
M364 VDD 82 160 VDD P12LL L=6E-08 W=1.2E-06
M365 VDD 160 BLXA[5] VDD P12LL L=6E-08 W=2E-06
M366 BLB[5] 161 VDD VDD P12LL L=6E-08 W=2E-06
M367 6 169 VDD VDD P12LL L=6E-08 W=2E-06
M368 161 83 VDD VDD P12LL L=6E-08 W=1.2E-06
M369 VDD 166 172 VDD P12LL L=6E-08 W=8E-07
M370 BLXB[5] 161 BLB[5] VDD P12LL L=6E-08 W=2E-06
M371 VDD 169 6 VDD P12LL L=6E-08 W=2E-06
M372 163 YXB[5] VDD VDD P12LL L=6E-08 W=4E-07
M373 BLB[5] 83 46 VDD P12LL L=6E-08 W=3E-07
M374 BLXB[5] 83 48 VDD P12LL L=6E-08 W=3E-07
M375 166 172 VDD VDD P12LL L=3E-07 W=1.2E-07
M376 VDD 161 BLXB[5] VDD P12LL L=6E-08 W=2E-06
M377 46 83 BLB[5] VDD P12LL L=6E-08 W=3E-07
M378 48 83 BLXB[5] VDD P12LL L=6E-08 W=3E-07
M379 VDD 163 83 VDD P12LL L=6E-08 W=1.2E-06
M380 VDD 150 165 VDD P12LL L=6E-08 W=1E-06
M381 BLB[4] 87 46 VDD P12LL L=6E-08 W=3E-07
M382 BLXB[4] 87 48 VDD P12LL L=6E-08 W=3E-07
M383 87 170 VDD VDD P12LL L=6E-08 W=1.2E-06
M384 169 165 VDD VDD P12LL L=6E-08 W=8E-07
M385 86 CLKB 166 VDD P12LL L=6E-08 W=7E-07
M386 VDD DATAB 164 VDD P12LL L=6E-08 W=4E-07
M387 168 164 VDD VDD P12LL L=3E-07 W=4E-07
M388 VDD 168 167 VDD P12LL L=2E-07 W=4E-07
M389 86 167 VDD VDD P12LL L=6E-08 W=3.5E-07
M390 VDD 167 86 VDD P12LL L=6E-08 W=3.5E-07
M391 BLXB[4] 174 VDD VDD P12LL L=6E-08 W=2E-06
M392 46 87 BLB[4] VDD P12LL L=6E-08 W=3E-07
M393 48 87 BLXB[4] VDD P12LL L=6E-08 W=3E-07
M394 173 172 VDD VDD P12LL L=6E-08 W=4E-07
M395 VDD 173 169 VDD P12LL L=6E-08 W=8E-07
M396 VDD VDD DATAB VDD P12LL L=6E-08 W=2E-07
M397 VDD YXB[4] 170 VDD P12LL L=6E-08 W=4E-07
M398 BLB[4] 174 BLXB[4] VDD P12LL L=6E-08 W=2E-06
M399 VDD 87 174 VDD P12LL L=6E-08 W=1.2E-06
M400 VDD 174 BLB[4] VDD P12LL L=6E-08 W=2E-06
M401 BLB[6] 175 VDD VDD P12LL L=6E-08 W=2E-06
M402 175 88 VDD VDD P12LL L=6E-08 W=1.2E-06
M403 VDD SACK1B 176 VDD P12LL L=6E-08 W=4E-07
M404 BLXB[6] 175 BLB[6] VDD P12LL L=6E-08 W=2E-06
M405 178 YXB[6] VDD VDD P12LL L=6E-08 W=4E-07
M406 BLB[6] 88 46 VDD P12LL L=6E-08 W=3E-07
M407 BLXB[6] 88 48 VDD P12LL L=6E-08 W=3E-07
M408 179 176 VDD VDD P12LL L=6E-08 W=1E-06
M409 VDD 175 BLXB[6] VDD P12LL L=6E-08 W=2E-06
M410 46 88 BLB[6] VDD P12LL L=6E-08 W=3E-07
M411 48 88 BLXB[6] VDD P12LL L=6E-08 W=3E-07
M412 VDD 178 88 VDD P12LL L=6E-08 W=1.2E-06
M413 92 97 48 VDD P12LL L=6E-08 W=7E-07
M414 48 97 92 VDD P12LL L=6E-08 W=7E-07
M415 BLB[7] 94 46 VDD P12LL L=6E-08 W=3E-07
M416 BLXB[7] 94 48 VDD P12LL L=6E-08 W=3E-07
M417 94 180 VDD VDD P12LL L=6E-08 W=1.2E-06
M418 VDD 92 96 VDD P12LL L=1E-07 W=4E-07
M419 VDD 189 48 VDD P12LL L=6E-08 W=5E-07
M420 48 189 VDD VDD P12LL L=6E-08 W=5E-07
M421 46 189 48 VDD P12LL L=6E-08 W=5E-07
M422 BLXB[7] 182 VDD VDD P12LL L=6E-08 W=2E-06
M423 46 94 BLB[7] VDD P12LL L=6E-08 W=3E-07
M424 48 94 BLXB[7] VDD P12LL L=6E-08 W=3E-07
M425 96 92 VDD VDD P12LL L=1E-07 W=4E-07
M426 VDD YXB[7] 180 VDD P12LL L=6E-08 W=4E-07
M427 183 92 VDD VDD P12LL L=6E-08 W=1E-06
M428 BLB[7] 182 BLXB[7] VDD P12LL L=6E-08 W=2E-06
M429 VDD 185 DOUTB VDD P12LL L=6E-08 W=1.5E-06
M430 VDD 185 183 VDD P12LL L=6E-08 W=1E-06
M431 VDD 94 182 VDD P12LL L=6E-08 W=1.2E-06
M432 VDD 182 BLB[7] VDD P12LL L=6E-08 W=2E-06
M433 BLXA[7] 184 VDD VDD P12LL L=6E-08 W=2E-06
M434 DOUTB 185 VDD VDD P12LL L=6E-08 W=1.5E-06
M435 185 183 VDD VDD P12LL L=6E-08 W=1E-06
M436 184 95 VDD VDD P12LL L=6E-08 W=1.2E-06
M437 96 97 46 VDD P12LL L=6E-08 W=7E-07
M438 46 97 96 VDD P12LL L=6E-08 W=7E-07
M439 VDD 189 46 VDD P12LL L=6E-08 W=5E-07
M440 46 189 VDD VDD P12LL L=6E-08 W=5E-07
M441 48 189 46 VDD P12LL L=6E-08 W=5E-07
M442 BLA[7] 184 BLXA[7] VDD P12LL L=6E-08 W=2E-06
M443 VDD 96 185 VDD P12LL L=6E-08 W=1E-06
M444 VDD 96 92 VDD P12LL L=1E-07 W=4E-07
M445 188 YXA[7] VDD VDD P12LL L=6E-08 W=4E-07
M446 BLXA[7] 95 32 VDD P12LL L=6E-08 W=3E-07
M447 BLA[7] 95 50 VDD P12LL L=6E-08 W=3E-07
M448 VDD 184 BLA[7] VDD P12LL L=6E-08 W=2E-06
M449 92 96 VDD VDD P12LL L=1E-07 W=4E-07
M450 32 95 BLXA[7] VDD P12LL L=6E-08 W=3E-07
M451 50 95 BLA[7] VDD P12LL L=6E-08 W=3E-07
M452 VDD 188 95 VDD P12LL L=6E-08 W=1.2E-06
M453 VDD 193 97 VDD P12LL L=6E-08 W=1E-06
M454 BLXA[6] 100 32 VDD P12LL L=6E-08 W=3E-07
M455 BLA[6] 100 50 VDD P12LL L=6E-08 W=3E-07
M456 100 190 VDD VDD P12LL L=6E-08 W=1.2E-06
M457 BLA[6] 194 VDD VDD P12LL L=6E-08 W=2E-06
M458 VDD 192 189 VDD P12LL L=6E-08 W=1.6E-06
M459 193 SACK1B VDD VDD P12LL L=6E-08 W=4E-07
M460 32 100 BLXA[6] VDD P12LL L=6E-08 W=3E-07
M461 50 100 BLA[6] VDD P12LL L=6E-08 W=3E-07
M462 VDD YXA[6] 190 VDD P12LL L=6E-08 W=4E-07
M463 BLXA[6] 194 BLA[6] VDD P12LL L=6E-08 W=2E-06
M464 192 SACK4B VDD VDD P12LL L=6E-08 W=8E-07
M465 VDD SACK4B 193 VDD P12LL L=6E-08 W=4E-07
M466 VDD 100 194 VDD P12LL L=6E-08 W=1.2E-06
M467 VDD 194 BLXA[6] VDD P12LL L=6E-08 W=2E-06
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    S55NLLGDPH_X512Y8D16_BW_Y512X8CELL_BW
* View Name:    schematic
************************************************************************

.SUBCKT S55NLLGDPH_X512Y8D16_BW_Y512X8CELL_BW BWENA BWENB CLKA CLKB CLKXA CLKXB DATAA DATAB DOUTA DOUTB
+RDWLA[3] RDWLA[2] RDWLA[1] RDWLA[0] RDWLB[3] RDWLB[2] RDWLB[1] RDWLB[0] RWLA[0] RWLA[1]
+RWLB[0] RWLB[1] SACK1A SACK1B SACK4A SACK4B VDD VSS WEA WEB
+WLA[511] WLA[510] WLA[509] WLA[508] WLA[507] WLA[506] WLA[505] WLA[504] WLA[503] WLA[502]
+WLA[501] WLA[500] WLA[499] WLA[498] WLA[497] WLA[496] WLA[495] WLA[494] WLA[493] WLA[492]
+WLA[491] WLA[490] WLA[489] WLA[488] WLA[487] WLA[486] WLA[485] WLA[484] WLA[483] WLA[482]
+WLA[481] WLA[480] WLA[479] WLA[478] WLA[477] WLA[476] WLA[475] WLA[474] WLA[473] WLA[472]
+WLA[471] WLA[470] WLA[469] WLA[468] WLA[467] WLA[466] WLA[465] WLA[464] WLA[463] WLA[462]
+WLA[461] WLA[460] WLA[459] WLA[458] WLA[457] WLA[456] WLA[455] WLA[454] WLA[453] WLA[452]
+WLA[451] WLA[450] WLA[449] WLA[448] WLA[447] WLA[446] WLA[445] WLA[444] WLA[443] WLA[442]
+WLA[441] WLA[440] WLA[439] WLA[438] WLA[437] WLA[436] WLA[435] WLA[434] WLA[433] WLA[432]
+WLA[431] WLA[430] WLA[429] WLA[428] WLA[427] WLA[426] WLA[425] WLA[424] WLA[423] WLA[422]
+WLA[421] WLA[420] WLA[419] WLA[418] WLA[417] WLA[416] WLA[415] WLA[414] WLA[413] WLA[412]
+WLA[411] WLA[410] WLA[409] WLA[408] WLA[407] WLA[406] WLA[405] WLA[404] WLA[403] WLA[402]
+WLA[401] WLA[400] WLA[399] WLA[398] WLA[397] WLA[396] WLA[395] WLA[394] WLA[393] WLA[392]
+WLA[391] WLA[390] WLA[389] WLA[388] WLA[387] WLA[386] WLA[385] WLA[384] WLA[383] WLA[382]
+WLA[381] WLA[380] WLA[379] WLA[378] WLA[377] WLA[376] WLA[375] WLA[374] WLA[373] WLA[372]
+WLA[371] WLA[370] WLA[369] WLA[368] WLA[367] WLA[366] WLA[365] WLA[364] WLA[363] WLA[362]
+WLA[361] WLA[360] WLA[359] WLA[358] WLA[357] WLA[356] WLA[355] WLA[354] WLA[353] WLA[352]
+WLA[351] WLA[350] WLA[349] WLA[348] WLA[347] WLA[346] WLA[345] WLA[344] WLA[343] WLA[342]
+WLA[341] WLA[340] WLA[339] WLA[338] WLA[337] WLA[336] WLA[335] WLA[334] WLA[333] WLA[332]
+WLA[331] WLA[330] WLA[329] WLA[328] WLA[327] WLA[326] WLA[325] WLA[324] WLA[323] WLA[322]
+WLA[321] WLA[320] WLA[319] WLA[318] WLA[317] WLA[316] WLA[315] WLA[314] WLA[313] WLA[312]
+WLA[311] WLA[310] WLA[309] WLA[308] WLA[307] WLA[306] WLA[305] WLA[304] WLA[303] WLA[302]
+WLA[301] WLA[300] WLA[299] WLA[298] WLA[297] WLA[296] WLA[295] WLA[294] WLA[293] WLA[292]
+WLA[291] WLA[290] WLA[289] WLA[288] WLA[287] WLA[286] WLA[285] WLA[284] WLA[283] WLA[282]
+WLA[281] WLA[280] WLA[279] WLA[278] WLA[277] WLA[276] WLA[275] WLA[274] WLA[273] WLA[272]
+WLA[271] WLA[270] WLA[269] WLA[268] WLA[267] WLA[266] WLA[265] WLA[264] WLA[263] WLA[262]
+WLA[261] WLA[260] WLA[259] WLA[258] WLA[257] WLA[256] WLA[255] WLA[254] WLA[253] WLA[252]
+WLA[251] WLA[250] WLA[249] WLA[248] WLA[247] WLA[246] WLA[245] WLA[244] WLA[243] WLA[242]
+WLA[241] WLA[240] WLA[239] WLA[238] WLA[237] WLA[236] WLA[235] WLA[234] WLA[233] WLA[232]
+WLA[231] WLA[230] WLA[229] WLA[228] WLA[227] WLA[226] WLA[225] WLA[224] WLA[223] WLA[222]
+WLA[221] WLA[220] WLA[219] WLA[218] WLA[217] WLA[216] WLA[215] WLA[214] WLA[213] WLA[212]
+WLA[211] WLA[210] WLA[209] WLA[208] WLA[207] WLA[206] WLA[205] WLA[204] WLA[203] WLA[202]
+WLA[201] WLA[200] WLA[199] WLA[198] WLA[197] WLA[196] WLA[195] WLA[194] WLA[193] WLA[192]
+WLA[191] WLA[190] WLA[189] WLA[188] WLA[187] WLA[186] WLA[185] WLA[184] WLA[183] WLA[182]
+WLA[181] WLA[180] WLA[179] WLA[178] WLA[177] WLA[176] WLA[175] WLA[174] WLA[173] WLA[172]
+WLA[171] WLA[170] WLA[169] WLA[168] WLA[167] WLA[166] WLA[165] WLA[164] WLA[163] WLA[162]
+WLA[161] WLA[160] WLA[159] WLA[158] WLA[157] WLA[156] WLA[155] WLA[154] WLA[153] WLA[152]
+WLA[151] WLA[150] WLA[149] WLA[148] WLA[147] WLA[146] WLA[145] WLA[144] WLA[143] WLA[142]
+WLA[141] WLA[140] WLA[139] WLA[138] WLA[137] WLA[136] WLA[135] WLA[134] WLA[133] WLA[132]
+WLA[131] WLA[130] WLA[129] WLA[128] WLA[127] WLA[126] WLA[125] WLA[124] WLA[123] WLA[122]
+WLA[121] WLA[120] WLA[119] WLA[118] WLA[117] WLA[116] WLA[115] WLA[114] WLA[113] WLA[112]
+WLA[111] WLA[110] WLA[109] WLA[108] WLA[107] WLA[106] WLA[105] WLA[104] WLA[103] WLA[102]
+WLA[101] WLA[100] WLA[99] WLA[98] WLA[97] WLA[96] WLA[95] WLA[94] WLA[93] WLA[92]
+WLA[91] WLA[90] WLA[89] WLA[88] WLA[87] WLA[86] WLA[85] WLA[84] WLA[83] WLA[82]
+WLA[81] WLA[80] WLA[79] WLA[78] WLA[77] WLA[76] WLA[75] WLA[74] WLA[73] WLA[72]
+WLA[71] WLA[70] WLA[69] WLA[68] WLA[67] WLA[66] WLA[65] WLA[64] WLA[63] WLA[62]
+WLA[61] WLA[60] WLA[59] WLA[58] WLA[57] WLA[56] WLA[55] WLA[54] WLA[53] WLA[52]
+WLA[51] WLA[50] WLA[49] WLA[48] WLA[47] WLA[46] WLA[45] WLA[44] WLA[43] WLA[42]
+WLA[41] WLA[40] WLA[39] WLA[38] WLA[37] WLA[36] WLA[35] WLA[34] WLA[33] WLA[32]
+WLA[31] WLA[30] WLA[29] WLA[28] WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22]
+WLA[21] WLA[20] WLA[19] WLA[18] WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12]
+WLA[11] WLA[10] WLA[9] WLA[8] WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2]
+WLA[1] WLA[0] WLB[511] WLB[510] WLB[509] WLB[508] WLB[507] WLB[506] WLB[505] WLB[504]
+WLB[503] WLB[502] WLB[501] WLB[500] WLB[499] WLB[498] WLB[497] WLB[496] WLB[495] WLB[494]
+WLB[493] WLB[492] WLB[491] WLB[490] WLB[489] WLB[488] WLB[487] WLB[486] WLB[485] WLB[484]
+WLB[483] WLB[482] WLB[481] WLB[480] WLB[479] WLB[478] WLB[477] WLB[476] WLB[475] WLB[474]
+WLB[473] WLB[472] WLB[471] WLB[470] WLB[469] WLB[468] WLB[467] WLB[466] WLB[465] WLB[464]
+WLB[463] WLB[462] WLB[461] WLB[460] WLB[459] WLB[458] WLB[457] WLB[456] WLB[455] WLB[454]
+WLB[453] WLB[452] WLB[451] WLB[450] WLB[449] WLB[448] WLB[447] WLB[446] WLB[445] WLB[444]
+WLB[443] WLB[442] WLB[441] WLB[440] WLB[439] WLB[438] WLB[437] WLB[436] WLB[435] WLB[434]
+WLB[433] WLB[432] WLB[431] WLB[430] WLB[429] WLB[428] WLB[427] WLB[426] WLB[425] WLB[424]
+WLB[423] WLB[422] WLB[421] WLB[420] WLB[419] WLB[418] WLB[417] WLB[416] WLB[415] WLB[414]
+WLB[413] WLB[412] WLB[411] WLB[410] WLB[409] WLB[408] WLB[407] WLB[406] WLB[405] WLB[404]
+WLB[403] WLB[402] WLB[401] WLB[400] WLB[399] WLB[398] WLB[397] WLB[396] WLB[395] WLB[394]
+WLB[393] WLB[392] WLB[391] WLB[390] WLB[389] WLB[388] WLB[387] WLB[386] WLB[385] WLB[384]
+WLB[383] WLB[382] WLB[381] WLB[380] WLB[379] WLB[378] WLB[377] WLB[376] WLB[375] WLB[374]
+WLB[373] WLB[372] WLB[371] WLB[370] WLB[369] WLB[368] WLB[367] WLB[366] WLB[365] WLB[364]
+WLB[363] WLB[362] WLB[361] WLB[360] WLB[359] WLB[358] WLB[357] WLB[356] WLB[355] WLB[354]
+WLB[353] WLB[352] WLB[351] WLB[350] WLB[349] WLB[348] WLB[347] WLB[346] WLB[345] WLB[344]
+WLB[343] WLB[342] WLB[341] WLB[340] WLB[339] WLB[338] WLB[337] WLB[336] WLB[335] WLB[334]
+WLB[333] WLB[332] WLB[331] WLB[330] WLB[329] WLB[328] WLB[327] WLB[326] WLB[325] WLB[324]
+WLB[323] WLB[322] WLB[321] WLB[320] WLB[319] WLB[318] WLB[317] WLB[316] WLB[315] WLB[314]
+WLB[313] WLB[312] WLB[311] WLB[310] WLB[309] WLB[308] WLB[307] WLB[306] WLB[305] WLB[304]
+WLB[303] WLB[302] WLB[301] WLB[300] WLB[299] WLB[298] WLB[297] WLB[296] WLB[295] WLB[294]
+WLB[293] WLB[292] WLB[291] WLB[290] WLB[289] WLB[288] WLB[287] WLB[286] WLB[285] WLB[284]
+WLB[283] WLB[282] WLB[281] WLB[280] WLB[279] WLB[278] WLB[277] WLB[276] WLB[275] WLB[274]
+WLB[273] WLB[272] WLB[271] WLB[270] WLB[269] WLB[268] WLB[267] WLB[266] WLB[265] WLB[264]
+WLB[263] WLB[262] WLB[261] WLB[260] WLB[259] WLB[258] WLB[257] WLB[256] WLB[255] WLB[254]
+WLB[253] WLB[252] WLB[251] WLB[250] WLB[249] WLB[248] WLB[247] WLB[246] WLB[245] WLB[244]
+WLB[243] WLB[242] WLB[241] WLB[240] WLB[239] WLB[238] WLB[237] WLB[236] WLB[235] WLB[234]
+WLB[233] WLB[232] WLB[231] WLB[230] WLB[229] WLB[228] WLB[227] WLB[226] WLB[225] WLB[224]
+WLB[223] WLB[222] WLB[221] WLB[220] WLB[219] WLB[218] WLB[217] WLB[216] WLB[215] WLB[214]
+WLB[213] WLB[212] WLB[211] WLB[210] WLB[209] WLB[208] WLB[207] WLB[206] WLB[205] WLB[204]
+WLB[203] WLB[202] WLB[201] WLB[200] WLB[199] WLB[198] WLB[197] WLB[196] WLB[195] WLB[194]
+WLB[193] WLB[192] WLB[191] WLB[190] WLB[189] WLB[188] WLB[187] WLB[186] WLB[185] WLB[184]
+WLB[183] WLB[182] WLB[181] WLB[180] WLB[179] WLB[178] WLB[177] WLB[176] WLB[175] WLB[174]
+WLB[173] WLB[172] WLB[171] WLB[170] WLB[169] WLB[168] WLB[167] WLB[166] WLB[165] WLB[164]
+WLB[163] WLB[162] WLB[161] WLB[160] WLB[159] WLB[158] WLB[157] WLB[156] WLB[155] WLB[154]
+WLB[153] WLB[152] WLB[151] WLB[150] WLB[149] WLB[148] WLB[147] WLB[146] WLB[145] WLB[144]
+WLB[143] WLB[142] WLB[141] WLB[140] WLB[139] WLB[138] WLB[137] WLB[136] WLB[135] WLB[134]
+WLB[133] WLB[132] WLB[131] WLB[130] WLB[129] WLB[128] WLB[127] WLB[126] WLB[125] WLB[124]
+WLB[123] WLB[122] WLB[121] WLB[120] WLB[119] WLB[118] WLB[117] WLB[116] WLB[115] WLB[114]
+WLB[113] WLB[112] WLB[111] WLB[110] WLB[109] WLB[108] WLB[107] WLB[106] WLB[105] WLB[104]
+WLB[103] WLB[102] WLB[101] WLB[100] WLB[99] WLB[98] WLB[97] WLB[96] WLB[95] WLB[94]
+WLB[93] WLB[92] WLB[91] WLB[90] WLB[89] WLB[88] WLB[87] WLB[86] WLB[85] WLB[84]
+WLB[83] WLB[82] WLB[81] WLB[80] WLB[79] WLB[78] WLB[77] WLB[76] WLB[75] WLB[74]
+WLB[73] WLB[72] WLB[71] WLB[70] WLB[69] WLB[68] WLB[67] WLB[66] WLB[65] WLB[64]
+WLB[63] WLB[62] WLB[61] WLB[60] WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54]
+WLB[53] WLB[52] WLB[51] WLB[50] WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44]
+WLB[43] WLB[42] WLB[41] WLB[40] WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34]
+WLB[33] WLB[32] WLB[31] WLB[30] WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24]
+WLB[23] WLB[22] WLB[21] WLB[20] WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14]
+WLB[13] WLB[12] WLB[11] WLB[10] WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4]
+WLB[3] WLB[2] WLB[1] WLB[0] YXA[7] YXA[6] YXA[5] YXA[4] YXA[3] YXA[2]
+YXA[1] YXA[0] YXB[7] YXB[6] YXB[5] YXB[4] YXB[3] YXB[2] YXB[1] YXB[0]
XI0 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] RDWLA[3] RDWLA[2] RDWLA[1] RDWLA[0] RDWLB[3] RDWLB[2] RDWLB[1] RDWLB[0]
+RWLA[0] RWLA[1] RWLB[0] RWLB[1] VDD VSS WLA[511] WLA[510] WLA[509] WLA[508]
+WLA[507] WLA[506] WLA[505] WLA[504] WLA[503] WLA[502] WLA[501] WLA[500] WLA[499] WLA[498]
+WLA[497] WLA[496] WLA[495] WLA[494] WLA[493] WLA[492] WLA[491] WLA[490] WLA[489] WLA[488]
+WLA[487] WLA[486] WLA[485] WLA[484] WLA[483] WLA[482] WLA[481] WLA[480] WLA[479] WLA[478]
+WLA[477] WLA[476] WLA[475] WLA[474] WLA[473] WLA[472] WLA[471] WLA[470] WLA[469] WLA[468]
+WLA[467] WLA[466] WLA[465] WLA[464] WLA[463] WLA[462] WLA[461] WLA[460] WLA[459] WLA[458]
+WLA[457] WLA[456] WLA[455] WLA[454] WLA[453] WLA[452] WLA[451] WLA[450] WLA[449] WLA[448]
+WLA[447] WLA[446] WLA[445] WLA[444] WLA[443] WLA[442] WLA[441] WLA[440] WLA[439] WLA[438]
+WLA[437] WLA[436] WLA[435] WLA[434] WLA[433] WLA[432] WLA[431] WLA[430] WLA[429] WLA[428]
+WLA[427] WLA[426] WLA[425] WLA[424] WLA[423] WLA[422] WLA[421] WLA[420] WLA[419] WLA[418]
+WLA[417] WLA[416] WLA[415] WLA[414] WLA[413] WLA[412] WLA[411] WLA[410] WLA[409] WLA[408]
+WLA[407] WLA[406] WLA[405] WLA[404] WLA[403] WLA[402] WLA[401] WLA[400] WLA[399] WLA[398]
+WLA[397] WLA[396] WLA[395] WLA[394] WLA[393] WLA[392] WLA[391] WLA[390] WLA[389] WLA[388]
+WLA[387] WLA[386] WLA[385] WLA[384] WLA[383] WLA[382] WLA[381] WLA[380] WLA[379] WLA[378]
+WLA[377] WLA[376] WLA[375] WLA[374] WLA[373] WLA[372] WLA[371] WLA[370] WLA[369] WLA[368]
+WLA[367] WLA[366] WLA[365] WLA[364] WLA[363] WLA[362] WLA[361] WLA[360] WLA[359] WLA[358]
+WLA[357] WLA[356] WLA[355] WLA[354] WLA[353] WLA[352] WLA[351] WLA[350] WLA[349] WLA[348]
+WLA[347] WLA[346] WLA[345] WLA[344] WLA[343] WLA[342] WLA[341] WLA[340] WLA[339] WLA[338]
+WLA[337] WLA[336] WLA[335] WLA[334] WLA[333] WLA[332] WLA[331] WLA[330] WLA[329] WLA[328]
+WLA[327] WLA[326] WLA[325] WLA[324] WLA[323] WLA[322] WLA[321] WLA[320] WLA[319] WLA[318]
+WLA[317] WLA[316] WLA[315] WLA[314] WLA[313] WLA[312] WLA[311] WLA[310] WLA[309] WLA[308]
+WLA[307] WLA[306] WLA[305] WLA[304] WLA[303] WLA[302] WLA[301] WLA[300] WLA[299] WLA[298]
+WLA[297] WLA[296] WLA[295] WLA[294] WLA[293] WLA[292] WLA[291] WLA[290] WLA[289] WLA[288]
+WLA[287] WLA[286] WLA[285] WLA[284] WLA[283] WLA[282] WLA[281] WLA[280] WLA[279] WLA[278]
+WLA[277] WLA[276] WLA[275] WLA[274] WLA[273] WLA[272] WLA[271] WLA[270] WLA[269] WLA[268]
+WLA[267] WLA[266] WLA[265] WLA[264] WLA[263] WLA[262] WLA[261] WLA[260] WLA[259] WLA[258]
+WLA[257] WLA[256] WLA[255] WLA[254] WLA[253] WLA[252] WLA[251] WLA[250] WLA[249] WLA[248]
+WLA[247] WLA[246] WLA[245] WLA[244] WLA[243] WLA[242] WLA[241] WLA[240] WLA[239] WLA[238]
+WLA[237] WLA[236] WLA[235] WLA[234] WLA[233] WLA[232] WLA[231] WLA[230] WLA[229] WLA[228]
+WLA[227] WLA[226] WLA[225] WLA[224] WLA[223] WLA[222] WLA[221] WLA[220] WLA[219] WLA[218]
+WLA[217] WLA[216] WLA[215] WLA[214] WLA[213] WLA[212] WLA[211] WLA[210] WLA[209] WLA[208]
+WLA[207] WLA[206] WLA[205] WLA[204] WLA[203] WLA[202] WLA[201] WLA[200] WLA[199] WLA[198]
+WLA[197] WLA[196] WLA[195] WLA[194] WLA[193] WLA[192] WLA[191] WLA[190] WLA[189] WLA[188]
+WLA[187] WLA[186] WLA[185] WLA[184] WLA[183] WLA[182] WLA[181] WLA[180] WLA[179] WLA[178]
+WLA[177] WLA[176] WLA[175] WLA[174] WLA[173] WLA[172] WLA[171] WLA[170] WLA[169] WLA[168]
+WLA[167] WLA[166] WLA[165] WLA[164] WLA[163] WLA[162] WLA[161] WLA[160] WLA[159] WLA[158]
+WLA[157] WLA[156] WLA[155] WLA[154] WLA[153] WLA[152] WLA[151] WLA[150] WLA[149] WLA[148]
+WLA[147] WLA[146] WLA[145] WLA[144] WLA[143] WLA[142] WLA[141] WLA[140] WLA[139] WLA[138]
+WLA[137] WLA[136] WLA[135] WLA[134] WLA[133] WLA[132] WLA[131] WLA[130] WLA[129] WLA[128]
+WLA[127] WLA[126] WLA[125] WLA[124] WLA[123] WLA[122] WLA[121] WLA[120] WLA[119] WLA[118]
+WLA[117] WLA[116] WLA[115] WLA[114] WLA[113] WLA[112] WLA[111] WLA[110] WLA[109] WLA[108]
+WLA[107] WLA[106] WLA[105] WLA[104] WLA[103] WLA[102] WLA[101] WLA[100] WLA[99] WLA[98]
+WLA[97] WLA[96] WLA[95] WLA[94] WLA[93] WLA[92] WLA[91] WLA[90] WLA[89] WLA[88]
+WLA[87] WLA[86] WLA[85] WLA[84] WLA[83] WLA[82] WLA[81] WLA[80] WLA[79] WLA[78]
+WLA[77] WLA[76] WLA[75] WLA[74] WLA[73] WLA[72] WLA[71] WLA[70] WLA[69] WLA[68]
+WLA[67] WLA[66] WLA[65] WLA[64] WLA[63] WLA[62] WLA[61] WLA[60] WLA[59] WLA[58]
+WLA[57] WLA[56] WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48]
+WLA[47] WLA[46] WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38]
+WLA[37] WLA[36] WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28]
+WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18]
+WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8]
+WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] WLB[511] WLB[510]
+WLB[509] WLB[508] WLB[507] WLB[506] WLB[505] WLB[504] WLB[503] WLB[502] WLB[501] WLB[500]
+WLB[499] WLB[498] WLB[497] WLB[496] WLB[495] WLB[494] WLB[493] WLB[492] WLB[491] WLB[490]
+WLB[489] WLB[488] WLB[487] WLB[486] WLB[485] WLB[484] WLB[483] WLB[482] WLB[481] WLB[480]
+WLB[479] WLB[478] WLB[477] WLB[476] WLB[475] WLB[474] WLB[473] WLB[472] WLB[471] WLB[470]
+WLB[469] WLB[468] WLB[467] WLB[466] WLB[465] WLB[464] WLB[463] WLB[462] WLB[461] WLB[460]
+WLB[459] WLB[458] WLB[457] WLB[456] WLB[455] WLB[454] WLB[453] WLB[452] WLB[451] WLB[450]
+WLB[449] WLB[448] WLB[447] WLB[446] WLB[445] WLB[444] WLB[443] WLB[442] WLB[441] WLB[440]
+WLB[439] WLB[438] WLB[437] WLB[436] WLB[435] WLB[434] WLB[433] WLB[432] WLB[431] WLB[430]
+WLB[429] WLB[428] WLB[427] WLB[426] WLB[425] WLB[424] WLB[423] WLB[422] WLB[421] WLB[420]
+WLB[419] WLB[418] WLB[417] WLB[416] WLB[415] WLB[414] WLB[413] WLB[412] WLB[411] WLB[410]
+WLB[409] WLB[408] WLB[407] WLB[406] WLB[405] WLB[404] WLB[403] WLB[402] WLB[401] WLB[400]
+WLB[399] WLB[398] WLB[397] WLB[396] WLB[395] WLB[394] WLB[393] WLB[392] WLB[391] WLB[390]
+WLB[389] WLB[388] WLB[387] WLB[386] WLB[385] WLB[384] WLB[383] WLB[382] WLB[381] WLB[380]
+WLB[379] WLB[378] WLB[377] WLB[376] WLB[375] WLB[374] WLB[373] WLB[372] WLB[371] WLB[370]
+WLB[369] WLB[368] WLB[367] WLB[366] WLB[365] WLB[364] WLB[363] WLB[362] WLB[361] WLB[360]
+WLB[359] WLB[358] WLB[357] WLB[356] WLB[355] WLB[354] WLB[353] WLB[352] WLB[351] WLB[350]
+WLB[349] WLB[348] WLB[347] WLB[346] WLB[345] WLB[344] WLB[343] WLB[342] WLB[341] WLB[340]
+WLB[339] WLB[338] WLB[337] WLB[336] WLB[335] WLB[334] WLB[333] WLB[332] WLB[331] WLB[330]
+WLB[329] WLB[328] WLB[327] WLB[326] WLB[325] WLB[324] WLB[323] WLB[322] WLB[321] WLB[320]
+WLB[319] WLB[318] WLB[317] WLB[316] WLB[315] WLB[314] WLB[313] WLB[312] WLB[311] WLB[310]
+WLB[309] WLB[308] WLB[307] WLB[306] WLB[305] WLB[304] WLB[303] WLB[302] WLB[301] WLB[300]
+WLB[299] WLB[298] WLB[297] WLB[296] WLB[295] WLB[294] WLB[293] WLB[292] WLB[291] WLB[290]
+WLB[289] WLB[288] WLB[287] WLB[286] WLB[285] WLB[284] WLB[283] WLB[282] WLB[281] WLB[280]
+WLB[279] WLB[278] WLB[277] WLB[276] WLB[275] WLB[274] WLB[273] WLB[272] WLB[271] WLB[270]
+WLB[269] WLB[268] WLB[267] WLB[266] WLB[265] WLB[264] WLB[263] WLB[262] WLB[261] WLB[260]
+WLB[259] WLB[258] WLB[257] WLB[256] WLB[255] WLB[254] WLB[253] WLB[252] WLB[251] WLB[250]
+WLB[249] WLB[248] WLB[247] WLB[246] WLB[245] WLB[244] WLB[243] WLB[242] WLB[241] WLB[240]
+WLB[239] WLB[238] WLB[237] WLB[236] WLB[235] WLB[234] WLB[233] WLB[232] WLB[231] WLB[230]
+WLB[229] WLB[228] WLB[227] WLB[226] WLB[225] WLB[224] WLB[223] WLB[222] WLB[221] WLB[220]
+WLB[219] WLB[218] WLB[217] WLB[216] WLB[215] WLB[214] WLB[213] WLB[212] WLB[211] WLB[210]
+WLB[209] WLB[208] WLB[207] WLB[206] WLB[205] WLB[204] WLB[203] WLB[202] WLB[201] WLB[200]
+WLB[199] WLB[198] WLB[197] WLB[196] WLB[195] WLB[194] WLB[193] WLB[192] WLB[191] WLB[190]
+WLB[189] WLB[188] WLB[187] WLB[186] WLB[185] WLB[184] WLB[183] WLB[182] WLB[181] WLB[180]
+WLB[179] WLB[178] WLB[177] WLB[176] WLB[175] WLB[174] WLB[173] WLB[172] WLB[171] WLB[170]
+WLB[169] WLB[168] WLB[167] WLB[166] WLB[165] WLB[164] WLB[163] WLB[162] WLB[161] WLB[160]
+WLB[159] WLB[158] WLB[157] WLB[156] WLB[155] WLB[154] WLB[153] WLB[152] WLB[151] WLB[150]
+WLB[149] WLB[148] WLB[147] WLB[146] WLB[145] WLB[144] WLB[143] WLB[142] WLB[141] WLB[140]
+WLB[139] WLB[138] WLB[137] WLB[136] WLB[135] WLB[134] WLB[133] WLB[132] WLB[131] WLB[130]
+WLB[129] WLB[128] WLB[127] WLB[126] WLB[125] WLB[124] WLB[123] WLB[122] WLB[121] WLB[120]
+WLB[119] WLB[118] WLB[117] WLB[116] WLB[115] WLB[114] WLB[113] WLB[112] WLB[111] WLB[110]
+WLB[109] WLB[108] WLB[107] WLB[106] WLB[105] WLB[104] WLB[103] WLB[102] WLB[101] WLB[100]
+WLB[99] WLB[98] WLB[97] WLB[96] WLB[95] WLB[94] WLB[93] WLB[92] WLB[91] WLB[90]
+WLB[89] WLB[88] WLB[87] WLB[86] WLB[85] WLB[84] WLB[83] WLB[82] WLB[81] WLB[80]
+WLB[79] WLB[78] WLB[77] WLB[76] WLB[75] WLB[74] WLB[73] WLB[72] WLB[71] WLB[70]
+WLB[69] WLB[68] WLB[67] WLB[66] WLB[65] WLB[64] WLB[63] WLB[62] WLB[61] WLB[60]
+WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54] WLB[53] WLB[52] WLB[51] WLB[50]
+WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44] WLB[43] WLB[42] WLB[41] WLB[40]
+WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34] WLB[33] WLB[32] WLB[31] WLB[30]
+WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24] WLB[23] WLB[22] WLB[21] WLB[20]
+WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14] WLB[13] WLB[12] WLB[11] WLB[10]
+WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4] WLB[3] WLB[2] WLB[1] WLB[0] S55NLLGDPH_X512Y8D16_BW_ARRAY512X8
XI1 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] BWENA BWENB CLKA CLKB CLKXA CLKXB DATAA DATAB
+DOUTA DOUTB SACK1A SACK1B SACK4A SACK4B VDD VSS WEA WEB
+YXA[7] YXA[6] YXA[5] YXA[4] YXA[3] YXA[2] YXA[1] YXA[0] YXB[7] YXB[6]
+YXB[5] YXB[4] YXB[3] YXB[2] YXB[1] YXB[0] S55NLLGDPH_X512Y8D16_BW_YMX8SAWRA_B_BW
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    S55NLLGDPH_X512Y8D16_BW_BITCELL68X8A_MID
* View Name:    schematic
************************************************************************

.SUBCKT S55NLLGDPH_X512Y8D16_BW_BITCELL68X8A_MID BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] RDWLA[3] RDWLA[2] RDWLA[1] RDWLA[0] RDWLA_MID[3] RDWLA_MID[2] RDWLA_MID[1] RDWLA_MID[0]
+RDWLB[3] RDWLB[2] RDWLB[1] RDWLB[0] RDWLB_MID[3] RDWLB_MID[2] RDWLB_MID[1] RDWLB_MID[0] VDD VSS
+WLA[63] WLA[62] WLA[61] WLA[60] WLA[59] WLA[58] WLA[57] WLA[56] WLA[55] WLA[54]
+WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48] WLA[47] WLA[46] WLA[45] WLA[44]
+WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38] WLA[37] WLA[36] WLA[35] WLA[34]
+WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28] WLA[27] WLA[26] WLA[25] WLA[24]
+WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18] WLA[17] WLA[16] WLA[15] WLA[14]
+WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8] WLA[7] WLA[6] WLA[5] WLA[4]
+WLA[3] WLA[2] WLA[1] WLA[0] WLB[63] WLB[62] WLB[61] WLB[60] WLB[59] WLB[58]
+WLB[57] WLB[56] WLB[55] WLB[54] WLB[53] WLB[52] WLB[51] WLB[50] WLB[49] WLB[48]
+WLB[47] WLB[46] WLB[45] WLB[44] WLB[43] WLB[42] WLB[41] WLB[40] WLB[39] WLB[38]
+WLB[37] WLB[36] WLB[35] WLB[34] WLB[33] WLB[32] WLB[31] WLB[30] WLB[29] WLB[28]
+WLB[27] WLB[26] WLB[25] WLB[24] WLB[23] WLB[22] WLB[21] WLB[20] WLB[19] WLB[18]
+WLB[17] WLB[16] WLB[15] WLB[14] WLB[13] WLB[12] WLB[11] WLB[10] WLB[9] WLB[8]
+WLB[7] WLB[6] WLB[5] WLB[4] WLB[3] WLB[2] WLB[1] WLB[0]
XI0 BLB[0] STRAP[0] BLXB[0] STRAPX[0] VDD VSS RDWLA[3] RDWLA[2] RDWLA[1] RDWLA[0]
+RDWLB[3] RDWLB[2] RDWLB[1] RDWLB[0] S55NLLGDPH_X512Y8D16_BW_BITCELL2X2_STWL
XI1 BLB[0] BLXB[0] VDD VSS S55NLLGDPH_X512Y8D16_BW_BLSTRAP
XI2 STRAP[0] STRAPX[0] VDD VSS S55NLLGDPH_X512Y8D16_BW_BLSTRAP
XI3 BLB[1] STRAP[1] BLXB[1] STRAPX[1] VDD VSS RDWLA[3] RDWLA[2] RDWLA[1] RDWLA[0]
+RDWLB[3] RDWLB[2] RDWLB[1] RDWLB[0] S55NLLGDPH_X512Y8D16_BW_BITCELL2X2_STWL
XI4 BLB[1] BLXB[1] VDD VSS S55NLLGDPH_X512Y8D16_BW_BLSTRAP
XI5 STRAP[1] STRAPX[1] VDD VSS S55NLLGDPH_X512Y8D16_BW_BLSTRAP
XI6 BLB[2] STRAP[2] BLXB[2] STRAPX[2] VDD VSS RDWLA[3] RDWLA[2] RDWLA[1] RDWLA[0]
+RDWLB[3] RDWLB[2] RDWLB[1] RDWLB[0] S55NLLGDPH_X512Y8D16_BW_BITCELL2X2_STWL
XI7 BLB[2] BLXB[2] VDD VSS S55NLLGDPH_X512Y8D16_BW_BLSTRAP
XI8 STRAP[2] STRAPX[2] VDD VSS S55NLLGDPH_X512Y8D16_BW_BLSTRAP
XI9 BLB[3] STRAP[3] BLXB[3] STRAPX[3] VDD VSS RDWLA[3] RDWLA[2] RDWLA[1] RDWLA[0]
+RDWLB[3] RDWLB[2] RDWLB[1] RDWLB[0] S55NLLGDPH_X512Y8D16_BW_BITCELL2X2_STWL
XI10 BLB[3] BLXB[3] VDD VSS S55NLLGDPH_X512Y8D16_BW_BLSTRAP
XI11 STRAP[3] STRAPX[3] VDD VSS S55NLLGDPH_X512Y8D16_BW_BLSTRAP
XI12 BLB[4] STRAP[4] BLXB[4] STRAPX[4] VDD VSS RDWLA[3] RDWLA[2] RDWLA[1] RDWLA[0]
+RDWLB[3] RDWLB[2] RDWLB[1] RDWLB[0] S55NLLGDPH_X512Y8D16_BW_BITCELL2X2_STWL
XI13 BLB[4] BLXB[4] VDD VSS S55NLLGDPH_X512Y8D16_BW_BLSTRAP
XI14 STRAP[4] STRAPX[4] VDD VSS S55NLLGDPH_X512Y8D16_BW_BLSTRAP
XI15 BLB[5] STRAP[5] BLXB[5] STRAPX[5] VDD VSS RDWLA[3] RDWLA[2] RDWLA[1] RDWLA[0]
+RDWLB[3] RDWLB[2] RDWLB[1] RDWLB[0] S55NLLGDPH_X512Y8D16_BW_BITCELL2X2_STWL
XI16 BLB[5] BLXB[5] VDD VSS S55NLLGDPH_X512Y8D16_BW_BLSTRAP
XI17 STRAP[5] STRAPX[5] VDD VSS S55NLLGDPH_X512Y8D16_BW_BLSTRAP
XI18 BLB[6] STRAP[6] BLXB[6] STRAPX[6] VDD VSS RDWLA_MID[3] RDWLA_MID[2] RDWLA_MID[1] RDWLA_MID[0]
+RDWLB_MID[3] RDWLB_MID[2] RDWLB_MID[1] RDWLB_MID[0] S55NLLGDPH_X512Y8D16_BW_BITCELL2X2_STWL
XI19 BLB[6] BLXB[6] VDD VSS S55NLLGDPH_X512Y8D16_BW_BLSTRAP
XI20 STRAP[6] STRAPX[6] VDD VSS S55NLLGDPH_X512Y8D16_BW_BLSTRAP
XI21 BLB[7] STRAP[7] BLXB[7] STRAPX[7] VDD VSS RDWLA[3] RDWLA[2] RDWLA[1] RDWLA[0]
+RDWLB[3] RDWLB[2] RDWLB[1] RDWLB[0] S55NLLGDPH_X512Y8D16_BW_BITCELL2X2_STWL
XI22 BLB[7] BLXB[7] VDD VSS S55NLLGDPH_X512Y8D16_BW_BLSTRAP
XI23 STRAP[7] STRAPX[7] VDD VSS S55NLLGDPH_X512Y8D16_BW_BLSTRAP
XI24 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[1] WLA[0] WLB[1] WLB[0] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI25 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[3] WLA[2] WLB[3] WLB[2] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI26 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[5] WLA[4] WLB[5] WLB[4] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI27 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[7] WLA[6] WLB[7] WLB[6] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI28 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[9] WLA[8] WLB[9] WLB[8] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI29 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[11] WLA[10] WLB[11] WLB[10] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI30 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[13] WLA[12] WLB[13] WLB[12] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI31 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[15] WLA[14] WLB[15] WLB[14] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI32 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[17] WLA[16] WLB[17] WLB[16] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI33 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[19] WLA[18] WLB[19] WLB[18] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI34 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[21] WLA[20] WLB[21] WLB[20] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI35 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[23] WLA[22] WLB[23] WLB[22] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI36 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[25] WLA[24] WLB[25] WLB[24] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI37 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[27] WLA[26] WLB[27] WLB[26] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI38 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[29] WLA[28] WLB[29] WLB[28] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI39 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[31] WLA[30] WLB[31] WLB[30] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI40 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[33] WLA[32] WLB[33] WLB[32] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI41 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[35] WLA[34] WLB[35] WLB[34] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI42 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[37] WLA[36] WLB[37] WLB[36] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI43 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[39] WLA[38] WLB[39] WLB[38] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI44 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[41] WLA[40] WLB[41] WLB[40] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI45 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[43] WLA[42] WLB[43] WLB[42] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI46 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[45] WLA[44] WLB[45] WLB[44] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI47 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[47] WLA[46] WLB[47] WLB[46] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI48 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[49] WLA[48] WLB[49] WLB[48] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI49 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[51] WLA[50] WLB[51] WLB[50] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI50 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[53] WLA[52] WLB[53] WLB[52] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI51 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[55] WLA[54] WLB[55] WLB[54] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI52 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[57] WLA[56] WLB[57] WLB[56] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI53 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[59] WLA[58] WLB[59] WLB[58] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI54 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[61] WLA[60] WLB[61] WLB[60] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
XI55 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[63] WLA[62] WLB[63] WLB[62] S55NLLGDPH_X512Y8D16_BW_BITCELL2X8
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    S55NLLGDPH_X512Y8D16_BW_ARRAY512X8_MID
* View Name:    schematic
************************************************************************

.SUBCKT S55NLLGDPH_X512Y8D16_BW_ARRAY512X8_MID BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] RDWLA[3] RDWLA[2] RDWLA[1] RDWLA[0] RDWLA_MID[3] RDWLA_MID[2] RDWLA_MID[1] RDWLA_MID[0]
+RDWLB[3] RDWLB[2] RDWLB[1] RDWLB[0] RDWLB_MID[3] RDWLB_MID[2] RDWLB_MID[1] RDWLB_MID[0] RWLA[0] RWLA[1]
+RWLB[0] RWLB[1] VDD VSS WLA[511] WLA[510] WLA[509] WLA[508] WLA[507] WLA[506]
+WLA[505] WLA[504] WLA[503] WLA[502] WLA[501] WLA[500] WLA[499] WLA[498] WLA[497] WLA[496]
+WLA[495] WLA[494] WLA[493] WLA[492] WLA[491] WLA[490] WLA[489] WLA[488] WLA[487] WLA[486]
+WLA[485] WLA[484] WLA[483] WLA[482] WLA[481] WLA[480] WLA[479] WLA[478] WLA[477] WLA[476]
+WLA[475] WLA[474] WLA[473] WLA[472] WLA[471] WLA[470] WLA[469] WLA[468] WLA[467] WLA[466]
+WLA[465] WLA[464] WLA[463] WLA[462] WLA[461] WLA[460] WLA[459] WLA[458] WLA[457] WLA[456]
+WLA[455] WLA[454] WLA[453] WLA[452] WLA[451] WLA[450] WLA[449] WLA[448] WLA[447] WLA[446]
+WLA[445] WLA[444] WLA[443] WLA[442] WLA[441] WLA[440] WLA[439] WLA[438] WLA[437] WLA[436]
+WLA[435] WLA[434] WLA[433] WLA[432] WLA[431] WLA[430] WLA[429] WLA[428] WLA[427] WLA[426]
+WLA[425] WLA[424] WLA[423] WLA[422] WLA[421] WLA[420] WLA[419] WLA[418] WLA[417] WLA[416]
+WLA[415] WLA[414] WLA[413] WLA[412] WLA[411] WLA[410] WLA[409] WLA[408] WLA[407] WLA[406]
+WLA[405] WLA[404] WLA[403] WLA[402] WLA[401] WLA[400] WLA[399] WLA[398] WLA[397] WLA[396]
+WLA[395] WLA[394] WLA[393] WLA[392] WLA[391] WLA[390] WLA[389] WLA[388] WLA[387] WLA[386]
+WLA[385] WLA[384] WLA[383] WLA[382] WLA[381] WLA[380] WLA[379] WLA[378] WLA[377] WLA[376]
+WLA[375] WLA[374] WLA[373] WLA[372] WLA[371] WLA[370] WLA[369] WLA[368] WLA[367] WLA[366]
+WLA[365] WLA[364] WLA[363] WLA[362] WLA[361] WLA[360] WLA[359] WLA[358] WLA[357] WLA[356]
+WLA[355] WLA[354] WLA[353] WLA[352] WLA[351] WLA[350] WLA[349] WLA[348] WLA[347] WLA[346]
+WLA[345] WLA[344] WLA[343] WLA[342] WLA[341] WLA[340] WLA[339] WLA[338] WLA[337] WLA[336]
+WLA[335] WLA[334] WLA[333] WLA[332] WLA[331] WLA[330] WLA[329] WLA[328] WLA[327] WLA[326]
+WLA[325] WLA[324] WLA[323] WLA[322] WLA[321] WLA[320] WLA[319] WLA[318] WLA[317] WLA[316]
+WLA[315] WLA[314] WLA[313] WLA[312] WLA[311] WLA[310] WLA[309] WLA[308] WLA[307] WLA[306]
+WLA[305] WLA[304] WLA[303] WLA[302] WLA[301] WLA[300] WLA[299] WLA[298] WLA[297] WLA[296]
+WLA[295] WLA[294] WLA[293] WLA[292] WLA[291] WLA[290] WLA[289] WLA[288] WLA[287] WLA[286]
+WLA[285] WLA[284] WLA[283] WLA[282] WLA[281] WLA[280] WLA[279] WLA[278] WLA[277] WLA[276]
+WLA[275] WLA[274] WLA[273] WLA[272] WLA[271] WLA[270] WLA[269] WLA[268] WLA[267] WLA[266]
+WLA[265] WLA[264] WLA[263] WLA[262] WLA[261] WLA[260] WLA[259] WLA[258] WLA[257] WLA[256]
+WLA[255] WLA[254] WLA[253] WLA[252] WLA[251] WLA[250] WLA[249] WLA[248] WLA[247] WLA[246]
+WLA[245] WLA[244] WLA[243] WLA[242] WLA[241] WLA[240] WLA[239] WLA[238] WLA[237] WLA[236]
+WLA[235] WLA[234] WLA[233] WLA[232] WLA[231] WLA[230] WLA[229] WLA[228] WLA[227] WLA[226]
+WLA[225] WLA[224] WLA[223] WLA[222] WLA[221] WLA[220] WLA[219] WLA[218] WLA[217] WLA[216]
+WLA[215] WLA[214] WLA[213] WLA[212] WLA[211] WLA[210] WLA[209] WLA[208] WLA[207] WLA[206]
+WLA[205] WLA[204] WLA[203] WLA[202] WLA[201] WLA[200] WLA[199] WLA[198] WLA[197] WLA[196]
+WLA[195] WLA[194] WLA[193] WLA[192] WLA[191] WLA[190] WLA[189] WLA[188] WLA[187] WLA[186]
+WLA[185] WLA[184] WLA[183] WLA[182] WLA[181] WLA[180] WLA[179] WLA[178] WLA[177] WLA[176]
+WLA[175] WLA[174] WLA[173] WLA[172] WLA[171] WLA[170] WLA[169] WLA[168] WLA[167] WLA[166]
+WLA[165] WLA[164] WLA[163] WLA[162] WLA[161] WLA[160] WLA[159] WLA[158] WLA[157] WLA[156]
+WLA[155] WLA[154] WLA[153] WLA[152] WLA[151] WLA[150] WLA[149] WLA[148] WLA[147] WLA[146]
+WLA[145] WLA[144] WLA[143] WLA[142] WLA[141] WLA[140] WLA[139] WLA[138] WLA[137] WLA[136]
+WLA[135] WLA[134] WLA[133] WLA[132] WLA[131] WLA[130] WLA[129] WLA[128] WLA[127] WLA[126]
+WLA[125] WLA[124] WLA[123] WLA[122] WLA[121] WLA[120] WLA[119] WLA[118] WLA[117] WLA[116]
+WLA[115] WLA[114] WLA[113] WLA[112] WLA[111] WLA[110] WLA[109] WLA[108] WLA[107] WLA[106]
+WLA[105] WLA[104] WLA[103] WLA[102] WLA[101] WLA[100] WLA[99] WLA[98] WLA[97] WLA[96]
+WLA[95] WLA[94] WLA[93] WLA[92] WLA[91] WLA[90] WLA[89] WLA[88] WLA[87] WLA[86]
+WLA[85] WLA[84] WLA[83] WLA[82] WLA[81] WLA[80] WLA[79] WLA[78] WLA[77] WLA[76]
+WLA[75] WLA[74] WLA[73] WLA[72] WLA[71] WLA[70] WLA[69] WLA[68] WLA[67] WLA[66]
+WLA[65] WLA[64] WLA[63] WLA[62] WLA[61] WLA[60] WLA[59] WLA[58] WLA[57] WLA[56]
+WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48] WLA[47] WLA[46]
+WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38] WLA[37] WLA[36]
+WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28] WLA[27] WLA[26]
+WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18] WLA[17] WLA[16]
+WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8] WLA[7] WLA[6]
+WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] WLB[511] WLB[510] WLB[509] WLB[508]
+WLB[507] WLB[506] WLB[505] WLB[504] WLB[503] WLB[502] WLB[501] WLB[500] WLB[499] WLB[498]
+WLB[497] WLB[496] WLB[495] WLB[494] WLB[493] WLB[492] WLB[491] WLB[490] WLB[489] WLB[488]
+WLB[487] WLB[486] WLB[485] WLB[484] WLB[483] WLB[482] WLB[481] WLB[480] WLB[479] WLB[478]
+WLB[477] WLB[476] WLB[475] WLB[474] WLB[473] WLB[472] WLB[471] WLB[470] WLB[469] WLB[468]
+WLB[467] WLB[466] WLB[465] WLB[464] WLB[463] WLB[462] WLB[461] WLB[460] WLB[459] WLB[458]
+WLB[457] WLB[456] WLB[455] WLB[454] WLB[453] WLB[452] WLB[451] WLB[450] WLB[449] WLB[448]
+WLB[447] WLB[446] WLB[445] WLB[444] WLB[443] WLB[442] WLB[441] WLB[440] WLB[439] WLB[438]
+WLB[437] WLB[436] WLB[435] WLB[434] WLB[433] WLB[432] WLB[431] WLB[430] WLB[429] WLB[428]
+WLB[427] WLB[426] WLB[425] WLB[424] WLB[423] WLB[422] WLB[421] WLB[420] WLB[419] WLB[418]
+WLB[417] WLB[416] WLB[415] WLB[414] WLB[413] WLB[412] WLB[411] WLB[410] WLB[409] WLB[408]
+WLB[407] WLB[406] WLB[405] WLB[404] WLB[403] WLB[402] WLB[401] WLB[400] WLB[399] WLB[398]
+WLB[397] WLB[396] WLB[395] WLB[394] WLB[393] WLB[392] WLB[391] WLB[390] WLB[389] WLB[388]
+WLB[387] WLB[386] WLB[385] WLB[384] WLB[383] WLB[382] WLB[381] WLB[380] WLB[379] WLB[378]
+WLB[377] WLB[376] WLB[375] WLB[374] WLB[373] WLB[372] WLB[371] WLB[370] WLB[369] WLB[368]
+WLB[367] WLB[366] WLB[365] WLB[364] WLB[363] WLB[362] WLB[361] WLB[360] WLB[359] WLB[358]
+WLB[357] WLB[356] WLB[355] WLB[354] WLB[353] WLB[352] WLB[351] WLB[350] WLB[349] WLB[348]
+WLB[347] WLB[346] WLB[345] WLB[344] WLB[343] WLB[342] WLB[341] WLB[340] WLB[339] WLB[338]
+WLB[337] WLB[336] WLB[335] WLB[334] WLB[333] WLB[332] WLB[331] WLB[330] WLB[329] WLB[328]
+WLB[327] WLB[326] WLB[325] WLB[324] WLB[323] WLB[322] WLB[321] WLB[320] WLB[319] WLB[318]
+WLB[317] WLB[316] WLB[315] WLB[314] WLB[313] WLB[312] WLB[311] WLB[310] WLB[309] WLB[308]
+WLB[307] WLB[306] WLB[305] WLB[304] WLB[303] WLB[302] WLB[301] WLB[300] WLB[299] WLB[298]
+WLB[297] WLB[296] WLB[295] WLB[294] WLB[293] WLB[292] WLB[291] WLB[290] WLB[289] WLB[288]
+WLB[287] WLB[286] WLB[285] WLB[284] WLB[283] WLB[282] WLB[281] WLB[280] WLB[279] WLB[278]
+WLB[277] WLB[276] WLB[275] WLB[274] WLB[273] WLB[272] WLB[271] WLB[270] WLB[269] WLB[268]
+WLB[267] WLB[266] WLB[265] WLB[264] WLB[263] WLB[262] WLB[261] WLB[260] WLB[259] WLB[258]
+WLB[257] WLB[256] WLB[255] WLB[254] WLB[253] WLB[252] WLB[251] WLB[250] WLB[249] WLB[248]
+WLB[247] WLB[246] WLB[245] WLB[244] WLB[243] WLB[242] WLB[241] WLB[240] WLB[239] WLB[238]
+WLB[237] WLB[236] WLB[235] WLB[234] WLB[233] WLB[232] WLB[231] WLB[230] WLB[229] WLB[228]
+WLB[227] WLB[226] WLB[225] WLB[224] WLB[223] WLB[222] WLB[221] WLB[220] WLB[219] WLB[218]
+WLB[217] WLB[216] WLB[215] WLB[214] WLB[213] WLB[212] WLB[211] WLB[210] WLB[209] WLB[208]
+WLB[207] WLB[206] WLB[205] WLB[204] WLB[203] WLB[202] WLB[201] WLB[200] WLB[199] WLB[198]
+WLB[197] WLB[196] WLB[195] WLB[194] WLB[193] WLB[192] WLB[191] WLB[190] WLB[189] WLB[188]
+WLB[187] WLB[186] WLB[185] WLB[184] WLB[183] WLB[182] WLB[181] WLB[180] WLB[179] WLB[178]
+WLB[177] WLB[176] WLB[175] WLB[174] WLB[173] WLB[172] WLB[171] WLB[170] WLB[169] WLB[168]
+WLB[167] WLB[166] WLB[165] WLB[164] WLB[163] WLB[162] WLB[161] WLB[160] WLB[159] WLB[158]
+WLB[157] WLB[156] WLB[155] WLB[154] WLB[153] WLB[152] WLB[151] WLB[150] WLB[149] WLB[148]
+WLB[147] WLB[146] WLB[145] WLB[144] WLB[143] WLB[142] WLB[141] WLB[140] WLB[139] WLB[138]
+WLB[137] WLB[136] WLB[135] WLB[134] WLB[133] WLB[132] WLB[131] WLB[130] WLB[129] WLB[128]
+WLB[127] WLB[126] WLB[125] WLB[124] WLB[123] WLB[122] WLB[121] WLB[120] WLB[119] WLB[118]
+WLB[117] WLB[116] WLB[115] WLB[114] WLB[113] WLB[112] WLB[111] WLB[110] WLB[109] WLB[108]
+WLB[107] WLB[106] WLB[105] WLB[104] WLB[103] WLB[102] WLB[101] WLB[100] WLB[99] WLB[98]
+WLB[97] WLB[96] WLB[95] WLB[94] WLB[93] WLB[92] WLB[91] WLB[90] WLB[89] WLB[88]
+WLB[87] WLB[86] WLB[85] WLB[84] WLB[83] WLB[82] WLB[81] WLB[80] WLB[79] WLB[78]
+WLB[77] WLB[76] WLB[75] WLB[74] WLB[73] WLB[72] WLB[71] WLB[70] WLB[69] WLB[68]
+WLB[67] WLB[66] WLB[65] WLB[64] WLB[63] WLB[62] WLB[61] WLB[60] WLB[59] WLB[58]
+WLB[57] WLB[56] WLB[55] WLB[54] WLB[53] WLB[52] WLB[51] WLB[50] WLB[49] WLB[48]
+WLB[47] WLB[46] WLB[45] WLB[44] WLB[43] WLB[42] WLB[41] WLB[40] WLB[39] WLB[38]
+WLB[37] WLB[36] WLB[35] WLB[34] WLB[33] WLB[32] WLB[31] WLB[30] WLB[29] WLB[28]
+WLB[27] WLB[26] WLB[25] WLB[24] WLB[23] WLB[22] WLB[21] WLB[20] WLB[19] WLB[18]
+WLB[17] WLB[16] WLB[15] WLB[14] WLB[13] WLB[12] WLB[11] WLB[10] WLB[9] WLB[8]
+WLB[7] WLB[6] WLB[5] WLB[4] WLB[3] WLB[2] WLB[1] WLB[0]
XI0 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] RWLA[0] RWLA[1] RWLB[0] RWLB[1] VDD VSS WLA[63] WLA[62]
+WLA[61] WLA[60] WLA[59] WLA[58] WLA[57] WLA[56] WLA[55] WLA[54] WLA[53] WLA[52]
+WLA[51] WLA[50] WLA[49] WLA[48] WLA[47] WLA[46] WLA[45] WLA[44] WLA[43] WLA[42]
+WLA[41] WLA[40] WLA[39] WLA[38] WLA[37] WLA[36] WLA[35] WLA[34] WLA[33] WLA[32]
+WLA[31] WLA[30] WLA[29] WLA[28] WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22]
+WLA[21] WLA[20] WLA[19] WLA[18] WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12]
+WLA[11] WLA[10] WLA[9] WLA[8] WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2]
+WLA[1] WLA[0] WLB[63] WLB[62] WLB[61] WLB[60] WLB[59] WLB[58] WLB[57] WLB[56]
+WLB[55] WLB[54] WLB[53] WLB[52] WLB[51] WLB[50] WLB[49] WLB[48] WLB[47] WLB[46]
+WLB[45] WLB[44] WLB[43] WLB[42] WLB[41] WLB[40] WLB[39] WLB[38] WLB[37] WLB[36]
+WLB[35] WLB[34] WLB[33] WLB[32] WLB[31] WLB[30] WLB[29] WLB[28] WLB[27] WLB[26]
+WLB[25] WLB[24] WLB[23] WLB[22] WLB[21] WLB[20] WLB[19] WLB[18] WLB[17] WLB[16]
+WLB[15] WLB[14] WLB[13] WLB[12] WLB[11] WLB[10] WLB[9] WLB[8] WLB[7] WLB[6]
+WLB[5] WLB[4] WLB[3] WLB[2] WLB[1] WLB[0] S55NLLGDPH_X512Y8D16_BW_BITCELL66X8B_RED
XI1 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[127] WLA[126] WLA[125] WLA[124] WLA[123] WLA[122]
+WLA[121] WLA[120] WLA[119] WLA[118] WLA[117] WLA[116] WLA[115] WLA[114] WLA[113] WLA[112]
+WLA[111] WLA[110] WLA[109] WLA[108] WLA[107] WLA[106] WLA[105] WLA[104] WLA[103] WLA[102]
+WLA[101] WLA[100] WLA[99] WLA[98] WLA[97] WLA[96] WLA[95] WLA[94] WLA[93] WLA[92]
+WLA[91] WLA[90] WLA[89] WLA[88] WLA[87] WLA[86] WLA[85] WLA[84] WLA[83] WLA[82]
+WLA[81] WLA[80] WLA[79] WLA[78] WLA[77] WLA[76] WLA[75] WLA[74] WLA[73] WLA[72]
+WLA[71] WLA[70] WLA[69] WLA[68] WLA[67] WLA[66] WLA[65] WLA[64] WLB[127] WLB[126]
+WLB[125] WLB[124] WLB[123] WLB[122] WLB[121] WLB[120] WLB[119] WLB[118] WLB[117] WLB[116]
+WLB[115] WLB[114] WLB[113] WLB[112] WLB[111] WLB[110] WLB[109] WLB[108] WLB[107] WLB[106]
+WLB[105] WLB[104] WLB[103] WLB[102] WLB[101] WLB[100] WLB[99] WLB[98] WLB[97] WLB[96]
+WLB[95] WLB[94] WLB[93] WLB[92] WLB[91] WLB[90] WLB[89] WLB[88] WLB[87] WLB[86]
+WLB[85] WLB[84] WLB[83] WLB[82] WLB[81] WLB[80] WLB[79] WLB[78] WLB[77] WLB[76]
+WLB[75] WLB[74] WLB[73] WLB[72] WLB[71] WLB[70] WLB[69] WLB[68] WLB[67] WLB[66]
+WLB[65] WLB[64] S55NLLGDPH_X512Y8D16_BW_BITCELL64X8A
XI2 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[191] WLA[190] WLA[189] WLA[188] WLA[187] WLA[186]
+WLA[185] WLA[184] WLA[183] WLA[182] WLA[181] WLA[180] WLA[179] WLA[178] WLA[177] WLA[176]
+WLA[175] WLA[174] WLA[173] WLA[172] WLA[171] WLA[170] WLA[169] WLA[168] WLA[167] WLA[166]
+WLA[165] WLA[164] WLA[163] WLA[162] WLA[161] WLA[160] WLA[159] WLA[158] WLA[157] WLA[156]
+WLA[155] WLA[154] WLA[153] WLA[152] WLA[151] WLA[150] WLA[149] WLA[148] WLA[147] WLA[146]
+WLA[145] WLA[144] WLA[143] WLA[142] WLA[141] WLA[140] WLA[139] WLA[138] WLA[137] WLA[136]
+WLA[135] WLA[134] WLA[133] WLA[132] WLA[131] WLA[130] WLA[129] WLA[128] WLB[191] WLB[190]
+WLB[189] WLB[188] WLB[187] WLB[186] WLB[185] WLB[184] WLB[183] WLB[182] WLB[181] WLB[180]
+WLB[179] WLB[178] WLB[177] WLB[176] WLB[175] WLB[174] WLB[173] WLB[172] WLB[171] WLB[170]
+WLB[169] WLB[168] WLB[167] WLB[166] WLB[165] WLB[164] WLB[163] WLB[162] WLB[161] WLB[160]
+WLB[159] WLB[158] WLB[157] WLB[156] WLB[155] WLB[154] WLB[153] WLB[152] WLB[151] WLB[150]
+WLB[149] WLB[148] WLB[147] WLB[146] WLB[145] WLB[144] WLB[143] WLB[142] WLB[141] WLB[140]
+WLB[139] WLB[138] WLB[137] WLB[136] WLB[135] WLB[134] WLB[133] WLB[132] WLB[131] WLB[130]
+WLB[129] WLB[128] S55NLLGDPH_X512Y8D16_BW_BITCELL64X8B
XI3 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] VDD VSS WLA[255] WLA[254] WLA[253] WLA[252] WLA[251] WLA[250]
+WLA[249] WLA[248] WLA[247] WLA[246] WLA[245] WLA[244] WLA[243] WLA[242] WLA[241] WLA[240]
+WLA[239] WLA[238] WLA[237] WLA[236] WLA[235] WLA[234] WLA[233] WLA[232] WLA[231] WLA[230]
+WLA[229] WLA[228] WLA[227] WLA[226] WLA[225] WLA[224] WLA[223] WLA[222] WLA[221] WLA[220]
+WLA[219] WLA[218] WLA[217] WLA[216] WLA[215] WLA[214] WLA[213] WLA[212] WLA[211] WLA[210]
+WLA[209] WLA[208] WLA[207] WLA[206] WLA[205] WLA[204] WLA[203] WLA[202] WLA[201] WLA[200]
+WLA[199] WLA[198] WLA[197] WLA[196] WLA[195] WLA[194] WLA[193] WLA[192] WLB[255] WLB[254]
+WLB[253] WLB[252] WLB[251] WLB[250] WLB[249] WLB[248] WLB[247] WLB[246] WLB[245] WLB[244]
+WLB[243] WLB[242] WLB[241] WLB[240] WLB[239] WLB[238] WLB[237] WLB[236] WLB[235] WLB[234]
+WLB[233] WLB[232] WLB[231] WLB[230] WLB[229] WLB[228] WLB[227] WLB[226] WLB[225] WLB[224]
+WLB[223] WLB[222] WLB[221] WLB[220] WLB[219] WLB[218] WLB[217] WLB[216] WLB[215] WLB[214]
+WLB[213] WLB[212] WLB[211] WLB[210] WLB[209] WLB[208] WLB[207] WLB[206] WLB[205] WLB[204]
+WLB[203] WLB[202] WLB[201] WLB[200] WLB[199] WLB[198] WLB[197] WLB[196] WLB[195] WLB[194]
+WLB[193] WLB[192] S55NLLGDPH_X512Y8D16_BW_BITCELL64X8A
XI4 BLXA[7] BLXA[6] BLXA[5] BLXA[4] BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6]
+BLXB[5] BLXB[4] BLXB[3] BLXB[2] BLXB[1] BLXB[0] BLA[7] BLA[6] BLA[5] BLA[4]
+BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6] BLB[5] BLB[4] BLB[3] BLB[2]
+BLB[1] BLB[0] VDD VSS WLA[319] WLA[318] WLA[317] WLA[316] WLA[315] WLA[314]
+WLA[313] WLA[312] WLA[311] WLA[310] WLA[309] WLA[308] WLA[307] WLA[306] WLA[305] WLA[304]
+WLA[303] WLA[302] WLA[301] WLA[300] WLA[299] WLA[298] WLA[297] WLA[296] WLA[295] WLA[294]
+WLA[293] WLA[292] WLA[291] WLA[290] WLA[289] WLA[288] WLA[287] WLA[286] WLA[285] WLA[284]
+WLA[283] WLA[282] WLA[281] WLA[280] WLA[279] WLA[278] WLA[277] WLA[276] WLA[275] WLA[274]
+WLA[273] WLA[272] WLA[271] WLA[270] WLA[269] WLA[268] WLA[267] WLA[266] WLA[265] WLA[264]
+WLA[263] WLA[262] WLA[261] WLA[260] WLA[259] WLA[258] WLA[257] WLA[256] WLB[319] WLB[318]
+WLB[317] WLB[316] WLB[315] WLB[314] WLB[313] WLB[312] WLB[311] WLB[310] WLB[309] WLB[308]
+WLB[307] WLB[306] WLB[305] WLB[304] WLB[303] WLB[302] WLB[301] WLB[300] WLB[299] WLB[298]
+WLB[297] WLB[296] WLB[295] WLB[294] WLB[293] WLB[292] WLB[291] WLB[290] WLB[289] WLB[288]
+WLB[287] WLB[286] WLB[285] WLB[284] WLB[283] WLB[282] WLB[281] WLB[280] WLB[279] WLB[278]
+WLB[277] WLB[276] WLB[275] WLB[274] WLB[273] WLB[272] WLB[271] WLB[270] WLB[269] WLB[268]
+WLB[267] WLB[266] WLB[265] WLB[264] WLB[263] WLB[262] WLB[261] WLB[260] WLB[259] WLB[258]
+WLB[257] WLB[256] S55NLLGDPH_X512Y8D16_BW_BITCELL64X8B
XI5 BLXA[7] BLXA[6] BLXA[5] BLXA[4] BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6]
+BLXB[5] BLXB[4] BLXB[3] BLXB[2] BLXB[1] BLXB[0] BLA[7] BLA[6] BLA[5] BLA[4]
+BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6] BLB[5] BLB[4] BLB[3] BLB[2]
+BLB[1] BLB[0] VDD VSS WLA[383] WLA[382] WLA[381] WLA[380] WLA[379] WLA[378]
+WLA[377] WLA[376] WLA[375] WLA[374] WLA[373] WLA[372] WLA[371] WLA[370] WLA[369] WLA[368]
+WLA[367] WLA[366] WLA[365] WLA[364] WLA[363] WLA[362] WLA[361] WLA[360] WLA[359] WLA[358]
+WLA[357] WLA[356] WLA[355] WLA[354] WLA[353] WLA[352] WLA[351] WLA[350] WLA[349] WLA[348]
+WLA[347] WLA[346] WLA[345] WLA[344] WLA[343] WLA[342] WLA[341] WLA[340] WLA[339] WLA[338]
+WLA[337] WLA[336] WLA[335] WLA[334] WLA[333] WLA[332] WLA[331] WLA[330] WLA[329] WLA[328]
+WLA[327] WLA[326] WLA[325] WLA[324] WLA[323] WLA[322] WLA[321] WLA[320] WLB[383] WLB[382]
+WLB[381] WLB[380] WLB[379] WLB[378] WLB[377] WLB[376] WLB[375] WLB[374] WLB[373] WLB[372]
+WLB[371] WLB[370] WLB[369] WLB[368] WLB[367] WLB[366] WLB[365] WLB[364] WLB[363] WLB[362]
+WLB[361] WLB[360] WLB[359] WLB[358] WLB[357] WLB[356] WLB[355] WLB[354] WLB[353] WLB[352]
+WLB[351] WLB[350] WLB[349] WLB[348] WLB[347] WLB[346] WLB[345] WLB[344] WLB[343] WLB[342]
+WLB[341] WLB[340] WLB[339] WLB[338] WLB[337] WLB[336] WLB[335] WLB[334] WLB[333] WLB[332]
+WLB[331] WLB[330] WLB[329] WLB[328] WLB[327] WLB[326] WLB[325] WLB[324] WLB[323] WLB[322]
+WLB[321] WLB[320] S55NLLGDPH_X512Y8D16_BW_BITCELL64X8A
XI6 BLXA[7] BLXA[6] BLXA[5] BLXA[4] BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6]
+BLXB[5] BLXB[4] BLXB[3] BLXB[2] BLXB[1] BLXB[0] BLA[7] BLA[6] BLA[5] BLA[4]
+BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6] BLB[5] BLB[4] BLB[3] BLB[2]
+BLB[1] BLB[0] VDD VSS WLA[447] WLA[446] WLA[445] WLA[444] WLA[443] WLA[442]
+WLA[441] WLA[440] WLA[439] WLA[438] WLA[437] WLA[436] WLA[435] WLA[434] WLA[433] WLA[432]
+WLA[431] WLA[430] WLA[429] WLA[428] WLA[427] WLA[426] WLA[425] WLA[424] WLA[423] WLA[422]
+WLA[421] WLA[420] WLA[419] WLA[418] WLA[417] WLA[416] WLA[415] WLA[414] WLA[413] WLA[412]
+WLA[411] WLA[410] WLA[409] WLA[408] WLA[407] WLA[406] WLA[405] WLA[404] WLA[403] WLA[402]
+WLA[401] WLA[400] WLA[399] WLA[398] WLA[397] WLA[396] WLA[395] WLA[394] WLA[393] WLA[392]
+WLA[391] WLA[390] WLA[389] WLA[388] WLA[387] WLA[386] WLA[385] WLA[384] WLB[447] WLB[446]
+WLB[445] WLB[444] WLB[443] WLB[442] WLB[441] WLB[440] WLB[439] WLB[438] WLB[437] WLB[436]
+WLB[435] WLB[434] WLB[433] WLB[432] WLB[431] WLB[430] WLB[429] WLB[428] WLB[427] WLB[426]
+WLB[425] WLB[424] WLB[423] WLB[422] WLB[421] WLB[420] WLB[419] WLB[418] WLB[417] WLB[416]
+WLB[415] WLB[414] WLB[413] WLB[412] WLB[411] WLB[410] WLB[409] WLB[408] WLB[407] WLB[406]
+WLB[405] WLB[404] WLB[403] WLB[402] WLB[401] WLB[400] WLB[399] WLB[398] WLB[397] WLB[396]
+WLB[395] WLB[394] WLB[393] WLB[392] WLB[391] WLB[390] WLB[389] WLB[388] WLB[387] WLB[386]
+WLB[385] WLB[384] S55NLLGDPH_X512Y8D16_BW_BITCELL64X8B
XI7 BLXA[7] BLXA[6] BLXA[5] BLXA[4] BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6]
+BLXB[5] BLXB[4] BLXB[3] BLXB[2] BLXB[1] BLXB[0] BLA[7] BLA[6] BLA[5] BLA[4]
+BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6] BLB[5] BLB[4] BLB[3] BLB[2]
+BLB[1] BLB[0] RDWLA[3] RDWLA[2] RDWLA[1] RDWLA[0] RDWLA_MID[3] RDWLA_MID[2] RDWLA_MID[1] RDWLA_MID[0]
+RDWLB[3] RDWLB[2] RDWLB[1] RDWLB[0] RDWLB_MID[3] RDWLB_MID[2] RDWLB_MID[1] RDWLB_MID[0] VDD VSS
+WLA[511] WLA[510] WLA[509] WLA[508] WLA[507] WLA[506] WLA[505] WLA[504] WLA[503] WLA[502]
+WLA[501] WLA[500] WLA[499] WLA[498] WLA[497] WLA[496] WLA[495] WLA[494] WLA[493] WLA[492]
+WLA[491] WLA[490] WLA[489] WLA[488] WLA[487] WLA[486] WLA[485] WLA[484] WLA[483] WLA[482]
+WLA[481] WLA[480] WLA[479] WLA[478] WLA[477] WLA[476] WLA[475] WLA[474] WLA[473] WLA[472]
+WLA[471] WLA[470] WLA[469] WLA[468] WLA[467] WLA[466] WLA[465] WLA[464] WLA[463] WLA[462]
+WLA[461] WLA[460] WLA[459] WLA[458] WLA[457] WLA[456] WLA[455] WLA[454] WLA[453] WLA[452]
+WLA[451] WLA[450] WLA[449] WLA[448] WLB[511] WLB[510] WLB[509] WLB[508] WLB[507] WLB[506]
+WLB[505] WLB[504] WLB[503] WLB[502] WLB[501] WLB[500] WLB[499] WLB[498] WLB[497] WLB[496]
+WLB[495] WLB[494] WLB[493] WLB[492] WLB[491] WLB[490] WLB[489] WLB[488] WLB[487] WLB[486]
+WLB[485] WLB[484] WLB[483] WLB[482] WLB[481] WLB[480] WLB[479] WLB[478] WLB[477] WLB[476]
+WLB[475] WLB[474] WLB[473] WLB[472] WLB[471] WLB[470] WLB[469] WLB[468] WLB[467] WLB[466]
+WLB[465] WLB[464] WLB[463] WLB[462] WLB[461] WLB[460] WLB[459] WLB[458] WLB[457] WLB[456]
+WLB[455] WLB[454] WLB[453] WLB[452] WLB[451] WLB[450] WLB[449] WLB[448] S55NLLGDPH_X512Y8D16_BW_BITCELL68X8A_MID
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    S55NLLGDPH_X512Y8D16_BW_Y512X8CELL_MID
* View Name:    schematic
************************************************************************

.SUBCKT S55NLLGDPH_X512Y8D16_BW_Y512X8CELL_MID BWENA BWENB CLKA CLKB CLKXA CLKXB DATAA DATAB DOUTA DOUTB
+RDWLA[3] RDWLA[2] RDWLA[1] RDWLA[0] RDWLA_MID[3] RDWLA_MID[2] RDWLA_MID[1] RDWLA_MID[0] RDWLB[3] RDWLB[2]
+RDWLB[1] RDWLB[0] RDWLB_MID[3] RDWLB_MID[2] RDWLB_MID[1] RDWLB_MID[0] RWLA[0] RWLA[1] RWLB[0] RWLB[1]
+SACK1A SACK1B SACK4A SACK4B VDD VSS WEA WEB WLA[511] WLA[510]
+WLA[509] WLA[508] WLA[507] WLA[506] WLA[505] WLA[504] WLA[503] WLA[502] WLA[501] WLA[500]
+WLA[499] WLA[498] WLA[497] WLA[496] WLA[495] WLA[494] WLA[493] WLA[492] WLA[491] WLA[490]
+WLA[489] WLA[488] WLA[487] WLA[486] WLA[485] WLA[484] WLA[483] WLA[482] WLA[481] WLA[480]
+WLA[479] WLA[478] WLA[477] WLA[476] WLA[475] WLA[474] WLA[473] WLA[472] WLA[471] WLA[470]
+WLA[469] WLA[468] WLA[467] WLA[466] WLA[465] WLA[464] WLA[463] WLA[462] WLA[461] WLA[460]
+WLA[459] WLA[458] WLA[457] WLA[456] WLA[455] WLA[454] WLA[453] WLA[452] WLA[451] WLA[450]
+WLA[449] WLA[448] WLA[447] WLA[446] WLA[445] WLA[444] WLA[443] WLA[442] WLA[441] WLA[440]
+WLA[439] WLA[438] WLA[437] WLA[436] WLA[435] WLA[434] WLA[433] WLA[432] WLA[431] WLA[430]
+WLA[429] WLA[428] WLA[427] WLA[426] WLA[425] WLA[424] WLA[423] WLA[422] WLA[421] WLA[420]
+WLA[419] WLA[418] WLA[417] WLA[416] WLA[415] WLA[414] WLA[413] WLA[412] WLA[411] WLA[410]
+WLA[409] WLA[408] WLA[407] WLA[406] WLA[405] WLA[404] WLA[403] WLA[402] WLA[401] WLA[400]
+WLA[399] WLA[398] WLA[397] WLA[396] WLA[395] WLA[394] WLA[393] WLA[392] WLA[391] WLA[390]
+WLA[389] WLA[388] WLA[387] WLA[386] WLA[385] WLA[384] WLA[383] WLA[382] WLA[381] WLA[380]
+WLA[379] WLA[378] WLA[377] WLA[376] WLA[375] WLA[374] WLA[373] WLA[372] WLA[371] WLA[370]
+WLA[369] WLA[368] WLA[367] WLA[366] WLA[365] WLA[364] WLA[363] WLA[362] WLA[361] WLA[360]
+WLA[359] WLA[358] WLA[357] WLA[356] WLA[355] WLA[354] WLA[353] WLA[352] WLA[351] WLA[350]
+WLA[349] WLA[348] WLA[347] WLA[346] WLA[345] WLA[344] WLA[343] WLA[342] WLA[341] WLA[340]
+WLA[339] WLA[338] WLA[337] WLA[336] WLA[335] WLA[334] WLA[333] WLA[332] WLA[331] WLA[330]
+WLA[329] WLA[328] WLA[327] WLA[326] WLA[325] WLA[324] WLA[323] WLA[322] WLA[321] WLA[320]
+WLA[319] WLA[318] WLA[317] WLA[316] WLA[315] WLA[314] WLA[313] WLA[312] WLA[311] WLA[310]
+WLA[309] WLA[308] WLA[307] WLA[306] WLA[305] WLA[304] WLA[303] WLA[302] WLA[301] WLA[300]
+WLA[299] WLA[298] WLA[297] WLA[296] WLA[295] WLA[294] WLA[293] WLA[292] WLA[291] WLA[290]
+WLA[289] WLA[288] WLA[287] WLA[286] WLA[285] WLA[284] WLA[283] WLA[282] WLA[281] WLA[280]
+WLA[279] WLA[278] WLA[277] WLA[276] WLA[275] WLA[274] WLA[273] WLA[272] WLA[271] WLA[270]
+WLA[269] WLA[268] WLA[267] WLA[266] WLA[265] WLA[264] WLA[263] WLA[262] WLA[261] WLA[260]
+WLA[259] WLA[258] WLA[257] WLA[256] WLA[255] WLA[254] WLA[253] WLA[252] WLA[251] WLA[250]
+WLA[249] WLA[248] WLA[247] WLA[246] WLA[245] WLA[244] WLA[243] WLA[242] WLA[241] WLA[240]
+WLA[239] WLA[238] WLA[237] WLA[236] WLA[235] WLA[234] WLA[233] WLA[232] WLA[231] WLA[230]
+WLA[229] WLA[228] WLA[227] WLA[226] WLA[225] WLA[224] WLA[223] WLA[222] WLA[221] WLA[220]
+WLA[219] WLA[218] WLA[217] WLA[216] WLA[215] WLA[214] WLA[213] WLA[212] WLA[211] WLA[210]
+WLA[209] WLA[208] WLA[207] WLA[206] WLA[205] WLA[204] WLA[203] WLA[202] WLA[201] WLA[200]
+WLA[199] WLA[198] WLA[197] WLA[196] WLA[195] WLA[194] WLA[193] WLA[192] WLA[191] WLA[190]
+WLA[189] WLA[188] WLA[187] WLA[186] WLA[185] WLA[184] WLA[183] WLA[182] WLA[181] WLA[180]
+WLA[179] WLA[178] WLA[177] WLA[176] WLA[175] WLA[174] WLA[173] WLA[172] WLA[171] WLA[170]
+WLA[169] WLA[168] WLA[167] WLA[166] WLA[165] WLA[164] WLA[163] WLA[162] WLA[161] WLA[160]
+WLA[159] WLA[158] WLA[157] WLA[156] WLA[155] WLA[154] WLA[153] WLA[152] WLA[151] WLA[150]
+WLA[149] WLA[148] WLA[147] WLA[146] WLA[145] WLA[144] WLA[143] WLA[142] WLA[141] WLA[140]
+WLA[139] WLA[138] WLA[137] WLA[136] WLA[135] WLA[134] WLA[133] WLA[132] WLA[131] WLA[130]
+WLA[129] WLA[128] WLA[127] WLA[126] WLA[125] WLA[124] WLA[123] WLA[122] WLA[121] WLA[120]
+WLA[119] WLA[118] WLA[117] WLA[116] WLA[115] WLA[114] WLA[113] WLA[112] WLA[111] WLA[110]
+WLA[109] WLA[108] WLA[107] WLA[106] WLA[105] WLA[104] WLA[103] WLA[102] WLA[101] WLA[100]
+WLA[99] WLA[98] WLA[97] WLA[96] WLA[95] WLA[94] WLA[93] WLA[92] WLA[91] WLA[90]
+WLA[89] WLA[88] WLA[87] WLA[86] WLA[85] WLA[84] WLA[83] WLA[82] WLA[81] WLA[80]
+WLA[79] WLA[78] WLA[77] WLA[76] WLA[75] WLA[74] WLA[73] WLA[72] WLA[71] WLA[70]
+WLA[69] WLA[68] WLA[67] WLA[66] WLA[65] WLA[64] WLA[63] WLA[62] WLA[61] WLA[60]
+WLA[59] WLA[58] WLA[57] WLA[56] WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50]
+WLA[49] WLA[48] WLA[47] WLA[46] WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40]
+WLA[39] WLA[38] WLA[37] WLA[36] WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30]
+WLA[29] WLA[28] WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20]
+WLA[19] WLA[18] WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10]
+WLA[9] WLA[8] WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0]
+WLB[511] WLB[510] WLB[509] WLB[508] WLB[507] WLB[506] WLB[505] WLB[504] WLB[503] WLB[502]
+WLB[501] WLB[500] WLB[499] WLB[498] WLB[497] WLB[496] WLB[495] WLB[494] WLB[493] WLB[492]
+WLB[491] WLB[490] WLB[489] WLB[488] WLB[487] WLB[486] WLB[485] WLB[484] WLB[483] WLB[482]
+WLB[481] WLB[480] WLB[479] WLB[478] WLB[477] WLB[476] WLB[475] WLB[474] WLB[473] WLB[472]
+WLB[471] WLB[470] WLB[469] WLB[468] WLB[467] WLB[466] WLB[465] WLB[464] WLB[463] WLB[462]
+WLB[461] WLB[460] WLB[459] WLB[458] WLB[457] WLB[456] WLB[455] WLB[454] WLB[453] WLB[452]
+WLB[451] WLB[450] WLB[449] WLB[448] WLB[447] WLB[446] WLB[445] WLB[444] WLB[443] WLB[442]
+WLB[441] WLB[440] WLB[439] WLB[438] WLB[437] WLB[436] WLB[435] WLB[434] WLB[433] WLB[432]
+WLB[431] WLB[430] WLB[429] WLB[428] WLB[427] WLB[426] WLB[425] WLB[424] WLB[423] WLB[422]
+WLB[421] WLB[420] WLB[419] WLB[418] WLB[417] WLB[416] WLB[415] WLB[414] WLB[413] WLB[412]
+WLB[411] WLB[410] WLB[409] WLB[408] WLB[407] WLB[406] WLB[405] WLB[404] WLB[403] WLB[402]
+WLB[401] WLB[400] WLB[399] WLB[398] WLB[397] WLB[396] WLB[395] WLB[394] WLB[393] WLB[392]
+WLB[391] WLB[390] WLB[389] WLB[388] WLB[387] WLB[386] WLB[385] WLB[384] WLB[383] WLB[382]
+WLB[381] WLB[380] WLB[379] WLB[378] WLB[377] WLB[376] WLB[375] WLB[374] WLB[373] WLB[372]
+WLB[371] WLB[370] WLB[369] WLB[368] WLB[367] WLB[366] WLB[365] WLB[364] WLB[363] WLB[362]
+WLB[361] WLB[360] WLB[359] WLB[358] WLB[357] WLB[356] WLB[355] WLB[354] WLB[353] WLB[352]
+WLB[351] WLB[350] WLB[349] WLB[348] WLB[347] WLB[346] WLB[345] WLB[344] WLB[343] WLB[342]
+WLB[341] WLB[340] WLB[339] WLB[338] WLB[337] WLB[336] WLB[335] WLB[334] WLB[333] WLB[332]
+WLB[331] WLB[330] WLB[329] WLB[328] WLB[327] WLB[326] WLB[325] WLB[324] WLB[323] WLB[322]
+WLB[321] WLB[320] WLB[319] WLB[318] WLB[317] WLB[316] WLB[315] WLB[314] WLB[313] WLB[312]
+WLB[311] WLB[310] WLB[309] WLB[308] WLB[307] WLB[306] WLB[305] WLB[304] WLB[303] WLB[302]
+WLB[301] WLB[300] WLB[299] WLB[298] WLB[297] WLB[296] WLB[295] WLB[294] WLB[293] WLB[292]
+WLB[291] WLB[290] WLB[289] WLB[288] WLB[287] WLB[286] WLB[285] WLB[284] WLB[283] WLB[282]
+WLB[281] WLB[280] WLB[279] WLB[278] WLB[277] WLB[276] WLB[275] WLB[274] WLB[273] WLB[272]
+WLB[271] WLB[270] WLB[269] WLB[268] WLB[267] WLB[266] WLB[265] WLB[264] WLB[263] WLB[262]
+WLB[261] WLB[260] WLB[259] WLB[258] WLB[257] WLB[256] WLB[255] WLB[254] WLB[253] WLB[252]
+WLB[251] WLB[250] WLB[249] WLB[248] WLB[247] WLB[246] WLB[245] WLB[244] WLB[243] WLB[242]
+WLB[241] WLB[240] WLB[239] WLB[238] WLB[237] WLB[236] WLB[235] WLB[234] WLB[233] WLB[232]
+WLB[231] WLB[230] WLB[229] WLB[228] WLB[227] WLB[226] WLB[225] WLB[224] WLB[223] WLB[222]
+WLB[221] WLB[220] WLB[219] WLB[218] WLB[217] WLB[216] WLB[215] WLB[214] WLB[213] WLB[212]
+WLB[211] WLB[210] WLB[209] WLB[208] WLB[207] WLB[206] WLB[205] WLB[204] WLB[203] WLB[202]
+WLB[201] WLB[200] WLB[199] WLB[198] WLB[197] WLB[196] WLB[195] WLB[194] WLB[193] WLB[192]
+WLB[191] WLB[190] WLB[189] WLB[188] WLB[187] WLB[186] WLB[185] WLB[184] WLB[183] WLB[182]
+WLB[181] WLB[180] WLB[179] WLB[178] WLB[177] WLB[176] WLB[175] WLB[174] WLB[173] WLB[172]
+WLB[171] WLB[170] WLB[169] WLB[168] WLB[167] WLB[166] WLB[165] WLB[164] WLB[163] WLB[162]
+WLB[161] WLB[160] WLB[159] WLB[158] WLB[157] WLB[156] WLB[155] WLB[154] WLB[153] WLB[152]
+WLB[151] WLB[150] WLB[149] WLB[148] WLB[147] WLB[146] WLB[145] WLB[144] WLB[143] WLB[142]
+WLB[141] WLB[140] WLB[139] WLB[138] WLB[137] WLB[136] WLB[135] WLB[134] WLB[133] WLB[132]
+WLB[131] WLB[130] WLB[129] WLB[128] WLB[127] WLB[126] WLB[125] WLB[124] WLB[123] WLB[122]
+WLB[121] WLB[120] WLB[119] WLB[118] WLB[117] WLB[116] WLB[115] WLB[114] WLB[113] WLB[112]
+WLB[111] WLB[110] WLB[109] WLB[108] WLB[107] WLB[106] WLB[105] WLB[104] WLB[103] WLB[102]
+WLB[101] WLB[100] WLB[99] WLB[98] WLB[97] WLB[96] WLB[95] WLB[94] WLB[93] WLB[92]
+WLB[91] WLB[90] WLB[89] WLB[88] WLB[87] WLB[86] WLB[85] WLB[84] WLB[83] WLB[82]
+WLB[81] WLB[80] WLB[79] WLB[78] WLB[77] WLB[76] WLB[75] WLB[74] WLB[73] WLB[72]
+WLB[71] WLB[70] WLB[69] WLB[68] WLB[67] WLB[66] WLB[65] WLB[64] WLB[63] WLB[62]
+WLB[61] WLB[60] WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54] WLB[53] WLB[52]
+WLB[51] WLB[50] WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44] WLB[43] WLB[42]
+WLB[41] WLB[40] WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34] WLB[33] WLB[32]
+WLB[31] WLB[30] WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24] WLB[23] WLB[22]
+WLB[21] WLB[20] WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14] WLB[13] WLB[12]
+WLB[11] WLB[10] WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4] WLB[3] WLB[2]
+WLB[1] WLB[0] YXA[7] YXA[6] YXA[5] YXA[4] YXA[3] YXA[2] YXA[1] YXA[0]
+YXB[7] YXB[6] YXB[5] YXB[4] YXB[3] YXB[2] YXB[1] YXB[0]
XI0 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] RDWLA[3] RDWLA[2] RDWLA[1] RDWLA[0] RDWLA_MID[3] RDWLA_MID[2] RDWLA_MID[1] RDWLA_MID[0]
+RDWLB[3] RDWLB[2] RDWLB[1] RDWLB[0] RDWLB_MID[3] RDWLB_MID[2] RDWLB_MID[1] RDWLB_MID[0] RWLA[0] RWLA[1]
+RWLB[0] RWLB[1] VDD VSS WLA[511] WLA[510] WLA[509] WLA[508] WLA[507] WLA[506]
+WLA[505] WLA[504] WLA[503] WLA[502] WLA[501] WLA[500] WLA[499] WLA[498] WLA[497] WLA[496]
+WLA[495] WLA[494] WLA[493] WLA[492] WLA[491] WLA[490] WLA[489] WLA[488] WLA[487] WLA[486]
+WLA[485] WLA[484] WLA[483] WLA[482] WLA[481] WLA[480] WLA[479] WLA[478] WLA[477] WLA[476]
+WLA[475] WLA[474] WLA[473] WLA[472] WLA[471] WLA[470] WLA[469] WLA[468] WLA[467] WLA[466]
+WLA[465] WLA[464] WLA[463] WLA[462] WLA[461] WLA[460] WLA[459] WLA[458] WLA[457] WLA[456]
+WLA[455] WLA[454] WLA[453] WLA[452] WLA[451] WLA[450] WLA[449] WLA[448] WLA[447] WLA[446]
+WLA[445] WLA[444] WLA[443] WLA[442] WLA[441] WLA[440] WLA[439] WLA[438] WLA[437] WLA[436]
+WLA[435] WLA[434] WLA[433] WLA[432] WLA[431] WLA[430] WLA[429] WLA[428] WLA[427] WLA[426]
+WLA[425] WLA[424] WLA[423] WLA[422] WLA[421] WLA[420] WLA[419] WLA[418] WLA[417] WLA[416]
+WLA[415] WLA[414] WLA[413] WLA[412] WLA[411] WLA[410] WLA[409] WLA[408] WLA[407] WLA[406]
+WLA[405] WLA[404] WLA[403] WLA[402] WLA[401] WLA[400] WLA[399] WLA[398] WLA[397] WLA[396]
+WLA[395] WLA[394] WLA[393] WLA[392] WLA[391] WLA[390] WLA[389] WLA[388] WLA[387] WLA[386]
+WLA[385] WLA[384] WLA[383] WLA[382] WLA[381] WLA[380] WLA[379] WLA[378] WLA[377] WLA[376]
+WLA[375] WLA[374] WLA[373] WLA[372] WLA[371] WLA[370] WLA[369] WLA[368] WLA[367] WLA[366]
+WLA[365] WLA[364] WLA[363] WLA[362] WLA[361] WLA[360] WLA[359] WLA[358] WLA[357] WLA[356]
+WLA[355] WLA[354] WLA[353] WLA[352] WLA[351] WLA[350] WLA[349] WLA[348] WLA[347] WLA[346]
+WLA[345] WLA[344] WLA[343] WLA[342] WLA[341] WLA[340] WLA[339] WLA[338] WLA[337] WLA[336]
+WLA[335] WLA[334] WLA[333] WLA[332] WLA[331] WLA[330] WLA[329] WLA[328] WLA[327] WLA[326]
+WLA[325] WLA[324] WLA[323] WLA[322] WLA[321] WLA[320] WLA[319] WLA[318] WLA[317] WLA[316]
+WLA[315] WLA[314] WLA[313] WLA[312] WLA[311] WLA[310] WLA[309] WLA[308] WLA[307] WLA[306]
+WLA[305] WLA[304] WLA[303] WLA[302] WLA[301] WLA[300] WLA[299] WLA[298] WLA[297] WLA[296]
+WLA[295] WLA[294] WLA[293] WLA[292] WLA[291] WLA[290] WLA[289] WLA[288] WLA[287] WLA[286]
+WLA[285] WLA[284] WLA[283] WLA[282] WLA[281] WLA[280] WLA[279] WLA[278] WLA[277] WLA[276]
+WLA[275] WLA[274] WLA[273] WLA[272] WLA[271] WLA[270] WLA[269] WLA[268] WLA[267] WLA[266]
+WLA[265] WLA[264] WLA[263] WLA[262] WLA[261] WLA[260] WLA[259] WLA[258] WLA[257] WLA[256]
+WLA[255] WLA[254] WLA[253] WLA[252] WLA[251] WLA[250] WLA[249] WLA[248] WLA[247] WLA[246]
+WLA[245] WLA[244] WLA[243] WLA[242] WLA[241] WLA[240] WLA[239] WLA[238] WLA[237] WLA[236]
+WLA[235] WLA[234] WLA[233] WLA[232] WLA[231] WLA[230] WLA[229] WLA[228] WLA[227] WLA[226]
+WLA[225] WLA[224] WLA[223] WLA[222] WLA[221] WLA[220] WLA[219] WLA[218] WLA[217] WLA[216]
+WLA[215] WLA[214] WLA[213] WLA[212] WLA[211] WLA[210] WLA[209] WLA[208] WLA[207] WLA[206]
+WLA[205] WLA[204] WLA[203] WLA[202] WLA[201] WLA[200] WLA[199] WLA[198] WLA[197] WLA[196]
+WLA[195] WLA[194] WLA[193] WLA[192] WLA[191] WLA[190] WLA[189] WLA[188] WLA[187] WLA[186]
+WLA[185] WLA[184] WLA[183] WLA[182] WLA[181] WLA[180] WLA[179] WLA[178] WLA[177] WLA[176]
+WLA[175] WLA[174] WLA[173] WLA[172] WLA[171] WLA[170] WLA[169] WLA[168] WLA[167] WLA[166]
+WLA[165] WLA[164] WLA[163] WLA[162] WLA[161] WLA[160] WLA[159] WLA[158] WLA[157] WLA[156]
+WLA[155] WLA[154] WLA[153] WLA[152] WLA[151] WLA[150] WLA[149] WLA[148] WLA[147] WLA[146]
+WLA[145] WLA[144] WLA[143] WLA[142] WLA[141] WLA[140] WLA[139] WLA[138] WLA[137] WLA[136]
+WLA[135] WLA[134] WLA[133] WLA[132] WLA[131] WLA[130] WLA[129] WLA[128] WLA[127] WLA[126]
+WLA[125] WLA[124] WLA[123] WLA[122] WLA[121] WLA[120] WLA[119] WLA[118] WLA[117] WLA[116]
+WLA[115] WLA[114] WLA[113] WLA[112] WLA[111] WLA[110] WLA[109] WLA[108] WLA[107] WLA[106]
+WLA[105] WLA[104] WLA[103] WLA[102] WLA[101] WLA[100] WLA[99] WLA[98] WLA[97] WLA[96]
+WLA[95] WLA[94] WLA[93] WLA[92] WLA[91] WLA[90] WLA[89] WLA[88] WLA[87] WLA[86]
+WLA[85] WLA[84] WLA[83] WLA[82] WLA[81] WLA[80] WLA[79] WLA[78] WLA[77] WLA[76]
+WLA[75] WLA[74] WLA[73] WLA[72] WLA[71] WLA[70] WLA[69] WLA[68] WLA[67] WLA[66]
+WLA[65] WLA[64] WLA[63] WLA[62] WLA[61] WLA[60] WLA[59] WLA[58] WLA[57] WLA[56]
+WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48] WLA[47] WLA[46]
+WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38] WLA[37] WLA[36]
+WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28] WLA[27] WLA[26]
+WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18] WLA[17] WLA[16]
+WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8] WLA[7] WLA[6]
+WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] WLB[511] WLB[510] WLB[509] WLB[508]
+WLB[507] WLB[506] WLB[505] WLB[504] WLB[503] WLB[502] WLB[501] WLB[500] WLB[499] WLB[498]
+WLB[497] WLB[496] WLB[495] WLB[494] WLB[493] WLB[492] WLB[491] WLB[490] WLB[489] WLB[488]
+WLB[487] WLB[486] WLB[485] WLB[484] WLB[483] WLB[482] WLB[481] WLB[480] WLB[479] WLB[478]
+WLB[477] WLB[476] WLB[475] WLB[474] WLB[473] WLB[472] WLB[471] WLB[470] WLB[469] WLB[468]
+WLB[467] WLB[466] WLB[465] WLB[464] WLB[463] WLB[462] WLB[461] WLB[460] WLB[459] WLB[458]
+WLB[457] WLB[456] WLB[455] WLB[454] WLB[453] WLB[452] WLB[451] WLB[450] WLB[449] WLB[448]
+WLB[447] WLB[446] WLB[445] WLB[444] WLB[443] WLB[442] WLB[441] WLB[440] WLB[439] WLB[438]
+WLB[437] WLB[436] WLB[435] WLB[434] WLB[433] WLB[432] WLB[431] WLB[430] WLB[429] WLB[428]
+WLB[427] WLB[426] WLB[425] WLB[424] WLB[423] WLB[422] WLB[421] WLB[420] WLB[419] WLB[418]
+WLB[417] WLB[416] WLB[415] WLB[414] WLB[413] WLB[412] WLB[411] WLB[410] WLB[409] WLB[408]
+WLB[407] WLB[406] WLB[405] WLB[404] WLB[403] WLB[402] WLB[401] WLB[400] WLB[399] WLB[398]
+WLB[397] WLB[396] WLB[395] WLB[394] WLB[393] WLB[392] WLB[391] WLB[390] WLB[389] WLB[388]
+WLB[387] WLB[386] WLB[385] WLB[384] WLB[383] WLB[382] WLB[381] WLB[380] WLB[379] WLB[378]
+WLB[377] WLB[376] WLB[375] WLB[374] WLB[373] WLB[372] WLB[371] WLB[370] WLB[369] WLB[368]
+WLB[367] WLB[366] WLB[365] WLB[364] WLB[363] WLB[362] WLB[361] WLB[360] WLB[359] WLB[358]
+WLB[357] WLB[356] WLB[355] WLB[354] WLB[353] WLB[352] WLB[351] WLB[350] WLB[349] WLB[348]
+WLB[347] WLB[346] WLB[345] WLB[344] WLB[343] WLB[342] WLB[341] WLB[340] WLB[339] WLB[338]
+WLB[337] WLB[336] WLB[335] WLB[334] WLB[333] WLB[332] WLB[331] WLB[330] WLB[329] WLB[328]
+WLB[327] WLB[326] WLB[325] WLB[324] WLB[323] WLB[322] WLB[321] WLB[320] WLB[319] WLB[318]
+WLB[317] WLB[316] WLB[315] WLB[314] WLB[313] WLB[312] WLB[311] WLB[310] WLB[309] WLB[308]
+WLB[307] WLB[306] WLB[305] WLB[304] WLB[303] WLB[302] WLB[301] WLB[300] WLB[299] WLB[298]
+WLB[297] WLB[296] WLB[295] WLB[294] WLB[293] WLB[292] WLB[291] WLB[290] WLB[289] WLB[288]
+WLB[287] WLB[286] WLB[285] WLB[284] WLB[283] WLB[282] WLB[281] WLB[280] WLB[279] WLB[278]
+WLB[277] WLB[276] WLB[275] WLB[274] WLB[273] WLB[272] WLB[271] WLB[270] WLB[269] WLB[268]
+WLB[267] WLB[266] WLB[265] WLB[264] WLB[263] WLB[262] WLB[261] WLB[260] WLB[259] WLB[258]
+WLB[257] WLB[256] WLB[255] WLB[254] WLB[253] WLB[252] WLB[251] WLB[250] WLB[249] WLB[248]
+WLB[247] WLB[246] WLB[245] WLB[244] WLB[243] WLB[242] WLB[241] WLB[240] WLB[239] WLB[238]
+WLB[237] WLB[236] WLB[235] WLB[234] WLB[233] WLB[232] WLB[231] WLB[230] WLB[229] WLB[228]
+WLB[227] WLB[226] WLB[225] WLB[224] WLB[223] WLB[222] WLB[221] WLB[220] WLB[219] WLB[218]
+WLB[217] WLB[216] WLB[215] WLB[214] WLB[213] WLB[212] WLB[211] WLB[210] WLB[209] WLB[208]
+WLB[207] WLB[206] WLB[205] WLB[204] WLB[203] WLB[202] WLB[201] WLB[200] WLB[199] WLB[198]
+WLB[197] WLB[196] WLB[195] WLB[194] WLB[193] WLB[192] WLB[191] WLB[190] WLB[189] WLB[188]
+WLB[187] WLB[186] WLB[185] WLB[184] WLB[183] WLB[182] WLB[181] WLB[180] WLB[179] WLB[178]
+WLB[177] WLB[176] WLB[175] WLB[174] WLB[173] WLB[172] WLB[171] WLB[170] WLB[169] WLB[168]
+WLB[167] WLB[166] WLB[165] WLB[164] WLB[163] WLB[162] WLB[161] WLB[160] WLB[159] WLB[158]
+WLB[157] WLB[156] WLB[155] WLB[154] WLB[153] WLB[152] WLB[151] WLB[150] WLB[149] WLB[148]
+WLB[147] WLB[146] WLB[145] WLB[144] WLB[143] WLB[142] WLB[141] WLB[140] WLB[139] WLB[138]
+WLB[137] WLB[136] WLB[135] WLB[134] WLB[133] WLB[132] WLB[131] WLB[130] WLB[129] WLB[128]
+WLB[127] WLB[126] WLB[125] WLB[124] WLB[123] WLB[122] WLB[121] WLB[120] WLB[119] WLB[118]
+WLB[117] WLB[116] WLB[115] WLB[114] WLB[113] WLB[112] WLB[111] WLB[110] WLB[109] WLB[108]
+WLB[107] WLB[106] WLB[105] WLB[104] WLB[103] WLB[102] WLB[101] WLB[100] WLB[99] WLB[98]
+WLB[97] WLB[96] WLB[95] WLB[94] WLB[93] WLB[92] WLB[91] WLB[90] WLB[89] WLB[88]
+WLB[87] WLB[86] WLB[85] WLB[84] WLB[83] WLB[82] WLB[81] WLB[80] WLB[79] WLB[78]
+WLB[77] WLB[76] WLB[75] WLB[74] WLB[73] WLB[72] WLB[71] WLB[70] WLB[69] WLB[68]
+WLB[67] WLB[66] WLB[65] WLB[64] WLB[63] WLB[62] WLB[61] WLB[60] WLB[59] WLB[58]
+WLB[57] WLB[56] WLB[55] WLB[54] WLB[53] WLB[52] WLB[51] WLB[50] WLB[49] WLB[48]
+WLB[47] WLB[46] WLB[45] WLB[44] WLB[43] WLB[42] WLB[41] WLB[40] WLB[39] WLB[38]
+WLB[37] WLB[36] WLB[35] WLB[34] WLB[33] WLB[32] WLB[31] WLB[30] WLB[29] WLB[28]
+WLB[27] WLB[26] WLB[25] WLB[24] WLB[23] WLB[22] WLB[21] WLB[20] WLB[19] WLB[18]
+WLB[17] WLB[16] WLB[15] WLB[14] WLB[13] WLB[12] WLB[11] WLB[10] WLB[9] WLB[8]
+WLB[7] WLB[6] WLB[5] WLB[4] WLB[3] WLB[2] WLB[1] WLB[0] S55NLLGDPH_X512Y8D16_BW_ARRAY512X8_MID
XI1 BLA[7] BLA[6] BLA[5] BLA[4] BLA[3] BLA[2] BLA[1] BLA[0] BLB[7] BLB[6]
+BLB[5] BLB[4] BLB[3] BLB[2] BLB[1] BLB[0] BLXA[7] BLXA[6] BLXA[5] BLXA[4]
+BLXA[3] BLXA[2] BLXA[1] BLXA[0] BLXB[7] BLXB[6] BLXB[5] BLXB[4] BLXB[3] BLXB[2]
+BLXB[1] BLXB[0] BWENA BWENB CLKA CLKB CLKXA CLKXB DATAA DATAB
+DOUTA DOUTB SACK1A SACK1B SACK4A SACK4B VDD VSS WEA WEB
+YXA[7] YXA[6] YXA[5] YXA[4] YXA[3] YXA[2] YXA[1] YXA[0] YXB[7] YXB[6]
+YXB[5] YXB[4] YXB[3] YXB[2] YXB[1] YXB[0] S55NLLGDPH_X512Y8D16_BW_YMX8SAWRA_B_BW
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    S55NLLGDPH_X512Y8D16_BW_Y512X8CELLX8_BW_LEFT
* View Name:    schematic
************************************************************************

.SUBCKT S55NLLGDPH_X512Y8D16_BW_Y512X8CELLX8_BW_LEFT BWENA[7] BWENA[6] BWENA[5] BWENA[4] BWENA[3] BWENA[2] BWENA[1] BWENA[0] BWENB[7] BWENB[6]
+BWENB[5] BWENB[4] BWENB[3] BWENB[2] BWENB[1] BWENB[0] CLKA CLKB CLKXA CLKXB
+DATAA[7] DATAA[6] DATAA[5] DATAA[4] DATAA[3] DATAA[2] DATAA[1] DATAA[0] DATAB[7] DATAB[6]
+DATAB[5] DATAB[4] DATAB[3] DATAB[2] DATAB[1] DATAB[0] DBL DOUTA[7] DOUTA[6] DOUTA[5]
+DOUTA[4] DOUTA[3] DOUTA[2] DOUTA[1] DOUTA[0] DOUTB[7] DOUTB[6] DOUTB[5] DOUTB[4] DOUTB[3]
+DOUTB[2] DOUTB[1] DOUTB[0] RWLA[0] RWLA[1] RWLB[0] RWLB[1] SACK1A SACK1B SACK4A
+SACK4B STWLA STWLB VDD VSS WEA WEB WLA[511] WLA[510] WLA[509]
+WLA[508] WLA[507] WLA[506] WLA[505] WLA[504] WLA[503] WLA[502] WLA[501] WLA[500] WLA[499]
+WLA[498] WLA[497] WLA[496] WLA[495] WLA[494] WLA[493] WLA[492] WLA[491] WLA[490] WLA[489]
+WLA[488] WLA[487] WLA[486] WLA[485] WLA[484] WLA[483] WLA[482] WLA[481] WLA[480] WLA[479]
+WLA[478] WLA[477] WLA[476] WLA[475] WLA[474] WLA[473] WLA[472] WLA[471] WLA[470] WLA[469]
+WLA[468] WLA[467] WLA[466] WLA[465] WLA[464] WLA[463] WLA[462] WLA[461] WLA[460] WLA[459]
+WLA[458] WLA[457] WLA[456] WLA[455] WLA[454] WLA[453] WLA[452] WLA[451] WLA[450] WLA[449]
+WLA[448] WLA[447] WLA[446] WLA[445] WLA[444] WLA[443] WLA[442] WLA[441] WLA[440] WLA[439]
+WLA[438] WLA[437] WLA[436] WLA[435] WLA[434] WLA[433] WLA[432] WLA[431] WLA[430] WLA[429]
+WLA[428] WLA[427] WLA[426] WLA[425] WLA[424] WLA[423] WLA[422] WLA[421] WLA[420] WLA[419]
+WLA[418] WLA[417] WLA[416] WLA[415] WLA[414] WLA[413] WLA[412] WLA[411] WLA[410] WLA[409]
+WLA[408] WLA[407] WLA[406] WLA[405] WLA[404] WLA[403] WLA[402] WLA[401] WLA[400] WLA[399]
+WLA[398] WLA[397] WLA[396] WLA[395] WLA[394] WLA[393] WLA[392] WLA[391] WLA[390] WLA[389]
+WLA[388] WLA[387] WLA[386] WLA[385] WLA[384] WLA[383] WLA[382] WLA[381] WLA[380] WLA[379]
+WLA[378] WLA[377] WLA[376] WLA[375] WLA[374] WLA[373] WLA[372] WLA[371] WLA[370] WLA[369]
+WLA[368] WLA[367] WLA[366] WLA[365] WLA[364] WLA[363] WLA[362] WLA[361] WLA[360] WLA[359]
+WLA[358] WLA[357] WLA[356] WLA[355] WLA[354] WLA[353] WLA[352] WLA[351] WLA[350] WLA[349]
+WLA[348] WLA[347] WLA[346] WLA[345] WLA[344] WLA[343] WLA[342] WLA[341] WLA[340] WLA[339]
+WLA[338] WLA[337] WLA[336] WLA[335] WLA[334] WLA[333] WLA[332] WLA[331] WLA[330] WLA[329]
+WLA[328] WLA[327] WLA[326] WLA[325] WLA[324] WLA[323] WLA[322] WLA[321] WLA[320] WLA[319]
+WLA[318] WLA[317] WLA[316] WLA[315] WLA[314] WLA[313] WLA[312] WLA[311] WLA[310] WLA[309]
+WLA[308] WLA[307] WLA[306] WLA[305] WLA[304] WLA[303] WLA[302] WLA[301] WLA[300] WLA[299]
+WLA[298] WLA[297] WLA[296] WLA[295] WLA[294] WLA[293] WLA[292] WLA[291] WLA[290] WLA[289]
+WLA[288] WLA[287] WLA[286] WLA[285] WLA[284] WLA[283] WLA[282] WLA[281] WLA[280] WLA[279]
+WLA[278] WLA[277] WLA[276] WLA[275] WLA[274] WLA[273] WLA[272] WLA[271] WLA[270] WLA[269]
+WLA[268] WLA[267] WLA[266] WLA[265] WLA[264] WLA[263] WLA[262] WLA[261] WLA[260] WLA[259]
+WLA[258] WLA[257] WLA[256] WLA[255] WLA[254] WLA[253] WLA[252] WLA[251] WLA[250] WLA[249]
+WLA[248] WLA[247] WLA[246] WLA[245] WLA[244] WLA[243] WLA[242] WLA[241] WLA[240] WLA[239]
+WLA[238] WLA[237] WLA[236] WLA[235] WLA[234] WLA[233] WLA[232] WLA[231] WLA[230] WLA[229]
+WLA[228] WLA[227] WLA[226] WLA[225] WLA[224] WLA[223] WLA[222] WLA[221] WLA[220] WLA[219]
+WLA[218] WLA[217] WLA[216] WLA[215] WLA[214] WLA[213] WLA[212] WLA[211] WLA[210] WLA[209]
+WLA[208] WLA[207] WLA[206] WLA[205] WLA[204] WLA[203] WLA[202] WLA[201] WLA[200] WLA[199]
+WLA[198] WLA[197] WLA[196] WLA[195] WLA[194] WLA[193] WLA[192] WLA[191] WLA[190] WLA[189]
+WLA[188] WLA[187] WLA[186] WLA[185] WLA[184] WLA[183] WLA[182] WLA[181] WLA[180] WLA[179]
+WLA[178] WLA[177] WLA[176] WLA[175] WLA[174] WLA[173] WLA[172] WLA[171] WLA[170] WLA[169]
+WLA[168] WLA[167] WLA[166] WLA[165] WLA[164] WLA[163] WLA[162] WLA[161] WLA[160] WLA[159]
+WLA[158] WLA[157] WLA[156] WLA[155] WLA[154] WLA[153] WLA[152] WLA[151] WLA[150] WLA[149]
+WLA[148] WLA[147] WLA[146] WLA[145] WLA[144] WLA[143] WLA[142] WLA[141] WLA[140] WLA[139]
+WLA[138] WLA[137] WLA[136] WLA[135] WLA[134] WLA[133] WLA[132] WLA[131] WLA[130] WLA[129]
+WLA[128] WLA[127] WLA[126] WLA[125] WLA[124] WLA[123] WLA[122] WLA[121] WLA[120] WLA[119]
+WLA[118] WLA[117] WLA[116] WLA[115] WLA[114] WLA[113] WLA[112] WLA[111] WLA[110] WLA[109]
+WLA[108] WLA[107] WLA[106] WLA[105] WLA[104] WLA[103] WLA[102] WLA[101] WLA[100] WLA[99]
+WLA[98] WLA[97] WLA[96] WLA[95] WLA[94] WLA[93] WLA[92] WLA[91] WLA[90] WLA[89]
+WLA[88] WLA[87] WLA[86] WLA[85] WLA[84] WLA[83] WLA[82] WLA[81] WLA[80] WLA[79]
+WLA[78] WLA[77] WLA[76] WLA[75] WLA[74] WLA[73] WLA[72] WLA[71] WLA[70] WLA[69]
+WLA[68] WLA[67] WLA[66] WLA[65] WLA[64] WLA[63] WLA[62] WLA[61] WLA[60] WLA[59]
+WLA[58] WLA[57] WLA[56] WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50] WLA[49]
+WLA[48] WLA[47] WLA[46] WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39]
+WLA[38] WLA[37] WLA[36] WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29]
+WLA[28] WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19]
+WLA[18] WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9]
+WLA[8] WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] WLB[511]
+WLB[510] WLB[509] WLB[508] WLB[507] WLB[506] WLB[505] WLB[504] WLB[503] WLB[502] WLB[501]
+WLB[500] WLB[499] WLB[498] WLB[497] WLB[496] WLB[495] WLB[494] WLB[493] WLB[492] WLB[491]
+WLB[490] WLB[489] WLB[488] WLB[487] WLB[486] WLB[485] WLB[484] WLB[483] WLB[482] WLB[481]
+WLB[480] WLB[479] WLB[478] WLB[477] WLB[476] WLB[475] WLB[474] WLB[473] WLB[472] WLB[471]
+WLB[470] WLB[469] WLB[468] WLB[467] WLB[466] WLB[465] WLB[464] WLB[463] WLB[462] WLB[461]
+WLB[460] WLB[459] WLB[458] WLB[457] WLB[456] WLB[455] WLB[454] WLB[453] WLB[452] WLB[451]
+WLB[450] WLB[449] WLB[448] WLB[447] WLB[446] WLB[445] WLB[444] WLB[443] WLB[442] WLB[441]
+WLB[440] WLB[439] WLB[438] WLB[437] WLB[436] WLB[435] WLB[434] WLB[433] WLB[432] WLB[431]
+WLB[430] WLB[429] WLB[428] WLB[427] WLB[426] WLB[425] WLB[424] WLB[423] WLB[422] WLB[421]
+WLB[420] WLB[419] WLB[418] WLB[417] WLB[416] WLB[415] WLB[414] WLB[413] WLB[412] WLB[411]
+WLB[410] WLB[409] WLB[408] WLB[407] WLB[406] WLB[405] WLB[404] WLB[403] WLB[402] WLB[401]
+WLB[400] WLB[399] WLB[398] WLB[397] WLB[396] WLB[395] WLB[394] WLB[393] WLB[392] WLB[391]
+WLB[390] WLB[389] WLB[388] WLB[387] WLB[386] WLB[385] WLB[384] WLB[383] WLB[382] WLB[381]
+WLB[380] WLB[379] WLB[378] WLB[377] WLB[376] WLB[375] WLB[374] WLB[373] WLB[372] WLB[371]
+WLB[370] WLB[369] WLB[368] WLB[367] WLB[366] WLB[365] WLB[364] WLB[363] WLB[362] WLB[361]
+WLB[360] WLB[359] WLB[358] WLB[357] WLB[356] WLB[355] WLB[354] WLB[353] WLB[352] WLB[351]
+WLB[350] WLB[349] WLB[348] WLB[347] WLB[346] WLB[345] WLB[344] WLB[343] WLB[342] WLB[341]
+WLB[340] WLB[339] WLB[338] WLB[337] WLB[336] WLB[335] WLB[334] WLB[333] WLB[332] WLB[331]
+WLB[330] WLB[329] WLB[328] WLB[327] WLB[326] WLB[325] WLB[324] WLB[323] WLB[322] WLB[321]
+WLB[320] WLB[319] WLB[318] WLB[317] WLB[316] WLB[315] WLB[314] WLB[313] WLB[312] WLB[311]
+WLB[310] WLB[309] WLB[308] WLB[307] WLB[306] WLB[305] WLB[304] WLB[303] WLB[302] WLB[301]
+WLB[300] WLB[299] WLB[298] WLB[297] WLB[296] WLB[295] WLB[294] WLB[293] WLB[292] WLB[291]
+WLB[290] WLB[289] WLB[288] WLB[287] WLB[286] WLB[285] WLB[284] WLB[283] WLB[282] WLB[281]
+WLB[280] WLB[279] WLB[278] WLB[277] WLB[276] WLB[275] WLB[274] WLB[273] WLB[272] WLB[271]
+WLB[270] WLB[269] WLB[268] WLB[267] WLB[266] WLB[265] WLB[264] WLB[263] WLB[262] WLB[261]
+WLB[260] WLB[259] WLB[258] WLB[257] WLB[256] WLB[255] WLB[254] WLB[253] WLB[252] WLB[251]
+WLB[250] WLB[249] WLB[248] WLB[247] WLB[246] WLB[245] WLB[244] WLB[243] WLB[242] WLB[241]
+WLB[240] WLB[239] WLB[238] WLB[237] WLB[236] WLB[235] WLB[234] WLB[233] WLB[232] WLB[231]
+WLB[230] WLB[229] WLB[228] WLB[227] WLB[226] WLB[225] WLB[224] WLB[223] WLB[222] WLB[221]
+WLB[220] WLB[219] WLB[218] WLB[217] WLB[216] WLB[215] WLB[214] WLB[213] WLB[212] WLB[211]
+WLB[210] WLB[209] WLB[208] WLB[207] WLB[206] WLB[205] WLB[204] WLB[203] WLB[202] WLB[201]
+WLB[200] WLB[199] WLB[198] WLB[197] WLB[196] WLB[195] WLB[194] WLB[193] WLB[192] WLB[191]
+WLB[190] WLB[189] WLB[188] WLB[187] WLB[186] WLB[185] WLB[184] WLB[183] WLB[182] WLB[181]
+WLB[180] WLB[179] WLB[178] WLB[177] WLB[176] WLB[175] WLB[174] WLB[173] WLB[172] WLB[171]
+WLB[170] WLB[169] WLB[168] WLB[167] WLB[166] WLB[165] WLB[164] WLB[163] WLB[162] WLB[161]
+WLB[160] WLB[159] WLB[158] WLB[157] WLB[156] WLB[155] WLB[154] WLB[153] WLB[152] WLB[151]
+WLB[150] WLB[149] WLB[148] WLB[147] WLB[146] WLB[145] WLB[144] WLB[143] WLB[142] WLB[141]
+WLB[140] WLB[139] WLB[138] WLB[137] WLB[136] WLB[135] WLB[134] WLB[133] WLB[132] WLB[131]
+WLB[130] WLB[129] WLB[128] WLB[127] WLB[126] WLB[125] WLB[124] WLB[123] WLB[122] WLB[121]
+WLB[120] WLB[119] WLB[118] WLB[117] WLB[116] WLB[115] WLB[114] WLB[113] WLB[112] WLB[111]
+WLB[110] WLB[109] WLB[108] WLB[107] WLB[106] WLB[105] WLB[104] WLB[103] WLB[102] WLB[101]
+WLB[100] WLB[99] WLB[98] WLB[97] WLB[96] WLB[95] WLB[94] WLB[93] WLB[92] WLB[91]
+WLB[90] WLB[89] WLB[88] WLB[87] WLB[86] WLB[85] WLB[84] WLB[83] WLB[82] WLB[81]
+WLB[80] WLB[79] WLB[78] WLB[77] WLB[76] WLB[75] WLB[74] WLB[73] WLB[72] WLB[71]
+WLB[70] WLB[69] WLB[68] WLB[67] WLB[66] WLB[65] WLB[64] WLB[63] WLB[62] WLB[61]
+WLB[60] WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54] WLB[53] WLB[52] WLB[51]
+WLB[50] WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44] WLB[43] WLB[42] WLB[41]
+WLB[40] WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34] WLB[33] WLB[32] WLB[31]
+WLB[30] WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24] WLB[23] WLB[22] WLB[21]
+WLB[20] WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14] WLB[13] WLB[12] WLB[11]
+WLB[10] WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4] WLB[3] WLB[2] WLB[1]
+WLB[0] YXA[7] YXA[6] YXA[5] YXA[4] YXA[3] YXA[2] YXA[1] YXA[0] YXB[7]
+YXB[6] YXB[5] YXB[4] YXB[3] YXB[2] YXB[1] YXB[0]
XI0 RWLA[0] RWLA[1] VDD VSS WLA[63] WLA[62] WLA[61] WLA[60] WLA[59] WLA[58]
+WLA[57] WLA[56] WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48]
+WLA[47] WLA[46] WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38]
+WLA[37] WLA[36] WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28]
+WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18]
+WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8]
+WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] S55NLLGDPH_X512Y8D16_BW_EDGECELL66B_RED_LEFT
XI1 VDD VSS WLA[127] WLA[126] WLA[125] WLA[124] WLA[123] WLA[122] WLA[121] WLA[120]
+WLA[119] WLA[118] WLA[117] WLA[116] WLA[115] WLA[114] WLA[113] WLA[112] WLA[111] WLA[110]
+WLA[109] WLA[108] WLA[107] WLA[106] WLA[105] WLA[104] WLA[103] WLA[102] WLA[101] WLA[100]
+WLA[99] WLA[98] WLA[97] WLA[96] WLA[95] WLA[94] WLA[93] WLA[92] WLA[91] WLA[90]
+WLA[89] WLA[88] WLA[87] WLA[86] WLA[85] WLA[84] WLA[83] WLA[82] WLA[81] WLA[80]
+WLA[79] WLA[78] WLA[77] WLA[76] WLA[75] WLA[74] WLA[73] WLA[72] WLA[71] WLA[70]
+WLA[69] WLA[68] WLA[67] WLA[66] WLA[65] WLA[64] S55NLLGDPH_X512Y8D16_BW_EDGECELL64A_LEFT
XI2 VDD VSS WLA[191] WLA[190] WLA[189] WLA[188] WLA[187] WLA[186] WLA[185] WLA[184]
+WLA[183] WLA[182] WLA[181] WLA[180] WLA[179] WLA[178] WLA[177] WLA[176] WLA[175] WLA[174]
+WLA[173] WLA[172] WLA[171] WLA[170] WLA[169] WLA[168] WLA[167] WLA[166] WLA[165] WLA[164]
+WLA[163] WLA[162] WLA[161] WLA[160] WLA[159] WLA[158] WLA[157] WLA[156] WLA[155] WLA[154]
+WLA[153] WLA[152] WLA[151] WLA[150] WLA[149] WLA[148] WLA[147] WLA[146] WLA[145] WLA[144]
+WLA[143] WLA[142] WLA[141] WLA[140] WLA[139] WLA[138] WLA[137] WLA[136] WLA[135] WLA[134]
+WLA[133] WLA[132] WLA[131] WLA[130] WLA[129] WLA[128] S55NLLGDPH_X512Y8D16_BW_EDGECELL64B_LEFT
XI3 VDD VSS WLA[255] WLA[254] WLA[253] WLA[252] WLA[251] WLA[250] WLA[249] WLA[248]
+WLA[247] WLA[246] WLA[245] WLA[244] WLA[243] WLA[242] WLA[241] WLA[240] WLA[239] WLA[238]
+WLA[237] WLA[236] WLA[235] WLA[234] WLA[233] WLA[232] WLA[231] WLA[230] WLA[229] WLA[228]
+WLA[227] WLA[226] WLA[225] WLA[224] WLA[223] WLA[222] WLA[221] WLA[220] WLA[219] WLA[218]
+WLA[217] WLA[216] WLA[215] WLA[214] WLA[213] WLA[212] WLA[211] WLA[210] WLA[209] WLA[208]
+WLA[207] WLA[206] WLA[205] WLA[204] WLA[203] WLA[202] WLA[201] WLA[200] WLA[199] WLA[198]
+WLA[197] WLA[196] WLA[195] WLA[194] WLA[193] WLA[192] S55NLLGDPH_X512Y8D16_BW_EDGECELL64A_LEFT
XI4 VDD VSS WLA[319] WLA[318] WLA[317] WLA[316] WLA[315] WLA[314] WLA[313] WLA[312]
+WLA[311] WLA[310] WLA[309] WLA[308] WLA[307] WLA[306] WLA[305] WLA[304] WLA[303] WLA[302]
+WLA[301] WLA[300] WLA[299] WLA[298] WLA[297] WLA[296] WLA[295] WLA[294] WLA[293] WLA[292]
+WLA[291] WLA[290] WLA[289] WLA[288] WLA[287] WLA[286] WLA[285] WLA[284] WLA[283] WLA[282]
+WLA[281] WLA[280] WLA[279] WLA[278] WLA[277] WLA[276] WLA[275] WLA[274] WLA[273] WLA[272]
+WLA[271] WLA[270] WLA[269] WLA[268] WLA[267] WLA[266] WLA[265] WLA[264] WLA[263] WLA[262]
+WLA[261] WLA[260] WLA[259] WLA[258] WLA[257] WLA[256] S55NLLGDPH_X512Y8D16_BW_EDGECELL64B_LEFT
XI5 VDD VSS WLA[383] WLA[382] WLA[381] WLA[380] WLA[379] WLA[378] WLA[377] WLA[376]
+WLA[375] WLA[374] WLA[373] WLA[372] WLA[371] WLA[370] WLA[369] WLA[368] WLA[367] WLA[366]
+WLA[365] WLA[364] WLA[363] WLA[362] WLA[361] WLA[360] WLA[359] WLA[358] WLA[357] WLA[356]
+WLA[355] WLA[354] WLA[353] WLA[352] WLA[351] WLA[350] WLA[349] WLA[348] WLA[347] WLA[346]
+WLA[345] WLA[344] WLA[343] WLA[342] WLA[341] WLA[340] WLA[339] WLA[338] WLA[337] WLA[336]
+WLA[335] WLA[334] WLA[333] WLA[332] WLA[331] WLA[330] WLA[329] WLA[328] WLA[327] WLA[326]
+WLA[325] WLA[324] WLA[323] WLA[322] WLA[321] WLA[320] S55NLLGDPH_X512Y8D16_BW_EDGECELL64A_LEFT
XI6 VDD VSS WLA[447] WLA[446] WLA[445] WLA[444] WLA[443] WLA[442] WLA[441] WLA[440]
+WLA[439] WLA[438] WLA[437] WLA[436] WLA[435] WLA[434] WLA[433] WLA[432] WLA[431] WLA[430]
+WLA[429] WLA[428] WLA[427] WLA[426] WLA[425] WLA[424] WLA[423] WLA[422] WLA[421] WLA[420]
+WLA[419] WLA[418] WLA[417] WLA[416] WLA[415] WLA[414] WLA[413] WLA[412] WLA[411] WLA[410]
+WLA[409] WLA[408] WLA[407] WLA[406] WLA[405] WLA[404] WLA[403] WLA[402] WLA[401] WLA[400]
+WLA[399] WLA[398] WLA[397] WLA[396] WLA[395] WLA[394] WLA[393] WLA[392] WLA[391] WLA[390]
+WLA[389] WLA[388] WLA[387] WLA[386] WLA[385] WLA[384] S55NLLGDPH_X512Y8D16_BW_EDGECELL64B_LEFT
XI7 VDD VSS WLA[511] WLA[510] WLA[509] WLA[508] WLA[507] WLA[506] WLA[505] WLA[504]
+WLA[503] WLA[502] WLA[501] WLA[500] WLA[499] WLA[498] WLA[497] WLA[496] WLA[495] WLA[494]
+WLA[493] WLA[492] WLA[491] WLA[490] WLA[489] WLA[488] WLA[487] WLA[486] WLA[485] WLA[484]
+WLA[483] WLA[482] WLA[481] WLA[480] WLA[479] WLA[478] WLA[477] WLA[476] WLA[475] WLA[474]
+WLA[473] WLA[472] WLA[471] WLA[470] WLA[469] WLA[468] WLA[467] WLA[466] WLA[465] WLA[464]
+WLA[463] WLA[462] WLA[461] WLA[460] WLA[459] WLA[458] WLA[457] WLA[456] WLA[455] WLA[454]
+WLA[453] WLA[452] WLA[451] WLA[450] WLA[449] WLA[448] S55NLLGDPH_X512Y8D16_BW_EDGECELL68A_TOP_LEFT
XI8 DBL RWLA[0] RWLA[1] VDD VSS WLA[63] WLA[62] WLA[61] WLA[60] WLA[59]
+WLA[58] WLA[57] WLA[56] WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50] WLA[49]
+WLA[48] WLA[47] WLA[46] WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39]
+WLA[38] WLA[37] WLA[36] WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29]
+WLA[28] WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19]
+WLA[18] WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9]
+WLA[8] WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST66B
XI9 DBL VDD VSS WLA[127] WLA[126] WLA[125] WLA[124] WLA[123] WLA[122] WLA[121]
+WLA[120] WLA[119] WLA[118] WLA[117] WLA[116] WLA[115] WLA[114] WLA[113] WLA[112] WLA[111]
+WLA[110] WLA[109] WLA[108] WLA[107] WLA[106] WLA[105] WLA[104] WLA[103] WLA[102] WLA[101]
+WLA[100] WLA[99] WLA[98] WLA[97] WLA[96] WLA[95] WLA[94] WLA[93] WLA[92] WLA[91]
+WLA[90] WLA[89] WLA[88] WLA[87] WLA[86] WLA[85] WLA[84] WLA[83] WLA[82] WLA[81]
+WLA[80] WLA[79] WLA[78] WLA[77] WLA[76] WLA[75] WLA[74] WLA[73] WLA[72] WLA[71]
+WLA[70] WLA[69] WLA[68] WLA[67] WLA[66] WLA[65] WLA[64] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST64A
XI10 DBL VDD VSS WLA[191] WLA[190] WLA[189] WLA[188] WLA[187] WLA[186] WLA[185]
+WLA[184] WLA[183] WLA[182] WLA[181] WLA[180] WLA[179] WLA[178] WLA[177] WLA[176] WLA[175]
+WLA[174] WLA[173] WLA[172] WLA[171] WLA[170] WLA[169] WLA[168] WLA[167] WLA[166] WLA[165]
+WLA[164] WLA[163] WLA[162] WLA[161] WLA[160] WLA[159] WLA[158] WLA[157] WLA[156] WLA[155]
+WLA[154] WLA[153] WLA[152] WLA[151] WLA[150] WLA[149] WLA[148] WLA[147] WLA[146] WLA[145]
+WLA[144] WLA[143] WLA[142] WLA[141] WLA[140] WLA[139] WLA[138] WLA[137] WLA[136] WLA[135]
+WLA[134] WLA[133] WLA[132] WLA[131] WLA[130] WLA[129] WLA[128] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST64B
XI11 DBL VDD VSS WLA[255] WLA[254] WLA[253] WLA[252] WLA[251] WLA[250] WLA[249]
+WLA[248] WLA[247] WLA[246] WLA[245] WLA[244] WLA[243] WLA[242] WLA[241] WLA[240] WLA[239]
+WLA[238] WLA[237] WLA[236] WLA[235] WLA[234] WLA[233] WLA[232] WLA[231] WLA[230] WLA[229]
+WLA[228] WLA[227] WLA[226] WLA[225] WLA[224] WLA[223] WLA[222] WLA[221] WLA[220] WLA[219]
+WLA[218] WLA[217] WLA[216] WLA[215] WLA[214] WLA[213] WLA[212] WLA[211] WLA[210] WLA[209]
+WLA[208] WLA[207] WLA[206] WLA[205] WLA[204] WLA[203] WLA[202] WLA[201] WLA[200] WLA[199]
+WLA[198] WLA[197] WLA[196] WLA[195] WLA[194] WLA[193] WLA[192] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST64A
XI12 DBL VDD VSS WLA[319] WLA[318] WLA[317] WLA[316] WLA[315] WLA[314] WLA[313]
+WLA[312] WLA[311] WLA[310] WLA[309] WLA[308] WLA[307] WLA[306] WLA[305] WLA[304] WLA[303]
+WLA[302] WLA[301] WLA[300] WLA[299] WLA[298] WLA[297] WLA[296] WLA[295] WLA[294] WLA[293]
+WLA[292] WLA[291] WLA[290] WLA[289] WLA[288] WLA[287] WLA[286] WLA[285] WLA[284] WLA[283]
+WLA[282] WLA[281] WLA[280] WLA[279] WLA[278] WLA[277] WLA[276] WLA[275] WLA[274] WLA[273]
+WLA[272] WLA[271] WLA[270] WLA[269] WLA[268] WLA[267] WLA[266] WLA[265] WLA[264] WLA[263]
+WLA[262] WLA[261] WLA[260] WLA[259] WLA[258] WLA[257] WLA[256] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST64B_TW_LEFT
XI13 DBL VDD VSS WLA[383] WLA[382] WLA[381] WLA[380] WLA[379] WLA[378] WLA[377]
+WLA[376] WLA[375] WLA[374] WLA[373] WLA[372] WLA[371] WLA[370] WLA[369] WLA[368] WLA[367]
+WLA[366] WLA[365] WLA[364] WLA[363] WLA[362] WLA[361] WLA[360] WLA[359] WLA[358] WLA[357]
+WLA[356] WLA[355] WLA[354] WLA[353] WLA[352] WLA[351] WLA[350] WLA[349] WLA[348] WLA[347]
+WLA[346] WLA[345] WLA[344] WLA[343] WLA[342] WLA[341] WLA[340] WLA[339] WLA[338] WLA[337]
+WLA[336] WLA[335] WLA[334] WLA[333] WLA[332] WLA[331] WLA[330] WLA[329] WLA[328] WLA[327]
+WLA[326] WLA[325] WLA[324] WLA[323] WLA[322] WLA[321] WLA[320] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST64A_TW_LEFT
XI14 DBL VDD VSS WLA[447] WLA[446] WLA[445] WLA[444] WLA[443] WLA[442] WLA[441]
+WLA[440] WLA[439] WLA[438] WLA[437] WLA[436] WLA[435] WLA[434] WLA[433] WLA[432] WLA[431]
+WLA[430] WLA[429] WLA[428] WLA[427] WLA[426] WLA[425] WLA[424] WLA[423] WLA[422] WLA[421]
+WLA[420] WLA[419] WLA[418] WLA[417] WLA[416] WLA[415] WLA[414] WLA[413] WLA[412] WLA[411]
+WLA[410] WLA[409] WLA[408] WLA[407] WLA[406] WLA[405] WLA[404] WLA[403] WLA[402] WLA[401]
+WLA[400] WLA[399] WLA[398] WLA[397] WLA[396] WLA[395] WLA[394] WLA[393] WLA[392] WLA[391]
+WLA[390] WLA[389] WLA[388] WLA[387] WLA[386] WLA[385] WLA[384] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST64B_TW_LEFT
XI15 DBL STWLA VDD VSS WLA[511] WLA[510] WLA[509] WLA[508] WLA[507] WLA[506]
+WLA[505] WLA[504] WLA[503] WLA[502] WLA[501] WLA[500] WLA[499] WLA[498] WLA[497] WLA[496]
+WLA[495] WLA[494] WLA[493] WLA[492] WLA[491] WLA[490] WLA[489] WLA[488] WLA[487] WLA[486]
+WLA[485] WLA[484] WLA[483] WLA[482] WLA[481] WLA[480] WLA[479] WLA[478] WLA[477] WLA[476]
+WLA[475] WLA[474] WLA[473] WLA[472] WLA[471] WLA[470] WLA[469] WLA[468] WLA[467] WLA[466]
+WLA[465] WLA[464] WLA[463] WLA[462] WLA[461] WLA[460] WLA[459] WLA[458] WLA[457] WLA[456]
+WLA[455] WLA[454] WLA[453] WLA[452] WLA[451] WLA[450] WLA[449] WLA[448] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST68A_TOP_TW_LEFT
XI16 BWENA[0] BWENB[0] CLKA CLKB CLKXA CLKXB DATAA[0] DATAB[0] DOUTA[0] DOUTB[0]
+VSS STWLA STWLA VSS STWLB VSS VSS VSS RWLA[0] RWLA[1]
+RWLB[0] RWLB[1] SACK1A SACK1B SACK4A SACK4B VDD VSS WEA WEB
+WLA[511] WLA[510] WLA[509] WLA[508] WLA[507] WLA[506] WLA[505] WLA[504] WLA[503] WLA[502]
+WLA[501] WLA[500] WLA[499] WLA[498] WLA[497] WLA[496] WLA[495] WLA[494] WLA[493] WLA[492]
+WLA[491] WLA[490] WLA[489] WLA[488] WLA[487] WLA[486] WLA[485] WLA[484] WLA[483] WLA[482]
+WLA[481] WLA[480] WLA[479] WLA[478] WLA[477] WLA[476] WLA[475] WLA[474] WLA[473] WLA[472]
+WLA[471] WLA[470] WLA[469] WLA[468] WLA[467] WLA[466] WLA[465] WLA[464] WLA[463] WLA[462]
+WLA[461] WLA[460] WLA[459] WLA[458] WLA[457] WLA[456] WLA[455] WLA[454] WLA[453] WLA[452]
+WLA[451] WLA[450] WLA[449] WLA[448] WLA[447] WLA[446] WLA[445] WLA[444] WLA[443] WLA[442]
+WLA[441] WLA[440] WLA[439] WLA[438] WLA[437] WLA[436] WLA[435] WLA[434] WLA[433] WLA[432]
+WLA[431] WLA[430] WLA[429] WLA[428] WLA[427] WLA[426] WLA[425] WLA[424] WLA[423] WLA[422]
+WLA[421] WLA[420] WLA[419] WLA[418] WLA[417] WLA[416] WLA[415] WLA[414] WLA[413] WLA[412]
+WLA[411] WLA[410] WLA[409] WLA[408] WLA[407] WLA[406] WLA[405] WLA[404] WLA[403] WLA[402]
+WLA[401] WLA[400] WLA[399] WLA[398] WLA[397] WLA[396] WLA[395] WLA[394] WLA[393] WLA[392]
+WLA[391] WLA[390] WLA[389] WLA[388] WLA[387] WLA[386] WLA[385] WLA[384] WLA[383] WLA[382]
+WLA[381] WLA[380] WLA[379] WLA[378] WLA[377] WLA[376] WLA[375] WLA[374] WLA[373] WLA[372]
+WLA[371] WLA[370] WLA[369] WLA[368] WLA[367] WLA[366] WLA[365] WLA[364] WLA[363] WLA[362]
+WLA[361] WLA[360] WLA[359] WLA[358] WLA[357] WLA[356] WLA[355] WLA[354] WLA[353] WLA[352]
+WLA[351] WLA[350] WLA[349] WLA[348] WLA[347] WLA[346] WLA[345] WLA[344] WLA[343] WLA[342]
+WLA[341] WLA[340] WLA[339] WLA[338] WLA[337] WLA[336] WLA[335] WLA[334] WLA[333] WLA[332]
+WLA[331] WLA[330] WLA[329] WLA[328] WLA[327] WLA[326] WLA[325] WLA[324] WLA[323] WLA[322]
+WLA[321] WLA[320] WLA[319] WLA[318] WLA[317] WLA[316] WLA[315] WLA[314] WLA[313] WLA[312]
+WLA[311] WLA[310] WLA[309] WLA[308] WLA[307] WLA[306] WLA[305] WLA[304] WLA[303] WLA[302]
+WLA[301] WLA[300] WLA[299] WLA[298] WLA[297] WLA[296] WLA[295] WLA[294] WLA[293] WLA[292]
+WLA[291] WLA[290] WLA[289] WLA[288] WLA[287] WLA[286] WLA[285] WLA[284] WLA[283] WLA[282]
+WLA[281] WLA[280] WLA[279] WLA[278] WLA[277] WLA[276] WLA[275] WLA[274] WLA[273] WLA[272]
+WLA[271] WLA[270] WLA[269] WLA[268] WLA[267] WLA[266] WLA[265] WLA[264] WLA[263] WLA[262]
+WLA[261] WLA[260] WLA[259] WLA[258] WLA[257] WLA[256] WLA[255] WLA[254] WLA[253] WLA[252]
+WLA[251] WLA[250] WLA[249] WLA[248] WLA[247] WLA[246] WLA[245] WLA[244] WLA[243] WLA[242]
+WLA[241] WLA[240] WLA[239] WLA[238] WLA[237] WLA[236] WLA[235] WLA[234] WLA[233] WLA[232]
+WLA[231] WLA[230] WLA[229] WLA[228] WLA[227] WLA[226] WLA[225] WLA[224] WLA[223] WLA[222]
+WLA[221] WLA[220] WLA[219] WLA[218] WLA[217] WLA[216] WLA[215] WLA[214] WLA[213] WLA[212]
+WLA[211] WLA[210] WLA[209] WLA[208] WLA[207] WLA[206] WLA[205] WLA[204] WLA[203] WLA[202]
+WLA[201] WLA[200] WLA[199] WLA[198] WLA[197] WLA[196] WLA[195] WLA[194] WLA[193] WLA[192]
+WLA[191] WLA[190] WLA[189] WLA[188] WLA[187] WLA[186] WLA[185] WLA[184] WLA[183] WLA[182]
+WLA[181] WLA[180] WLA[179] WLA[178] WLA[177] WLA[176] WLA[175] WLA[174] WLA[173] WLA[172]
+WLA[171] WLA[170] WLA[169] WLA[168] WLA[167] WLA[166] WLA[165] WLA[164] WLA[163] WLA[162]
+WLA[161] WLA[160] WLA[159] WLA[158] WLA[157] WLA[156] WLA[155] WLA[154] WLA[153] WLA[152]
+WLA[151] WLA[150] WLA[149] WLA[148] WLA[147] WLA[146] WLA[145] WLA[144] WLA[143] WLA[142]
+WLA[141] WLA[140] WLA[139] WLA[138] WLA[137] WLA[136] WLA[135] WLA[134] WLA[133] WLA[132]
+WLA[131] WLA[130] WLA[129] WLA[128] WLA[127] WLA[126] WLA[125] WLA[124] WLA[123] WLA[122]
+WLA[121] WLA[120] WLA[119] WLA[118] WLA[117] WLA[116] WLA[115] WLA[114] WLA[113] WLA[112]
+WLA[111] WLA[110] WLA[109] WLA[108] WLA[107] WLA[106] WLA[105] WLA[104] WLA[103] WLA[102]
+WLA[101] WLA[100] WLA[99] WLA[98] WLA[97] WLA[96] WLA[95] WLA[94] WLA[93] WLA[92]
+WLA[91] WLA[90] WLA[89] WLA[88] WLA[87] WLA[86] WLA[85] WLA[84] WLA[83] WLA[82]
+WLA[81] WLA[80] WLA[79] WLA[78] WLA[77] WLA[76] WLA[75] WLA[74] WLA[73] WLA[72]
+WLA[71] WLA[70] WLA[69] WLA[68] WLA[67] WLA[66] WLA[65] WLA[64] WLA[63] WLA[62]
+WLA[61] WLA[60] WLA[59] WLA[58] WLA[57] WLA[56] WLA[55] WLA[54] WLA[53] WLA[52]
+WLA[51] WLA[50] WLA[49] WLA[48] WLA[47] WLA[46] WLA[45] WLA[44] WLA[43] WLA[42]
+WLA[41] WLA[40] WLA[39] WLA[38] WLA[37] WLA[36] WLA[35] WLA[34] WLA[33] WLA[32]
+WLA[31] WLA[30] WLA[29] WLA[28] WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22]
+WLA[21] WLA[20] WLA[19] WLA[18] WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12]
+WLA[11] WLA[10] WLA[9] WLA[8] WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2]
+WLA[1] WLA[0] WLB[511] WLB[510] WLB[509] WLB[508] WLB[507] WLB[506] WLB[505] WLB[504]
+WLB[503] WLB[502] WLB[501] WLB[500] WLB[499] WLB[498] WLB[497] WLB[496] WLB[495] WLB[494]
+WLB[493] WLB[492] WLB[491] WLB[490] WLB[489] WLB[488] WLB[487] WLB[486] WLB[485] WLB[484]
+WLB[483] WLB[482] WLB[481] WLB[480] WLB[479] WLB[478] WLB[477] WLB[476] WLB[475] WLB[474]
+WLB[473] WLB[472] WLB[471] WLB[470] WLB[469] WLB[468] WLB[467] WLB[466] WLB[465] WLB[464]
+WLB[463] WLB[462] WLB[461] WLB[460] WLB[459] WLB[458] WLB[457] WLB[456] WLB[455] WLB[454]
+WLB[453] WLB[452] WLB[451] WLB[450] WLB[449] WLB[448] WLB[447] WLB[446] WLB[445] WLB[444]
+WLB[443] WLB[442] WLB[441] WLB[440] WLB[439] WLB[438] WLB[437] WLB[436] WLB[435] WLB[434]
+WLB[433] WLB[432] WLB[431] WLB[430] WLB[429] WLB[428] WLB[427] WLB[426] WLB[425] WLB[424]
+WLB[423] WLB[422] WLB[421] WLB[420] WLB[419] WLB[418] WLB[417] WLB[416] WLB[415] WLB[414]
+WLB[413] WLB[412] WLB[411] WLB[410] WLB[409] WLB[408] WLB[407] WLB[406] WLB[405] WLB[404]
+WLB[403] WLB[402] WLB[401] WLB[400] WLB[399] WLB[398] WLB[397] WLB[396] WLB[395] WLB[394]
+WLB[393] WLB[392] WLB[391] WLB[390] WLB[389] WLB[388] WLB[387] WLB[386] WLB[385] WLB[384]
+WLB[383] WLB[382] WLB[381] WLB[380] WLB[379] WLB[378] WLB[377] WLB[376] WLB[375] WLB[374]
+WLB[373] WLB[372] WLB[371] WLB[370] WLB[369] WLB[368] WLB[367] WLB[366] WLB[365] WLB[364]
+WLB[363] WLB[362] WLB[361] WLB[360] WLB[359] WLB[358] WLB[357] WLB[356] WLB[355] WLB[354]
+WLB[353] WLB[352] WLB[351] WLB[350] WLB[349] WLB[348] WLB[347] WLB[346] WLB[345] WLB[344]
+WLB[343] WLB[342] WLB[341] WLB[340] WLB[339] WLB[338] WLB[337] WLB[336] WLB[335] WLB[334]
+WLB[333] WLB[332] WLB[331] WLB[330] WLB[329] WLB[328] WLB[327] WLB[326] WLB[325] WLB[324]
+WLB[323] WLB[322] WLB[321] WLB[320] WLB[319] WLB[318] WLB[317] WLB[316] WLB[315] WLB[314]
+WLB[313] WLB[312] WLB[311] WLB[310] WLB[309] WLB[308] WLB[307] WLB[306] WLB[305] WLB[304]
+WLB[303] WLB[302] WLB[301] WLB[300] WLB[299] WLB[298] WLB[297] WLB[296] WLB[295] WLB[294]
+WLB[293] WLB[292] WLB[291] WLB[290] WLB[289] WLB[288] WLB[287] WLB[286] WLB[285] WLB[284]
+WLB[283] WLB[282] WLB[281] WLB[280] WLB[279] WLB[278] WLB[277] WLB[276] WLB[275] WLB[274]
+WLB[273] WLB[272] WLB[271] WLB[270] WLB[269] WLB[268] WLB[267] WLB[266] WLB[265] WLB[264]
+WLB[263] WLB[262] WLB[261] WLB[260] WLB[259] WLB[258] WLB[257] WLB[256] WLB[255] WLB[254]
+WLB[253] WLB[252] WLB[251] WLB[250] WLB[249] WLB[248] WLB[247] WLB[246] WLB[245] WLB[244]
+WLB[243] WLB[242] WLB[241] WLB[240] WLB[239] WLB[238] WLB[237] WLB[236] WLB[235] WLB[234]
+WLB[233] WLB[232] WLB[231] WLB[230] WLB[229] WLB[228] WLB[227] WLB[226] WLB[225] WLB[224]
+WLB[223] WLB[222] WLB[221] WLB[220] WLB[219] WLB[218] WLB[217] WLB[216] WLB[215] WLB[214]
+WLB[213] WLB[212] WLB[211] WLB[210] WLB[209] WLB[208] WLB[207] WLB[206] WLB[205] WLB[204]
+WLB[203] WLB[202] WLB[201] WLB[200] WLB[199] WLB[198] WLB[197] WLB[196] WLB[195] WLB[194]
+WLB[193] WLB[192] WLB[191] WLB[190] WLB[189] WLB[188] WLB[187] WLB[186] WLB[185] WLB[184]
+WLB[183] WLB[182] WLB[181] WLB[180] WLB[179] WLB[178] WLB[177] WLB[176] WLB[175] WLB[174]
+WLB[173] WLB[172] WLB[171] WLB[170] WLB[169] WLB[168] WLB[167] WLB[166] WLB[165] WLB[164]
+WLB[163] WLB[162] WLB[161] WLB[160] WLB[159] WLB[158] WLB[157] WLB[156] WLB[155] WLB[154]
+WLB[153] WLB[152] WLB[151] WLB[150] WLB[149] WLB[148] WLB[147] WLB[146] WLB[145] WLB[144]
+WLB[143] WLB[142] WLB[141] WLB[140] WLB[139] WLB[138] WLB[137] WLB[136] WLB[135] WLB[134]
+WLB[133] WLB[132] WLB[131] WLB[130] WLB[129] WLB[128] WLB[127] WLB[126] WLB[125] WLB[124]
+WLB[123] WLB[122] WLB[121] WLB[120] WLB[119] WLB[118] WLB[117] WLB[116] WLB[115] WLB[114]
+WLB[113] WLB[112] WLB[111] WLB[110] WLB[109] WLB[108] WLB[107] WLB[106] WLB[105] WLB[104]
+WLB[103] WLB[102] WLB[101] WLB[100] WLB[99] WLB[98] WLB[97] WLB[96] WLB[95] WLB[94]
+WLB[93] WLB[92] WLB[91] WLB[90] WLB[89] WLB[88] WLB[87] WLB[86] WLB[85] WLB[84]
+WLB[83] WLB[82] WLB[81] WLB[80] WLB[79] WLB[78] WLB[77] WLB[76] WLB[75] WLB[74]
+WLB[73] WLB[72] WLB[71] WLB[70] WLB[69] WLB[68] WLB[67] WLB[66] WLB[65] WLB[64]
+WLB[63] WLB[62] WLB[61] WLB[60] WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54]
+WLB[53] WLB[52] WLB[51] WLB[50] WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44]
+WLB[43] WLB[42] WLB[41] WLB[40] WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34]
+WLB[33] WLB[32] WLB[31] WLB[30] WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24]
+WLB[23] WLB[22] WLB[21] WLB[20] WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14]
+WLB[13] WLB[12] WLB[11] WLB[10] WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4]
+WLB[3] WLB[2] WLB[1] WLB[0] YXA[7] YXA[6] YXA[5] YXA[4] YXA[3] YXA[2]
+YXA[1] YXA[0] YXB[7] YXB[6] YXB[5] YXB[4] YXB[3] YXB[2] YXB[1] YXB[0] S55NLLGDPH_X512Y8D16_BW_Y512X8CELL_BW
XI17 BWENA[1] BWENB[1] CLKA CLKB CLKXA CLKXB DATAA[1] DATAB[1] DOUTA[1] DOUTB[1]
+VSS STWLA STWLA VSS STWLB VSS VSS VSS RWLA[0] RWLA[1]
+RWLB[0] RWLB[1] SACK1A SACK1B SACK4A SACK4B VDD VSS WEA WEB
+WLA[511] WLA[510] WLA[509] WLA[508] WLA[507] WLA[506] WLA[505] WLA[504] WLA[503] WLA[502]
+WLA[501] WLA[500] WLA[499] WLA[498] WLA[497] WLA[496] WLA[495] WLA[494] WLA[493] WLA[492]
+WLA[491] WLA[490] WLA[489] WLA[488] WLA[487] WLA[486] WLA[485] WLA[484] WLA[483] WLA[482]
+WLA[481] WLA[480] WLA[479] WLA[478] WLA[477] WLA[476] WLA[475] WLA[474] WLA[473] WLA[472]
+WLA[471] WLA[470] WLA[469] WLA[468] WLA[467] WLA[466] WLA[465] WLA[464] WLA[463] WLA[462]
+WLA[461] WLA[460] WLA[459] WLA[458] WLA[457] WLA[456] WLA[455] WLA[454] WLA[453] WLA[452]
+WLA[451] WLA[450] WLA[449] WLA[448] WLA[447] WLA[446] WLA[445] WLA[444] WLA[443] WLA[442]
+WLA[441] WLA[440] WLA[439] WLA[438] WLA[437] WLA[436] WLA[435] WLA[434] WLA[433] WLA[432]
+WLA[431] WLA[430] WLA[429] WLA[428] WLA[427] WLA[426] WLA[425] WLA[424] WLA[423] WLA[422]
+WLA[421] WLA[420] WLA[419] WLA[418] WLA[417] WLA[416] WLA[415] WLA[414] WLA[413] WLA[412]
+WLA[411] WLA[410] WLA[409] WLA[408] WLA[407] WLA[406] WLA[405] WLA[404] WLA[403] WLA[402]
+WLA[401] WLA[400] WLA[399] WLA[398] WLA[397] WLA[396] WLA[395] WLA[394] WLA[393] WLA[392]
+WLA[391] WLA[390] WLA[389] WLA[388] WLA[387] WLA[386] WLA[385] WLA[384] WLA[383] WLA[382]
+WLA[381] WLA[380] WLA[379] WLA[378] WLA[377] WLA[376] WLA[375] WLA[374] WLA[373] WLA[372]
+WLA[371] WLA[370] WLA[369] WLA[368] WLA[367] WLA[366] WLA[365] WLA[364] WLA[363] WLA[362]
+WLA[361] WLA[360] WLA[359] WLA[358] WLA[357] WLA[356] WLA[355] WLA[354] WLA[353] WLA[352]
+WLA[351] WLA[350] WLA[349] WLA[348] WLA[347] WLA[346] WLA[345] WLA[344] WLA[343] WLA[342]
+WLA[341] WLA[340] WLA[339] WLA[338] WLA[337] WLA[336] WLA[335] WLA[334] WLA[333] WLA[332]
+WLA[331] WLA[330] WLA[329] WLA[328] WLA[327] WLA[326] WLA[325] WLA[324] WLA[323] WLA[322]
+WLA[321] WLA[320] WLA[319] WLA[318] WLA[317] WLA[316] WLA[315] WLA[314] WLA[313] WLA[312]
+WLA[311] WLA[310] WLA[309] WLA[308] WLA[307] WLA[306] WLA[305] WLA[304] WLA[303] WLA[302]
+WLA[301] WLA[300] WLA[299] WLA[298] WLA[297] WLA[296] WLA[295] WLA[294] WLA[293] WLA[292]
+WLA[291] WLA[290] WLA[289] WLA[288] WLA[287] WLA[286] WLA[285] WLA[284] WLA[283] WLA[282]
+WLA[281] WLA[280] WLA[279] WLA[278] WLA[277] WLA[276] WLA[275] WLA[274] WLA[273] WLA[272]
+WLA[271] WLA[270] WLA[269] WLA[268] WLA[267] WLA[266] WLA[265] WLA[264] WLA[263] WLA[262]
+WLA[261] WLA[260] WLA[259] WLA[258] WLA[257] WLA[256] WLA[255] WLA[254] WLA[253] WLA[252]
+WLA[251] WLA[250] WLA[249] WLA[248] WLA[247] WLA[246] WLA[245] WLA[244] WLA[243] WLA[242]
+WLA[241] WLA[240] WLA[239] WLA[238] WLA[237] WLA[236] WLA[235] WLA[234] WLA[233] WLA[232]
+WLA[231] WLA[230] WLA[229] WLA[228] WLA[227] WLA[226] WLA[225] WLA[224] WLA[223] WLA[222]
+WLA[221] WLA[220] WLA[219] WLA[218] WLA[217] WLA[216] WLA[215] WLA[214] WLA[213] WLA[212]
+WLA[211] WLA[210] WLA[209] WLA[208] WLA[207] WLA[206] WLA[205] WLA[204] WLA[203] WLA[202]
+WLA[201] WLA[200] WLA[199] WLA[198] WLA[197] WLA[196] WLA[195] WLA[194] WLA[193] WLA[192]
+WLA[191] WLA[190] WLA[189] WLA[188] WLA[187] WLA[186] WLA[185] WLA[184] WLA[183] WLA[182]
+WLA[181] WLA[180] WLA[179] WLA[178] WLA[177] WLA[176] WLA[175] WLA[174] WLA[173] WLA[172]
+WLA[171] WLA[170] WLA[169] WLA[168] WLA[167] WLA[166] WLA[165] WLA[164] WLA[163] WLA[162]
+WLA[161] WLA[160] WLA[159] WLA[158] WLA[157] WLA[156] WLA[155] WLA[154] WLA[153] WLA[152]
+WLA[151] WLA[150] WLA[149] WLA[148] WLA[147] WLA[146] WLA[145] WLA[144] WLA[143] WLA[142]
+WLA[141] WLA[140] WLA[139] WLA[138] WLA[137] WLA[136] WLA[135] WLA[134] WLA[133] WLA[132]
+WLA[131] WLA[130] WLA[129] WLA[128] WLA[127] WLA[126] WLA[125] WLA[124] WLA[123] WLA[122]
+WLA[121] WLA[120] WLA[119] WLA[118] WLA[117] WLA[116] WLA[115] WLA[114] WLA[113] WLA[112]
+WLA[111] WLA[110] WLA[109] WLA[108] WLA[107] WLA[106] WLA[105] WLA[104] WLA[103] WLA[102]
+WLA[101] WLA[100] WLA[99] WLA[98] WLA[97] WLA[96] WLA[95] WLA[94] WLA[93] WLA[92]
+WLA[91] WLA[90] WLA[89] WLA[88] WLA[87] WLA[86] WLA[85] WLA[84] WLA[83] WLA[82]
+WLA[81] WLA[80] WLA[79] WLA[78] WLA[77] WLA[76] WLA[75] WLA[74] WLA[73] WLA[72]
+WLA[71] WLA[70] WLA[69] WLA[68] WLA[67] WLA[66] WLA[65] WLA[64] WLA[63] WLA[62]
+WLA[61] WLA[60] WLA[59] WLA[58] WLA[57] WLA[56] WLA[55] WLA[54] WLA[53] WLA[52]
+WLA[51] WLA[50] WLA[49] WLA[48] WLA[47] WLA[46] WLA[45] WLA[44] WLA[43] WLA[42]
+WLA[41] WLA[40] WLA[39] WLA[38] WLA[37] WLA[36] WLA[35] WLA[34] WLA[33] WLA[32]
+WLA[31] WLA[30] WLA[29] WLA[28] WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22]
+WLA[21] WLA[20] WLA[19] WLA[18] WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12]
+WLA[11] WLA[10] WLA[9] WLA[8] WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2]
+WLA[1] WLA[0] WLB[511] WLB[510] WLB[509] WLB[508] WLB[507] WLB[506] WLB[505] WLB[504]
+WLB[503] WLB[502] WLB[501] WLB[500] WLB[499] WLB[498] WLB[497] WLB[496] WLB[495] WLB[494]
+WLB[493] WLB[492] WLB[491] WLB[490] WLB[489] WLB[488] WLB[487] WLB[486] WLB[485] WLB[484]
+WLB[483] WLB[482] WLB[481] WLB[480] WLB[479] WLB[478] WLB[477] WLB[476] WLB[475] WLB[474]
+WLB[473] WLB[472] WLB[471] WLB[470] WLB[469] WLB[468] WLB[467] WLB[466] WLB[465] WLB[464]
+WLB[463] WLB[462] WLB[461] WLB[460] WLB[459] WLB[458] WLB[457] WLB[456] WLB[455] WLB[454]
+WLB[453] WLB[452] WLB[451] WLB[450] WLB[449] WLB[448] WLB[447] WLB[446] WLB[445] WLB[444]
+WLB[443] WLB[442] WLB[441] WLB[440] WLB[439] WLB[438] WLB[437] WLB[436] WLB[435] WLB[434]
+WLB[433] WLB[432] WLB[431] WLB[430] WLB[429] WLB[428] WLB[427] WLB[426] WLB[425] WLB[424]
+WLB[423] WLB[422] WLB[421] WLB[420] WLB[419] WLB[418] WLB[417] WLB[416] WLB[415] WLB[414]
+WLB[413] WLB[412] WLB[411] WLB[410] WLB[409] WLB[408] WLB[407] WLB[406] WLB[405] WLB[404]
+WLB[403] WLB[402] WLB[401] WLB[400] WLB[399] WLB[398] WLB[397] WLB[396] WLB[395] WLB[394]
+WLB[393] WLB[392] WLB[391] WLB[390] WLB[389] WLB[388] WLB[387] WLB[386] WLB[385] WLB[384]
+WLB[383] WLB[382] WLB[381] WLB[380] WLB[379] WLB[378] WLB[377] WLB[376] WLB[375] WLB[374]
+WLB[373] WLB[372] WLB[371] WLB[370] WLB[369] WLB[368] WLB[367] WLB[366] WLB[365] WLB[364]
+WLB[363] WLB[362] WLB[361] WLB[360] WLB[359] WLB[358] WLB[357] WLB[356] WLB[355] WLB[354]
+WLB[353] WLB[352] WLB[351] WLB[350] WLB[349] WLB[348] WLB[347] WLB[346] WLB[345] WLB[344]
+WLB[343] WLB[342] WLB[341] WLB[340] WLB[339] WLB[338] WLB[337] WLB[336] WLB[335] WLB[334]
+WLB[333] WLB[332] WLB[331] WLB[330] WLB[329] WLB[328] WLB[327] WLB[326] WLB[325] WLB[324]
+WLB[323] WLB[322] WLB[321] WLB[320] WLB[319] WLB[318] WLB[317] WLB[316] WLB[315] WLB[314]
+WLB[313] WLB[312] WLB[311] WLB[310] WLB[309] WLB[308] WLB[307] WLB[306] WLB[305] WLB[304]
+WLB[303] WLB[302] WLB[301] WLB[300] WLB[299] WLB[298] WLB[297] WLB[296] WLB[295] WLB[294]
+WLB[293] WLB[292] WLB[291] WLB[290] WLB[289] WLB[288] WLB[287] WLB[286] WLB[285] WLB[284]
+WLB[283] WLB[282] WLB[281] WLB[280] WLB[279] WLB[278] WLB[277] WLB[276] WLB[275] WLB[274]
+WLB[273] WLB[272] WLB[271] WLB[270] WLB[269] WLB[268] WLB[267] WLB[266] WLB[265] WLB[264]
+WLB[263] WLB[262] WLB[261] WLB[260] WLB[259] WLB[258] WLB[257] WLB[256] WLB[255] WLB[254]
+WLB[253] WLB[252] WLB[251] WLB[250] WLB[249] WLB[248] WLB[247] WLB[246] WLB[245] WLB[244]
+WLB[243] WLB[242] WLB[241] WLB[240] WLB[239] WLB[238] WLB[237] WLB[236] WLB[235] WLB[234]
+WLB[233] WLB[232] WLB[231] WLB[230] WLB[229] WLB[228] WLB[227] WLB[226] WLB[225] WLB[224]
+WLB[223] WLB[222] WLB[221] WLB[220] WLB[219] WLB[218] WLB[217] WLB[216] WLB[215] WLB[214]
+WLB[213] WLB[212] WLB[211] WLB[210] WLB[209] WLB[208] WLB[207] WLB[206] WLB[205] WLB[204]
+WLB[203] WLB[202] WLB[201] WLB[200] WLB[199] WLB[198] WLB[197] WLB[196] WLB[195] WLB[194]
+WLB[193] WLB[192] WLB[191] WLB[190] WLB[189] WLB[188] WLB[187] WLB[186] WLB[185] WLB[184]
+WLB[183] WLB[182] WLB[181] WLB[180] WLB[179] WLB[178] WLB[177] WLB[176] WLB[175] WLB[174]
+WLB[173] WLB[172] WLB[171] WLB[170] WLB[169] WLB[168] WLB[167] WLB[166] WLB[165] WLB[164]
+WLB[163] WLB[162] WLB[161] WLB[160] WLB[159] WLB[158] WLB[157] WLB[156] WLB[155] WLB[154]
+WLB[153] WLB[152] WLB[151] WLB[150] WLB[149] WLB[148] WLB[147] WLB[146] WLB[145] WLB[144]
+WLB[143] WLB[142] WLB[141] WLB[140] WLB[139] WLB[138] WLB[137] WLB[136] WLB[135] WLB[134]
+WLB[133] WLB[132] WLB[131] WLB[130] WLB[129] WLB[128] WLB[127] WLB[126] WLB[125] WLB[124]
+WLB[123] WLB[122] WLB[121] WLB[120] WLB[119] WLB[118] WLB[117] WLB[116] WLB[115] WLB[114]
+WLB[113] WLB[112] WLB[111] WLB[110] WLB[109] WLB[108] WLB[107] WLB[106] WLB[105] WLB[104]
+WLB[103] WLB[102] WLB[101] WLB[100] WLB[99] WLB[98] WLB[97] WLB[96] WLB[95] WLB[94]
+WLB[93] WLB[92] WLB[91] WLB[90] WLB[89] WLB[88] WLB[87] WLB[86] WLB[85] WLB[84]
+WLB[83] WLB[82] WLB[81] WLB[80] WLB[79] WLB[78] WLB[77] WLB[76] WLB[75] WLB[74]
+WLB[73] WLB[72] WLB[71] WLB[70] WLB[69] WLB[68] WLB[67] WLB[66] WLB[65] WLB[64]
+WLB[63] WLB[62] WLB[61] WLB[60] WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54]
+WLB[53] WLB[52] WLB[51] WLB[50] WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44]
+WLB[43] WLB[42] WLB[41] WLB[40] WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34]
+WLB[33] WLB[32] WLB[31] WLB[30] WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24]
+WLB[23] WLB[22] WLB[21] WLB[20] WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14]
+WLB[13] WLB[12] WLB[11] WLB[10] WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4]
+WLB[3] WLB[2] WLB[1] WLB[0] YXA[7] YXA[6] YXA[5] YXA[4] YXA[3] YXA[2]
+YXA[1] YXA[0] YXB[7] YXB[6] YXB[5] YXB[4] YXB[3] YXB[2] YXB[1] YXB[0] S55NLLGDPH_X512Y8D16_BW_Y512X8CELL_BW
XI18 BWENA[2] BWENB[2] CLKA CLKB CLKXA CLKXB DATAA[2] DATAB[2] DOUTA[2] DOUTB[2]
+VSS STWLA STWLA VSS STWLB VSS VSS VSS RWLA[0] RWLA[1]
+RWLB[0] RWLB[1] SACK1A SACK1B SACK4A SACK4B VDD VSS WEA WEB
+WLA[511] WLA[510] WLA[509] WLA[508] WLA[507] WLA[506] WLA[505] WLA[504] WLA[503] WLA[502]
+WLA[501] WLA[500] WLA[499] WLA[498] WLA[497] WLA[496] WLA[495] WLA[494] WLA[493] WLA[492]
+WLA[491] WLA[490] WLA[489] WLA[488] WLA[487] WLA[486] WLA[485] WLA[484] WLA[483] WLA[482]
+WLA[481] WLA[480] WLA[479] WLA[478] WLA[477] WLA[476] WLA[475] WLA[474] WLA[473] WLA[472]
+WLA[471] WLA[470] WLA[469] WLA[468] WLA[467] WLA[466] WLA[465] WLA[464] WLA[463] WLA[462]
+WLA[461] WLA[460] WLA[459] WLA[458] WLA[457] WLA[456] WLA[455] WLA[454] WLA[453] WLA[452]
+WLA[451] WLA[450] WLA[449] WLA[448] WLA[447] WLA[446] WLA[445] WLA[444] WLA[443] WLA[442]
+WLA[441] WLA[440] WLA[439] WLA[438] WLA[437] WLA[436] WLA[435] WLA[434] WLA[433] WLA[432]
+WLA[431] WLA[430] WLA[429] WLA[428] WLA[427] WLA[426] WLA[425] WLA[424] WLA[423] WLA[422]
+WLA[421] WLA[420] WLA[419] WLA[418] WLA[417] WLA[416] WLA[415] WLA[414] WLA[413] WLA[412]
+WLA[411] WLA[410] WLA[409] WLA[408] WLA[407] WLA[406] WLA[405] WLA[404] WLA[403] WLA[402]
+WLA[401] WLA[400] WLA[399] WLA[398] WLA[397] WLA[396] WLA[395] WLA[394] WLA[393] WLA[392]
+WLA[391] WLA[390] WLA[389] WLA[388] WLA[387] WLA[386] WLA[385] WLA[384] WLA[383] WLA[382]
+WLA[381] WLA[380] WLA[379] WLA[378] WLA[377] WLA[376] WLA[375] WLA[374] WLA[373] WLA[372]
+WLA[371] WLA[370] WLA[369] WLA[368] WLA[367] WLA[366] WLA[365] WLA[364] WLA[363] WLA[362]
+WLA[361] WLA[360] WLA[359] WLA[358] WLA[357] WLA[356] WLA[355] WLA[354] WLA[353] WLA[352]
+WLA[351] WLA[350] WLA[349] WLA[348] WLA[347] WLA[346] WLA[345] WLA[344] WLA[343] WLA[342]
+WLA[341] WLA[340] WLA[339] WLA[338] WLA[337] WLA[336] WLA[335] WLA[334] WLA[333] WLA[332]
+WLA[331] WLA[330] WLA[329] WLA[328] WLA[327] WLA[326] WLA[325] WLA[324] WLA[323] WLA[322]
+WLA[321] WLA[320] WLA[319] WLA[318] WLA[317] WLA[316] WLA[315] WLA[314] WLA[313] WLA[312]
+WLA[311] WLA[310] WLA[309] WLA[308] WLA[307] WLA[306] WLA[305] WLA[304] WLA[303] WLA[302]
+WLA[301] WLA[300] WLA[299] WLA[298] WLA[297] WLA[296] WLA[295] WLA[294] WLA[293] WLA[292]
+WLA[291] WLA[290] WLA[289] WLA[288] WLA[287] WLA[286] WLA[285] WLA[284] WLA[283] WLA[282]
+WLA[281] WLA[280] WLA[279] WLA[278] WLA[277] WLA[276] WLA[275] WLA[274] WLA[273] WLA[272]
+WLA[271] WLA[270] WLA[269] WLA[268] WLA[267] WLA[266] WLA[265] WLA[264] WLA[263] WLA[262]
+WLA[261] WLA[260] WLA[259] WLA[258] WLA[257] WLA[256] WLA[255] WLA[254] WLA[253] WLA[252]
+WLA[251] WLA[250] WLA[249] WLA[248] WLA[247] WLA[246] WLA[245] WLA[244] WLA[243] WLA[242]
+WLA[241] WLA[240] WLA[239] WLA[238] WLA[237] WLA[236] WLA[235] WLA[234] WLA[233] WLA[232]
+WLA[231] WLA[230] WLA[229] WLA[228] WLA[227] WLA[226] WLA[225] WLA[224] WLA[223] WLA[222]
+WLA[221] WLA[220] WLA[219] WLA[218] WLA[217] WLA[216] WLA[215] WLA[214] WLA[213] WLA[212]
+WLA[211] WLA[210] WLA[209] WLA[208] WLA[207] WLA[206] WLA[205] WLA[204] WLA[203] WLA[202]
+WLA[201] WLA[200] WLA[199] WLA[198] WLA[197] WLA[196] WLA[195] WLA[194] WLA[193] WLA[192]
+WLA[191] WLA[190] WLA[189] WLA[188] WLA[187] WLA[186] WLA[185] WLA[184] WLA[183] WLA[182]
+WLA[181] WLA[180] WLA[179] WLA[178] WLA[177] WLA[176] WLA[175] WLA[174] WLA[173] WLA[172]
+WLA[171] WLA[170] WLA[169] WLA[168] WLA[167] WLA[166] WLA[165] WLA[164] WLA[163] WLA[162]
+WLA[161] WLA[160] WLA[159] WLA[158] WLA[157] WLA[156] WLA[155] WLA[154] WLA[153] WLA[152]
+WLA[151] WLA[150] WLA[149] WLA[148] WLA[147] WLA[146] WLA[145] WLA[144] WLA[143] WLA[142]
+WLA[141] WLA[140] WLA[139] WLA[138] WLA[137] WLA[136] WLA[135] WLA[134] WLA[133] WLA[132]
+WLA[131] WLA[130] WLA[129] WLA[128] WLA[127] WLA[126] WLA[125] WLA[124] WLA[123] WLA[122]
+WLA[121] WLA[120] WLA[119] WLA[118] WLA[117] WLA[116] WLA[115] WLA[114] WLA[113] WLA[112]
+WLA[111] WLA[110] WLA[109] WLA[108] WLA[107] WLA[106] WLA[105] WLA[104] WLA[103] WLA[102]
+WLA[101] WLA[100] WLA[99] WLA[98] WLA[97] WLA[96] WLA[95] WLA[94] WLA[93] WLA[92]
+WLA[91] WLA[90] WLA[89] WLA[88] WLA[87] WLA[86] WLA[85] WLA[84] WLA[83] WLA[82]
+WLA[81] WLA[80] WLA[79] WLA[78] WLA[77] WLA[76] WLA[75] WLA[74] WLA[73] WLA[72]
+WLA[71] WLA[70] WLA[69] WLA[68] WLA[67] WLA[66] WLA[65] WLA[64] WLA[63] WLA[62]
+WLA[61] WLA[60] WLA[59] WLA[58] WLA[57] WLA[56] WLA[55] WLA[54] WLA[53] WLA[52]
+WLA[51] WLA[50] WLA[49] WLA[48] WLA[47] WLA[46] WLA[45] WLA[44] WLA[43] WLA[42]
+WLA[41] WLA[40] WLA[39] WLA[38] WLA[37] WLA[36] WLA[35] WLA[34] WLA[33] WLA[32]
+WLA[31] WLA[30] WLA[29] WLA[28] WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22]
+WLA[21] WLA[20] WLA[19] WLA[18] WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12]
+WLA[11] WLA[10] WLA[9] WLA[8] WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2]
+WLA[1] WLA[0] WLB[511] WLB[510] WLB[509] WLB[508] WLB[507] WLB[506] WLB[505] WLB[504]
+WLB[503] WLB[502] WLB[501] WLB[500] WLB[499] WLB[498] WLB[497] WLB[496] WLB[495] WLB[494]
+WLB[493] WLB[492] WLB[491] WLB[490] WLB[489] WLB[488] WLB[487] WLB[486] WLB[485] WLB[484]
+WLB[483] WLB[482] WLB[481] WLB[480] WLB[479] WLB[478] WLB[477] WLB[476] WLB[475] WLB[474]
+WLB[473] WLB[472] WLB[471] WLB[470] WLB[469] WLB[468] WLB[467] WLB[466] WLB[465] WLB[464]
+WLB[463] WLB[462] WLB[461] WLB[460] WLB[459] WLB[458] WLB[457] WLB[456] WLB[455] WLB[454]
+WLB[453] WLB[452] WLB[451] WLB[450] WLB[449] WLB[448] WLB[447] WLB[446] WLB[445] WLB[444]
+WLB[443] WLB[442] WLB[441] WLB[440] WLB[439] WLB[438] WLB[437] WLB[436] WLB[435] WLB[434]
+WLB[433] WLB[432] WLB[431] WLB[430] WLB[429] WLB[428] WLB[427] WLB[426] WLB[425] WLB[424]
+WLB[423] WLB[422] WLB[421] WLB[420] WLB[419] WLB[418] WLB[417] WLB[416] WLB[415] WLB[414]
+WLB[413] WLB[412] WLB[411] WLB[410] WLB[409] WLB[408] WLB[407] WLB[406] WLB[405] WLB[404]
+WLB[403] WLB[402] WLB[401] WLB[400] WLB[399] WLB[398] WLB[397] WLB[396] WLB[395] WLB[394]
+WLB[393] WLB[392] WLB[391] WLB[390] WLB[389] WLB[388] WLB[387] WLB[386] WLB[385] WLB[384]
+WLB[383] WLB[382] WLB[381] WLB[380] WLB[379] WLB[378] WLB[377] WLB[376] WLB[375] WLB[374]
+WLB[373] WLB[372] WLB[371] WLB[370] WLB[369] WLB[368] WLB[367] WLB[366] WLB[365] WLB[364]
+WLB[363] WLB[362] WLB[361] WLB[360] WLB[359] WLB[358] WLB[357] WLB[356] WLB[355] WLB[354]
+WLB[353] WLB[352] WLB[351] WLB[350] WLB[349] WLB[348] WLB[347] WLB[346] WLB[345] WLB[344]
+WLB[343] WLB[342] WLB[341] WLB[340] WLB[339] WLB[338] WLB[337] WLB[336] WLB[335] WLB[334]
+WLB[333] WLB[332] WLB[331] WLB[330] WLB[329] WLB[328] WLB[327] WLB[326] WLB[325] WLB[324]
+WLB[323] WLB[322] WLB[321] WLB[320] WLB[319] WLB[318] WLB[317] WLB[316] WLB[315] WLB[314]
+WLB[313] WLB[312] WLB[311] WLB[310] WLB[309] WLB[308] WLB[307] WLB[306] WLB[305] WLB[304]
+WLB[303] WLB[302] WLB[301] WLB[300] WLB[299] WLB[298] WLB[297] WLB[296] WLB[295] WLB[294]
+WLB[293] WLB[292] WLB[291] WLB[290] WLB[289] WLB[288] WLB[287] WLB[286] WLB[285] WLB[284]
+WLB[283] WLB[282] WLB[281] WLB[280] WLB[279] WLB[278] WLB[277] WLB[276] WLB[275] WLB[274]
+WLB[273] WLB[272] WLB[271] WLB[270] WLB[269] WLB[268] WLB[267] WLB[266] WLB[265] WLB[264]
+WLB[263] WLB[262] WLB[261] WLB[260] WLB[259] WLB[258] WLB[257] WLB[256] WLB[255] WLB[254]
+WLB[253] WLB[252] WLB[251] WLB[250] WLB[249] WLB[248] WLB[247] WLB[246] WLB[245] WLB[244]
+WLB[243] WLB[242] WLB[241] WLB[240] WLB[239] WLB[238] WLB[237] WLB[236] WLB[235] WLB[234]
+WLB[233] WLB[232] WLB[231] WLB[230] WLB[229] WLB[228] WLB[227] WLB[226] WLB[225] WLB[224]
+WLB[223] WLB[222] WLB[221] WLB[220] WLB[219] WLB[218] WLB[217] WLB[216] WLB[215] WLB[214]
+WLB[213] WLB[212] WLB[211] WLB[210] WLB[209] WLB[208] WLB[207] WLB[206] WLB[205] WLB[204]
+WLB[203] WLB[202] WLB[201] WLB[200] WLB[199] WLB[198] WLB[197] WLB[196] WLB[195] WLB[194]
+WLB[193] WLB[192] WLB[191] WLB[190] WLB[189] WLB[188] WLB[187] WLB[186] WLB[185] WLB[184]
+WLB[183] WLB[182] WLB[181] WLB[180] WLB[179] WLB[178] WLB[177] WLB[176] WLB[175] WLB[174]
+WLB[173] WLB[172] WLB[171] WLB[170] WLB[169] WLB[168] WLB[167] WLB[166] WLB[165] WLB[164]
+WLB[163] WLB[162] WLB[161] WLB[160] WLB[159] WLB[158] WLB[157] WLB[156] WLB[155] WLB[154]
+WLB[153] WLB[152] WLB[151] WLB[150] WLB[149] WLB[148] WLB[147] WLB[146] WLB[145] WLB[144]
+WLB[143] WLB[142] WLB[141] WLB[140] WLB[139] WLB[138] WLB[137] WLB[136] WLB[135] WLB[134]
+WLB[133] WLB[132] WLB[131] WLB[130] WLB[129] WLB[128] WLB[127] WLB[126] WLB[125] WLB[124]
+WLB[123] WLB[122] WLB[121] WLB[120] WLB[119] WLB[118] WLB[117] WLB[116] WLB[115] WLB[114]
+WLB[113] WLB[112] WLB[111] WLB[110] WLB[109] WLB[108] WLB[107] WLB[106] WLB[105] WLB[104]
+WLB[103] WLB[102] WLB[101] WLB[100] WLB[99] WLB[98] WLB[97] WLB[96] WLB[95] WLB[94]
+WLB[93] WLB[92] WLB[91] WLB[90] WLB[89] WLB[88] WLB[87] WLB[86] WLB[85] WLB[84]
+WLB[83] WLB[82] WLB[81] WLB[80] WLB[79] WLB[78] WLB[77] WLB[76] WLB[75] WLB[74]
+WLB[73] WLB[72] WLB[71] WLB[70] WLB[69] WLB[68] WLB[67] WLB[66] WLB[65] WLB[64]
+WLB[63] WLB[62] WLB[61] WLB[60] WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54]
+WLB[53] WLB[52] WLB[51] WLB[50] WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44]
+WLB[43] WLB[42] WLB[41] WLB[40] WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34]
+WLB[33] WLB[32] WLB[31] WLB[30] WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24]
+WLB[23] WLB[22] WLB[21] WLB[20] WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14]
+WLB[13] WLB[12] WLB[11] WLB[10] WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4]
+WLB[3] WLB[2] WLB[1] WLB[0] YXA[7] YXA[6] YXA[5] YXA[4] YXA[3] YXA[2]
+YXA[1] YXA[0] YXB[7] YXB[6] YXB[5] YXB[4] YXB[3] YXB[2] YXB[1] YXB[0] S55NLLGDPH_X512Y8D16_BW_Y512X8CELL_BW
XI19 BWENA[3] BWENB[3] CLKA CLKB CLKXA CLKXB DATAA[3] DATAB[3] DOUTA[3] DOUTB[3]
+VSS STWLA STWLA VSS VSS VSS VSS VSS STWLB VSS
+VSS VSS STWLB VSS VSS VSS RWLA[0] RWLA[1] RWLB[0] RWLB[1]
+SACK1A SACK1B SACK4A SACK4B VDD VSS WEA WEB WLA[511] WLA[510]
+WLA[509] WLA[508] WLA[507] WLA[506] WLA[505] WLA[504] WLA[503] WLA[502] WLA[501] WLA[500]
+WLA[499] WLA[498] WLA[497] WLA[496] WLA[495] WLA[494] WLA[493] WLA[492] WLA[491] WLA[490]
+WLA[489] WLA[488] WLA[487] WLA[486] WLA[485] WLA[484] WLA[483] WLA[482] WLA[481] WLA[480]
+WLA[479] WLA[478] WLA[477] WLA[476] WLA[475] WLA[474] WLA[473] WLA[472] WLA[471] WLA[470]
+WLA[469] WLA[468] WLA[467] WLA[466] WLA[465] WLA[464] WLA[463] WLA[462] WLA[461] WLA[460]
+WLA[459] WLA[458] WLA[457] WLA[456] WLA[455] WLA[454] WLA[453] WLA[452] WLA[451] WLA[450]
+WLA[449] WLA[448] WLA[447] WLA[446] WLA[445] WLA[444] WLA[443] WLA[442] WLA[441] WLA[440]
+WLA[439] WLA[438] WLA[437] WLA[436] WLA[435] WLA[434] WLA[433] WLA[432] WLA[431] WLA[430]
+WLA[429] WLA[428] WLA[427] WLA[426] WLA[425] WLA[424] WLA[423] WLA[422] WLA[421] WLA[420]
+WLA[419] WLA[418] WLA[417] WLA[416] WLA[415] WLA[414] WLA[413] WLA[412] WLA[411] WLA[410]
+WLA[409] WLA[408] WLA[407] WLA[406] WLA[405] WLA[404] WLA[403] WLA[402] WLA[401] WLA[400]
+WLA[399] WLA[398] WLA[397] WLA[396] WLA[395] WLA[394] WLA[393] WLA[392] WLA[391] WLA[390]
+WLA[389] WLA[388] WLA[387] WLA[386] WLA[385] WLA[384] WLA[383] WLA[382] WLA[381] WLA[380]
+WLA[379] WLA[378] WLA[377] WLA[376] WLA[375] WLA[374] WLA[373] WLA[372] WLA[371] WLA[370]
+WLA[369] WLA[368] WLA[367] WLA[366] WLA[365] WLA[364] WLA[363] WLA[362] WLA[361] WLA[360]
+WLA[359] WLA[358] WLA[357] WLA[356] WLA[355] WLA[354] WLA[353] WLA[352] WLA[351] WLA[350]
+WLA[349] WLA[348] WLA[347] WLA[346] WLA[345] WLA[344] WLA[343] WLA[342] WLA[341] WLA[340]
+WLA[339] WLA[338] WLA[337] WLA[336] WLA[335] WLA[334] WLA[333] WLA[332] WLA[331] WLA[330]
+WLA[329] WLA[328] WLA[327] WLA[326] WLA[325] WLA[324] WLA[323] WLA[322] WLA[321] WLA[320]
+WLA[319] WLA[318] WLA[317] WLA[316] WLA[315] WLA[314] WLA[313] WLA[312] WLA[311] WLA[310]
+WLA[309] WLA[308] WLA[307] WLA[306] WLA[305] WLA[304] WLA[303] WLA[302] WLA[301] WLA[300]
+WLA[299] WLA[298] WLA[297] WLA[296] WLA[295] WLA[294] WLA[293] WLA[292] WLA[291] WLA[290]
+WLA[289] WLA[288] WLA[287] WLA[286] WLA[285] WLA[284] WLA[283] WLA[282] WLA[281] WLA[280]
+WLA[279] WLA[278] WLA[277] WLA[276] WLA[275] WLA[274] WLA[273] WLA[272] WLA[271] WLA[270]
+WLA[269] WLA[268] WLA[267] WLA[266] WLA[265] WLA[264] WLA[263] WLA[262] WLA[261] WLA[260]
+WLA[259] WLA[258] WLA[257] WLA[256] WLA[255] WLA[254] WLA[253] WLA[252] WLA[251] WLA[250]
+WLA[249] WLA[248] WLA[247] WLA[246] WLA[245] WLA[244] WLA[243] WLA[242] WLA[241] WLA[240]
+WLA[239] WLA[238] WLA[237] WLA[236] WLA[235] WLA[234] WLA[233] WLA[232] WLA[231] WLA[230]
+WLA[229] WLA[228] WLA[227] WLA[226] WLA[225] WLA[224] WLA[223] WLA[222] WLA[221] WLA[220]
+WLA[219] WLA[218] WLA[217] WLA[216] WLA[215] WLA[214] WLA[213] WLA[212] WLA[211] WLA[210]
+WLA[209] WLA[208] WLA[207] WLA[206] WLA[205] WLA[204] WLA[203] WLA[202] WLA[201] WLA[200]
+WLA[199] WLA[198] WLA[197] WLA[196] WLA[195] WLA[194] WLA[193] WLA[192] WLA[191] WLA[190]
+WLA[189] WLA[188] WLA[187] WLA[186] WLA[185] WLA[184] WLA[183] WLA[182] WLA[181] WLA[180]
+WLA[179] WLA[178] WLA[177] WLA[176] WLA[175] WLA[174] WLA[173] WLA[172] WLA[171] WLA[170]
+WLA[169] WLA[168] WLA[167] WLA[166] WLA[165] WLA[164] WLA[163] WLA[162] WLA[161] WLA[160]
+WLA[159] WLA[158] WLA[157] WLA[156] WLA[155] WLA[154] WLA[153] WLA[152] WLA[151] WLA[150]
+WLA[149] WLA[148] WLA[147] WLA[146] WLA[145] WLA[144] WLA[143] WLA[142] WLA[141] WLA[140]
+WLA[139] WLA[138] WLA[137] WLA[136] WLA[135] WLA[134] WLA[133] WLA[132] WLA[131] WLA[130]
+WLA[129] WLA[128] WLA[127] WLA[126] WLA[125] WLA[124] WLA[123] WLA[122] WLA[121] WLA[120]
+WLA[119] WLA[118] WLA[117] WLA[116] WLA[115] WLA[114] WLA[113] WLA[112] WLA[111] WLA[110]
+WLA[109] WLA[108] WLA[107] WLA[106] WLA[105] WLA[104] WLA[103] WLA[102] WLA[101] WLA[100]
+WLA[99] WLA[98] WLA[97] WLA[96] WLA[95] WLA[94] WLA[93] WLA[92] WLA[91] WLA[90]
+WLA[89] WLA[88] WLA[87] WLA[86] WLA[85] WLA[84] WLA[83] WLA[82] WLA[81] WLA[80]
+WLA[79] WLA[78] WLA[77] WLA[76] WLA[75] WLA[74] WLA[73] WLA[72] WLA[71] WLA[70]
+WLA[69] WLA[68] WLA[67] WLA[66] WLA[65] WLA[64] WLA[63] WLA[62] WLA[61] WLA[60]
+WLA[59] WLA[58] WLA[57] WLA[56] WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50]
+WLA[49] WLA[48] WLA[47] WLA[46] WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40]
+WLA[39] WLA[38] WLA[37] WLA[36] WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30]
+WLA[29] WLA[28] WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20]
+WLA[19] WLA[18] WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10]
+WLA[9] WLA[8] WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0]
+WLB[511] WLB[510] WLB[509] WLB[508] WLB[507] WLB[506] WLB[505] WLB[504] WLB[503] WLB[502]
+WLB[501] WLB[500] WLB[499] WLB[498] WLB[497] WLB[496] WLB[495] WLB[494] WLB[493] WLB[492]
+WLB[491] WLB[490] WLB[489] WLB[488] WLB[487] WLB[486] WLB[485] WLB[484] WLB[483] WLB[482]
+WLB[481] WLB[480] WLB[479] WLB[478] WLB[477] WLB[476] WLB[475] WLB[474] WLB[473] WLB[472]
+WLB[471] WLB[470] WLB[469] WLB[468] WLB[467] WLB[466] WLB[465] WLB[464] WLB[463] WLB[462]
+WLB[461] WLB[460] WLB[459] WLB[458] WLB[457] WLB[456] WLB[455] WLB[454] WLB[453] WLB[452]
+WLB[451] WLB[450] WLB[449] WLB[448] WLB[447] WLB[446] WLB[445] WLB[444] WLB[443] WLB[442]
+WLB[441] WLB[440] WLB[439] WLB[438] WLB[437] WLB[436] WLB[435] WLB[434] WLB[433] WLB[432]
+WLB[431] WLB[430] WLB[429] WLB[428] WLB[427] WLB[426] WLB[425] WLB[424] WLB[423] WLB[422]
+WLB[421] WLB[420] WLB[419] WLB[418] WLB[417] WLB[416] WLB[415] WLB[414] WLB[413] WLB[412]
+WLB[411] WLB[410] WLB[409] WLB[408] WLB[407] WLB[406] WLB[405] WLB[404] WLB[403] WLB[402]
+WLB[401] WLB[400] WLB[399] WLB[398] WLB[397] WLB[396] WLB[395] WLB[394] WLB[393] WLB[392]
+WLB[391] WLB[390] WLB[389] WLB[388] WLB[387] WLB[386] WLB[385] WLB[384] WLB[383] WLB[382]
+WLB[381] WLB[380] WLB[379] WLB[378] WLB[377] WLB[376] WLB[375] WLB[374] WLB[373] WLB[372]
+WLB[371] WLB[370] WLB[369] WLB[368] WLB[367] WLB[366] WLB[365] WLB[364] WLB[363] WLB[362]
+WLB[361] WLB[360] WLB[359] WLB[358] WLB[357] WLB[356] WLB[355] WLB[354] WLB[353] WLB[352]
+WLB[351] WLB[350] WLB[349] WLB[348] WLB[347] WLB[346] WLB[345] WLB[344] WLB[343] WLB[342]
+WLB[341] WLB[340] WLB[339] WLB[338] WLB[337] WLB[336] WLB[335] WLB[334] WLB[333] WLB[332]
+WLB[331] WLB[330] WLB[329] WLB[328] WLB[327] WLB[326] WLB[325] WLB[324] WLB[323] WLB[322]
+WLB[321] WLB[320] WLB[319] WLB[318] WLB[317] WLB[316] WLB[315] WLB[314] WLB[313] WLB[312]
+WLB[311] WLB[310] WLB[309] WLB[308] WLB[307] WLB[306] WLB[305] WLB[304] WLB[303] WLB[302]
+WLB[301] WLB[300] WLB[299] WLB[298] WLB[297] WLB[296] WLB[295] WLB[294] WLB[293] WLB[292]
+WLB[291] WLB[290] WLB[289] WLB[288] WLB[287] WLB[286] WLB[285] WLB[284] WLB[283] WLB[282]
+WLB[281] WLB[280] WLB[279] WLB[278] WLB[277] WLB[276] WLB[275] WLB[274] WLB[273] WLB[272]
+WLB[271] WLB[270] WLB[269] WLB[268] WLB[267] WLB[266] WLB[265] WLB[264] WLB[263] WLB[262]
+WLB[261] WLB[260] WLB[259] WLB[258] WLB[257] WLB[256] WLB[255] WLB[254] WLB[253] WLB[252]
+WLB[251] WLB[250] WLB[249] WLB[248] WLB[247] WLB[246] WLB[245] WLB[244] WLB[243] WLB[242]
+WLB[241] WLB[240] WLB[239] WLB[238] WLB[237] WLB[236] WLB[235] WLB[234] WLB[233] WLB[232]
+WLB[231] WLB[230] WLB[229] WLB[228] WLB[227] WLB[226] WLB[225] WLB[224] WLB[223] WLB[222]
+WLB[221] WLB[220] WLB[219] WLB[218] WLB[217] WLB[216] WLB[215] WLB[214] WLB[213] WLB[212]
+WLB[211] WLB[210] WLB[209] WLB[208] WLB[207] WLB[206] WLB[205] WLB[204] WLB[203] WLB[202]
+WLB[201] WLB[200] WLB[199] WLB[198] WLB[197] WLB[196] WLB[195] WLB[194] WLB[193] WLB[192]
+WLB[191] WLB[190] WLB[189] WLB[188] WLB[187] WLB[186] WLB[185] WLB[184] WLB[183] WLB[182]
+WLB[181] WLB[180] WLB[179] WLB[178] WLB[177] WLB[176] WLB[175] WLB[174] WLB[173] WLB[172]
+WLB[171] WLB[170] WLB[169] WLB[168] WLB[167] WLB[166] WLB[165] WLB[164] WLB[163] WLB[162]
+WLB[161] WLB[160] WLB[159] WLB[158] WLB[157] WLB[156] WLB[155] WLB[154] WLB[153] WLB[152]
+WLB[151] WLB[150] WLB[149] WLB[148] WLB[147] WLB[146] WLB[145] WLB[144] WLB[143] WLB[142]
+WLB[141] WLB[140] WLB[139] WLB[138] WLB[137] WLB[136] WLB[135] WLB[134] WLB[133] WLB[132]
+WLB[131] WLB[130] WLB[129] WLB[128] WLB[127] WLB[126] WLB[125] WLB[124] WLB[123] WLB[122]
+WLB[121] WLB[120] WLB[119] WLB[118] WLB[117] WLB[116] WLB[115] WLB[114] WLB[113] WLB[112]
+WLB[111] WLB[110] WLB[109] WLB[108] WLB[107] WLB[106] WLB[105] WLB[104] WLB[103] WLB[102]
+WLB[101] WLB[100] WLB[99] WLB[98] WLB[97] WLB[96] WLB[95] WLB[94] WLB[93] WLB[92]
+WLB[91] WLB[90] WLB[89] WLB[88] WLB[87] WLB[86] WLB[85] WLB[84] WLB[83] WLB[82]
+WLB[81] WLB[80] WLB[79] WLB[78] WLB[77] WLB[76] WLB[75] WLB[74] WLB[73] WLB[72]
+WLB[71] WLB[70] WLB[69] WLB[68] WLB[67] WLB[66] WLB[65] WLB[64] WLB[63] WLB[62]
+WLB[61] WLB[60] WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54] WLB[53] WLB[52]
+WLB[51] WLB[50] WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44] WLB[43] WLB[42]
+WLB[41] WLB[40] WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34] WLB[33] WLB[32]
+WLB[31] WLB[30] WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24] WLB[23] WLB[22]
+WLB[21] WLB[20] WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14] WLB[13] WLB[12]
+WLB[11] WLB[10] WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4] WLB[3] WLB[2]
+WLB[1] WLB[0] YXA[7] YXA[6] YXA[5] YXA[4] YXA[3] YXA[2] YXA[1] YXA[0]
+YXB[7] YXB[6] YXB[5] YXB[4] YXB[3] YXB[2] YXB[1] YXB[0] S55NLLGDPH_X512Y8D16_BW_Y512X8CELL_MID
XI20 BWENA[4] BWENB[4] CLKA CLKB CLKXA CLKXB DATAA[4] DATAB[4] DOUTA[4] DOUTB[4]
+VSS VSS VSS VSS STWLB VSS VSS VSS RWLA[0] RWLA[1]
+RWLB[0] RWLB[1] SACK1A SACK1B SACK4A SACK4B VDD VSS WEA WEB
+WLA[511] WLA[510] WLA[509] WLA[508] WLA[507] WLA[506] WLA[505] WLA[504] WLA[503] WLA[502]
+WLA[501] WLA[500] WLA[499] WLA[498] WLA[497] WLA[496] WLA[495] WLA[494] WLA[493] WLA[492]
+WLA[491] WLA[490] WLA[489] WLA[488] WLA[487] WLA[486] WLA[485] WLA[484] WLA[483] WLA[482]
+WLA[481] WLA[480] WLA[479] WLA[478] WLA[477] WLA[476] WLA[475] WLA[474] WLA[473] WLA[472]
+WLA[471] WLA[470] WLA[469] WLA[468] WLA[467] WLA[466] WLA[465] WLA[464] WLA[463] WLA[462]
+WLA[461] WLA[460] WLA[459] WLA[458] WLA[457] WLA[456] WLA[455] WLA[454] WLA[453] WLA[452]
+WLA[451] WLA[450] WLA[449] WLA[448] WLA[447] WLA[446] WLA[445] WLA[444] WLA[443] WLA[442]
+WLA[441] WLA[440] WLA[439] WLA[438] WLA[437] WLA[436] WLA[435] WLA[434] WLA[433] WLA[432]
+WLA[431] WLA[430] WLA[429] WLA[428] WLA[427] WLA[426] WLA[425] WLA[424] WLA[423] WLA[422]
+WLA[421] WLA[420] WLA[419] WLA[418] WLA[417] WLA[416] WLA[415] WLA[414] WLA[413] WLA[412]
+WLA[411] WLA[410] WLA[409] WLA[408] WLA[407] WLA[406] WLA[405] WLA[404] WLA[403] WLA[402]
+WLA[401] WLA[400] WLA[399] WLA[398] WLA[397] WLA[396] WLA[395] WLA[394] WLA[393] WLA[392]
+WLA[391] WLA[390] WLA[389] WLA[388] WLA[387] WLA[386] WLA[385] WLA[384] WLA[383] WLA[382]
+WLA[381] WLA[380] WLA[379] WLA[378] WLA[377] WLA[376] WLA[375] WLA[374] WLA[373] WLA[372]
+WLA[371] WLA[370] WLA[369] WLA[368] WLA[367] WLA[366] WLA[365] WLA[364] WLA[363] WLA[362]
+WLA[361] WLA[360] WLA[359] WLA[358] WLA[357] WLA[356] WLA[355] WLA[354] WLA[353] WLA[352]
+WLA[351] WLA[350] WLA[349] WLA[348] WLA[347] WLA[346] WLA[345] WLA[344] WLA[343] WLA[342]
+WLA[341] WLA[340] WLA[339] WLA[338] WLA[337] WLA[336] WLA[335] WLA[334] WLA[333] WLA[332]
+WLA[331] WLA[330] WLA[329] WLA[328] WLA[327] WLA[326] WLA[325] WLA[324] WLA[323] WLA[322]
+WLA[321] WLA[320] WLA[319] WLA[318] WLA[317] WLA[316] WLA[315] WLA[314] WLA[313] WLA[312]
+WLA[311] WLA[310] WLA[309] WLA[308] WLA[307] WLA[306] WLA[305] WLA[304] WLA[303] WLA[302]
+WLA[301] WLA[300] WLA[299] WLA[298] WLA[297] WLA[296] WLA[295] WLA[294] WLA[293] WLA[292]
+WLA[291] WLA[290] WLA[289] WLA[288] WLA[287] WLA[286] WLA[285] WLA[284] WLA[283] WLA[282]
+WLA[281] WLA[280] WLA[279] WLA[278] WLA[277] WLA[276] WLA[275] WLA[274] WLA[273] WLA[272]
+WLA[271] WLA[270] WLA[269] WLA[268] WLA[267] WLA[266] WLA[265] WLA[264] WLA[263] WLA[262]
+WLA[261] WLA[260] WLA[259] WLA[258] WLA[257] WLA[256] WLA[255] WLA[254] WLA[253] WLA[252]
+WLA[251] WLA[250] WLA[249] WLA[248] WLA[247] WLA[246] WLA[245] WLA[244] WLA[243] WLA[242]
+WLA[241] WLA[240] WLA[239] WLA[238] WLA[237] WLA[236] WLA[235] WLA[234] WLA[233] WLA[232]
+WLA[231] WLA[230] WLA[229] WLA[228] WLA[227] WLA[226] WLA[225] WLA[224] WLA[223] WLA[222]
+WLA[221] WLA[220] WLA[219] WLA[218] WLA[217] WLA[216] WLA[215] WLA[214] WLA[213] WLA[212]
+WLA[211] WLA[210] WLA[209] WLA[208] WLA[207] WLA[206] WLA[205] WLA[204] WLA[203] WLA[202]
+WLA[201] WLA[200] WLA[199] WLA[198] WLA[197] WLA[196] WLA[195] WLA[194] WLA[193] WLA[192]
+WLA[191] WLA[190] WLA[189] WLA[188] WLA[187] WLA[186] WLA[185] WLA[184] WLA[183] WLA[182]
+WLA[181] WLA[180] WLA[179] WLA[178] WLA[177] WLA[176] WLA[175] WLA[174] WLA[173] WLA[172]
+WLA[171] WLA[170] WLA[169] WLA[168] WLA[167] WLA[166] WLA[165] WLA[164] WLA[163] WLA[162]
+WLA[161] WLA[160] WLA[159] WLA[158] WLA[157] WLA[156] WLA[155] WLA[154] WLA[153] WLA[152]
+WLA[151] WLA[150] WLA[149] WLA[148] WLA[147] WLA[146] WLA[145] WLA[144] WLA[143] WLA[142]
+WLA[141] WLA[140] WLA[139] WLA[138] WLA[137] WLA[136] WLA[135] WLA[134] WLA[133] WLA[132]
+WLA[131] WLA[130] WLA[129] WLA[128] WLA[127] WLA[126] WLA[125] WLA[124] WLA[123] WLA[122]
+WLA[121] WLA[120] WLA[119] WLA[118] WLA[117] WLA[116] WLA[115] WLA[114] WLA[113] WLA[112]
+WLA[111] WLA[110] WLA[109] WLA[108] WLA[107] WLA[106] WLA[105] WLA[104] WLA[103] WLA[102]
+WLA[101] WLA[100] WLA[99] WLA[98] WLA[97] WLA[96] WLA[95] WLA[94] WLA[93] WLA[92]
+WLA[91] WLA[90] WLA[89] WLA[88] WLA[87] WLA[86] WLA[85] WLA[84] WLA[83] WLA[82]
+WLA[81] WLA[80] WLA[79] WLA[78] WLA[77] WLA[76] WLA[75] WLA[74] WLA[73] WLA[72]
+WLA[71] WLA[70] WLA[69] WLA[68] WLA[67] WLA[66] WLA[65] WLA[64] WLA[63] WLA[62]
+WLA[61] WLA[60] WLA[59] WLA[58] WLA[57] WLA[56] WLA[55] WLA[54] WLA[53] WLA[52]
+WLA[51] WLA[50] WLA[49] WLA[48] WLA[47] WLA[46] WLA[45] WLA[44] WLA[43] WLA[42]
+WLA[41] WLA[40] WLA[39] WLA[38] WLA[37] WLA[36] WLA[35] WLA[34] WLA[33] WLA[32]
+WLA[31] WLA[30] WLA[29] WLA[28] WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22]
+WLA[21] WLA[20] WLA[19] WLA[18] WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12]
+WLA[11] WLA[10] WLA[9] WLA[8] WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2]
+WLA[1] WLA[0] WLB[511] WLB[510] WLB[509] WLB[508] WLB[507] WLB[506] WLB[505] WLB[504]
+WLB[503] WLB[502] WLB[501] WLB[500] WLB[499] WLB[498] WLB[497] WLB[496] WLB[495] WLB[494]
+WLB[493] WLB[492] WLB[491] WLB[490] WLB[489] WLB[488] WLB[487] WLB[486] WLB[485] WLB[484]
+WLB[483] WLB[482] WLB[481] WLB[480] WLB[479] WLB[478] WLB[477] WLB[476] WLB[475] WLB[474]
+WLB[473] WLB[472] WLB[471] WLB[470] WLB[469] WLB[468] WLB[467] WLB[466] WLB[465] WLB[464]
+WLB[463] WLB[462] WLB[461] WLB[460] WLB[459] WLB[458] WLB[457] WLB[456] WLB[455] WLB[454]
+WLB[453] WLB[452] WLB[451] WLB[450] WLB[449] WLB[448] WLB[447] WLB[446] WLB[445] WLB[444]
+WLB[443] WLB[442] WLB[441] WLB[440] WLB[439] WLB[438] WLB[437] WLB[436] WLB[435] WLB[434]
+WLB[433] WLB[432] WLB[431] WLB[430] WLB[429] WLB[428] WLB[427] WLB[426] WLB[425] WLB[424]
+WLB[423] WLB[422] WLB[421] WLB[420] WLB[419] WLB[418] WLB[417] WLB[416] WLB[415] WLB[414]
+WLB[413] WLB[412] WLB[411] WLB[410] WLB[409] WLB[408] WLB[407] WLB[406] WLB[405] WLB[404]
+WLB[403] WLB[402] WLB[401] WLB[400] WLB[399] WLB[398] WLB[397] WLB[396] WLB[395] WLB[394]
+WLB[393] WLB[392] WLB[391] WLB[390] WLB[389] WLB[388] WLB[387] WLB[386] WLB[385] WLB[384]
+WLB[383] WLB[382] WLB[381] WLB[380] WLB[379] WLB[378] WLB[377] WLB[376] WLB[375] WLB[374]
+WLB[373] WLB[372] WLB[371] WLB[370] WLB[369] WLB[368] WLB[367] WLB[366] WLB[365] WLB[364]
+WLB[363] WLB[362] WLB[361] WLB[360] WLB[359] WLB[358] WLB[357] WLB[356] WLB[355] WLB[354]
+WLB[353] WLB[352] WLB[351] WLB[350] WLB[349] WLB[348] WLB[347] WLB[346] WLB[345] WLB[344]
+WLB[343] WLB[342] WLB[341] WLB[340] WLB[339] WLB[338] WLB[337] WLB[336] WLB[335] WLB[334]
+WLB[333] WLB[332] WLB[331] WLB[330] WLB[329] WLB[328] WLB[327] WLB[326] WLB[325] WLB[324]
+WLB[323] WLB[322] WLB[321] WLB[320] WLB[319] WLB[318] WLB[317] WLB[316] WLB[315] WLB[314]
+WLB[313] WLB[312] WLB[311] WLB[310] WLB[309] WLB[308] WLB[307] WLB[306] WLB[305] WLB[304]
+WLB[303] WLB[302] WLB[301] WLB[300] WLB[299] WLB[298] WLB[297] WLB[296] WLB[295] WLB[294]
+WLB[293] WLB[292] WLB[291] WLB[290] WLB[289] WLB[288] WLB[287] WLB[286] WLB[285] WLB[284]
+WLB[283] WLB[282] WLB[281] WLB[280] WLB[279] WLB[278] WLB[277] WLB[276] WLB[275] WLB[274]
+WLB[273] WLB[272] WLB[271] WLB[270] WLB[269] WLB[268] WLB[267] WLB[266] WLB[265] WLB[264]
+WLB[263] WLB[262] WLB[261] WLB[260] WLB[259] WLB[258] WLB[257] WLB[256] WLB[255] WLB[254]
+WLB[253] WLB[252] WLB[251] WLB[250] WLB[249] WLB[248] WLB[247] WLB[246] WLB[245] WLB[244]
+WLB[243] WLB[242] WLB[241] WLB[240] WLB[239] WLB[238] WLB[237] WLB[236] WLB[235] WLB[234]
+WLB[233] WLB[232] WLB[231] WLB[230] WLB[229] WLB[228] WLB[227] WLB[226] WLB[225] WLB[224]
+WLB[223] WLB[222] WLB[221] WLB[220] WLB[219] WLB[218] WLB[217] WLB[216] WLB[215] WLB[214]
+WLB[213] WLB[212] WLB[211] WLB[210] WLB[209] WLB[208] WLB[207] WLB[206] WLB[205] WLB[204]
+WLB[203] WLB[202] WLB[201] WLB[200] WLB[199] WLB[198] WLB[197] WLB[196] WLB[195] WLB[194]
+WLB[193] WLB[192] WLB[191] WLB[190] WLB[189] WLB[188] WLB[187] WLB[186] WLB[185] WLB[184]
+WLB[183] WLB[182] WLB[181] WLB[180] WLB[179] WLB[178] WLB[177] WLB[176] WLB[175] WLB[174]
+WLB[173] WLB[172] WLB[171] WLB[170] WLB[169] WLB[168] WLB[167] WLB[166] WLB[165] WLB[164]
+WLB[163] WLB[162] WLB[161] WLB[160] WLB[159] WLB[158] WLB[157] WLB[156] WLB[155] WLB[154]
+WLB[153] WLB[152] WLB[151] WLB[150] WLB[149] WLB[148] WLB[147] WLB[146] WLB[145] WLB[144]
+WLB[143] WLB[142] WLB[141] WLB[140] WLB[139] WLB[138] WLB[137] WLB[136] WLB[135] WLB[134]
+WLB[133] WLB[132] WLB[131] WLB[130] WLB[129] WLB[128] WLB[127] WLB[126] WLB[125] WLB[124]
+WLB[123] WLB[122] WLB[121] WLB[120] WLB[119] WLB[118] WLB[117] WLB[116] WLB[115] WLB[114]
+WLB[113] WLB[112] WLB[111] WLB[110] WLB[109] WLB[108] WLB[107] WLB[106] WLB[105] WLB[104]
+WLB[103] WLB[102] WLB[101] WLB[100] WLB[99] WLB[98] WLB[97] WLB[96] WLB[95] WLB[94]
+WLB[93] WLB[92] WLB[91] WLB[90] WLB[89] WLB[88] WLB[87] WLB[86] WLB[85] WLB[84]
+WLB[83] WLB[82] WLB[81] WLB[80] WLB[79] WLB[78] WLB[77] WLB[76] WLB[75] WLB[74]
+WLB[73] WLB[72] WLB[71] WLB[70] WLB[69] WLB[68] WLB[67] WLB[66] WLB[65] WLB[64]
+WLB[63] WLB[62] WLB[61] WLB[60] WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54]
+WLB[53] WLB[52] WLB[51] WLB[50] WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44]
+WLB[43] WLB[42] WLB[41] WLB[40] WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34]
+WLB[33] WLB[32] WLB[31] WLB[30] WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24]
+WLB[23] WLB[22] WLB[21] WLB[20] WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14]
+WLB[13] WLB[12] WLB[11] WLB[10] WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4]
+WLB[3] WLB[2] WLB[1] WLB[0] YXA[7] YXA[6] YXA[5] YXA[4] YXA[3] YXA[2]
+YXA[1] YXA[0] YXB[7] YXB[6] YXB[5] YXB[4] YXB[3] YXB[2] YXB[1] YXB[0] S55NLLGDPH_X512Y8D16_BW_Y512X8CELL_BW
XI21 BWENA[5] BWENB[5] CLKA CLKB CLKXA CLKXB DATAA[5] DATAB[5] DOUTA[5] DOUTB[5]
+VSS VSS VSS VSS STWLB VSS VSS VSS RWLA[0] RWLA[1]
+RWLB[0] RWLB[1] SACK1A SACK1B SACK4A SACK4B VDD VSS WEA WEB
+WLA[511] WLA[510] WLA[509] WLA[508] WLA[507] WLA[506] WLA[505] WLA[504] WLA[503] WLA[502]
+WLA[501] WLA[500] WLA[499] WLA[498] WLA[497] WLA[496] WLA[495] WLA[494] WLA[493] WLA[492]
+WLA[491] WLA[490] WLA[489] WLA[488] WLA[487] WLA[486] WLA[485] WLA[484] WLA[483] WLA[482]
+WLA[481] WLA[480] WLA[479] WLA[478] WLA[477] WLA[476] WLA[475] WLA[474] WLA[473] WLA[472]
+WLA[471] WLA[470] WLA[469] WLA[468] WLA[467] WLA[466] WLA[465] WLA[464] WLA[463] WLA[462]
+WLA[461] WLA[460] WLA[459] WLA[458] WLA[457] WLA[456] WLA[455] WLA[454] WLA[453] WLA[452]
+WLA[451] WLA[450] WLA[449] WLA[448] WLA[447] WLA[446] WLA[445] WLA[444] WLA[443] WLA[442]
+WLA[441] WLA[440] WLA[439] WLA[438] WLA[437] WLA[436] WLA[435] WLA[434] WLA[433] WLA[432]
+WLA[431] WLA[430] WLA[429] WLA[428] WLA[427] WLA[426] WLA[425] WLA[424] WLA[423] WLA[422]
+WLA[421] WLA[420] WLA[419] WLA[418] WLA[417] WLA[416] WLA[415] WLA[414] WLA[413] WLA[412]
+WLA[411] WLA[410] WLA[409] WLA[408] WLA[407] WLA[406] WLA[405] WLA[404] WLA[403] WLA[402]
+WLA[401] WLA[400] WLA[399] WLA[398] WLA[397] WLA[396] WLA[395] WLA[394] WLA[393] WLA[392]
+WLA[391] WLA[390] WLA[389] WLA[388] WLA[387] WLA[386] WLA[385] WLA[384] WLA[383] WLA[382]
+WLA[381] WLA[380] WLA[379] WLA[378] WLA[377] WLA[376] WLA[375] WLA[374] WLA[373] WLA[372]
+WLA[371] WLA[370] WLA[369] WLA[368] WLA[367] WLA[366] WLA[365] WLA[364] WLA[363] WLA[362]
+WLA[361] WLA[360] WLA[359] WLA[358] WLA[357] WLA[356] WLA[355] WLA[354] WLA[353] WLA[352]
+WLA[351] WLA[350] WLA[349] WLA[348] WLA[347] WLA[346] WLA[345] WLA[344] WLA[343] WLA[342]
+WLA[341] WLA[340] WLA[339] WLA[338] WLA[337] WLA[336] WLA[335] WLA[334] WLA[333] WLA[332]
+WLA[331] WLA[330] WLA[329] WLA[328] WLA[327] WLA[326] WLA[325] WLA[324] WLA[323] WLA[322]
+WLA[321] WLA[320] WLA[319] WLA[318] WLA[317] WLA[316] WLA[315] WLA[314] WLA[313] WLA[312]
+WLA[311] WLA[310] WLA[309] WLA[308] WLA[307] WLA[306] WLA[305] WLA[304] WLA[303] WLA[302]
+WLA[301] WLA[300] WLA[299] WLA[298] WLA[297] WLA[296] WLA[295] WLA[294] WLA[293] WLA[292]
+WLA[291] WLA[290] WLA[289] WLA[288] WLA[287] WLA[286] WLA[285] WLA[284] WLA[283] WLA[282]
+WLA[281] WLA[280] WLA[279] WLA[278] WLA[277] WLA[276] WLA[275] WLA[274] WLA[273] WLA[272]
+WLA[271] WLA[270] WLA[269] WLA[268] WLA[267] WLA[266] WLA[265] WLA[264] WLA[263] WLA[262]
+WLA[261] WLA[260] WLA[259] WLA[258] WLA[257] WLA[256] WLA[255] WLA[254] WLA[253] WLA[252]
+WLA[251] WLA[250] WLA[249] WLA[248] WLA[247] WLA[246] WLA[245] WLA[244] WLA[243] WLA[242]
+WLA[241] WLA[240] WLA[239] WLA[238] WLA[237] WLA[236] WLA[235] WLA[234] WLA[233] WLA[232]
+WLA[231] WLA[230] WLA[229] WLA[228] WLA[227] WLA[226] WLA[225] WLA[224] WLA[223] WLA[222]
+WLA[221] WLA[220] WLA[219] WLA[218] WLA[217] WLA[216] WLA[215] WLA[214] WLA[213] WLA[212]
+WLA[211] WLA[210] WLA[209] WLA[208] WLA[207] WLA[206] WLA[205] WLA[204] WLA[203] WLA[202]
+WLA[201] WLA[200] WLA[199] WLA[198] WLA[197] WLA[196] WLA[195] WLA[194] WLA[193] WLA[192]
+WLA[191] WLA[190] WLA[189] WLA[188] WLA[187] WLA[186] WLA[185] WLA[184] WLA[183] WLA[182]
+WLA[181] WLA[180] WLA[179] WLA[178] WLA[177] WLA[176] WLA[175] WLA[174] WLA[173] WLA[172]
+WLA[171] WLA[170] WLA[169] WLA[168] WLA[167] WLA[166] WLA[165] WLA[164] WLA[163] WLA[162]
+WLA[161] WLA[160] WLA[159] WLA[158] WLA[157] WLA[156] WLA[155] WLA[154] WLA[153] WLA[152]
+WLA[151] WLA[150] WLA[149] WLA[148] WLA[147] WLA[146] WLA[145] WLA[144] WLA[143] WLA[142]
+WLA[141] WLA[140] WLA[139] WLA[138] WLA[137] WLA[136] WLA[135] WLA[134] WLA[133] WLA[132]
+WLA[131] WLA[130] WLA[129] WLA[128] WLA[127] WLA[126] WLA[125] WLA[124] WLA[123] WLA[122]
+WLA[121] WLA[120] WLA[119] WLA[118] WLA[117] WLA[116] WLA[115] WLA[114] WLA[113] WLA[112]
+WLA[111] WLA[110] WLA[109] WLA[108] WLA[107] WLA[106] WLA[105] WLA[104] WLA[103] WLA[102]
+WLA[101] WLA[100] WLA[99] WLA[98] WLA[97] WLA[96] WLA[95] WLA[94] WLA[93] WLA[92]
+WLA[91] WLA[90] WLA[89] WLA[88] WLA[87] WLA[86] WLA[85] WLA[84] WLA[83] WLA[82]
+WLA[81] WLA[80] WLA[79] WLA[78] WLA[77] WLA[76] WLA[75] WLA[74] WLA[73] WLA[72]
+WLA[71] WLA[70] WLA[69] WLA[68] WLA[67] WLA[66] WLA[65] WLA[64] WLA[63] WLA[62]
+WLA[61] WLA[60] WLA[59] WLA[58] WLA[57] WLA[56] WLA[55] WLA[54] WLA[53] WLA[52]
+WLA[51] WLA[50] WLA[49] WLA[48] WLA[47] WLA[46] WLA[45] WLA[44] WLA[43] WLA[42]
+WLA[41] WLA[40] WLA[39] WLA[38] WLA[37] WLA[36] WLA[35] WLA[34] WLA[33] WLA[32]
+WLA[31] WLA[30] WLA[29] WLA[28] WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22]
+WLA[21] WLA[20] WLA[19] WLA[18] WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12]
+WLA[11] WLA[10] WLA[9] WLA[8] WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2]
+WLA[1] WLA[0] WLB[511] WLB[510] WLB[509] WLB[508] WLB[507] WLB[506] WLB[505] WLB[504]
+WLB[503] WLB[502] WLB[501] WLB[500] WLB[499] WLB[498] WLB[497] WLB[496] WLB[495] WLB[494]
+WLB[493] WLB[492] WLB[491] WLB[490] WLB[489] WLB[488] WLB[487] WLB[486] WLB[485] WLB[484]
+WLB[483] WLB[482] WLB[481] WLB[480] WLB[479] WLB[478] WLB[477] WLB[476] WLB[475] WLB[474]
+WLB[473] WLB[472] WLB[471] WLB[470] WLB[469] WLB[468] WLB[467] WLB[466] WLB[465] WLB[464]
+WLB[463] WLB[462] WLB[461] WLB[460] WLB[459] WLB[458] WLB[457] WLB[456] WLB[455] WLB[454]
+WLB[453] WLB[452] WLB[451] WLB[450] WLB[449] WLB[448] WLB[447] WLB[446] WLB[445] WLB[444]
+WLB[443] WLB[442] WLB[441] WLB[440] WLB[439] WLB[438] WLB[437] WLB[436] WLB[435] WLB[434]
+WLB[433] WLB[432] WLB[431] WLB[430] WLB[429] WLB[428] WLB[427] WLB[426] WLB[425] WLB[424]
+WLB[423] WLB[422] WLB[421] WLB[420] WLB[419] WLB[418] WLB[417] WLB[416] WLB[415] WLB[414]
+WLB[413] WLB[412] WLB[411] WLB[410] WLB[409] WLB[408] WLB[407] WLB[406] WLB[405] WLB[404]
+WLB[403] WLB[402] WLB[401] WLB[400] WLB[399] WLB[398] WLB[397] WLB[396] WLB[395] WLB[394]
+WLB[393] WLB[392] WLB[391] WLB[390] WLB[389] WLB[388] WLB[387] WLB[386] WLB[385] WLB[384]
+WLB[383] WLB[382] WLB[381] WLB[380] WLB[379] WLB[378] WLB[377] WLB[376] WLB[375] WLB[374]
+WLB[373] WLB[372] WLB[371] WLB[370] WLB[369] WLB[368] WLB[367] WLB[366] WLB[365] WLB[364]
+WLB[363] WLB[362] WLB[361] WLB[360] WLB[359] WLB[358] WLB[357] WLB[356] WLB[355] WLB[354]
+WLB[353] WLB[352] WLB[351] WLB[350] WLB[349] WLB[348] WLB[347] WLB[346] WLB[345] WLB[344]
+WLB[343] WLB[342] WLB[341] WLB[340] WLB[339] WLB[338] WLB[337] WLB[336] WLB[335] WLB[334]
+WLB[333] WLB[332] WLB[331] WLB[330] WLB[329] WLB[328] WLB[327] WLB[326] WLB[325] WLB[324]
+WLB[323] WLB[322] WLB[321] WLB[320] WLB[319] WLB[318] WLB[317] WLB[316] WLB[315] WLB[314]
+WLB[313] WLB[312] WLB[311] WLB[310] WLB[309] WLB[308] WLB[307] WLB[306] WLB[305] WLB[304]
+WLB[303] WLB[302] WLB[301] WLB[300] WLB[299] WLB[298] WLB[297] WLB[296] WLB[295] WLB[294]
+WLB[293] WLB[292] WLB[291] WLB[290] WLB[289] WLB[288] WLB[287] WLB[286] WLB[285] WLB[284]
+WLB[283] WLB[282] WLB[281] WLB[280] WLB[279] WLB[278] WLB[277] WLB[276] WLB[275] WLB[274]
+WLB[273] WLB[272] WLB[271] WLB[270] WLB[269] WLB[268] WLB[267] WLB[266] WLB[265] WLB[264]
+WLB[263] WLB[262] WLB[261] WLB[260] WLB[259] WLB[258] WLB[257] WLB[256] WLB[255] WLB[254]
+WLB[253] WLB[252] WLB[251] WLB[250] WLB[249] WLB[248] WLB[247] WLB[246] WLB[245] WLB[244]
+WLB[243] WLB[242] WLB[241] WLB[240] WLB[239] WLB[238] WLB[237] WLB[236] WLB[235] WLB[234]
+WLB[233] WLB[232] WLB[231] WLB[230] WLB[229] WLB[228] WLB[227] WLB[226] WLB[225] WLB[224]
+WLB[223] WLB[222] WLB[221] WLB[220] WLB[219] WLB[218] WLB[217] WLB[216] WLB[215] WLB[214]
+WLB[213] WLB[212] WLB[211] WLB[210] WLB[209] WLB[208] WLB[207] WLB[206] WLB[205] WLB[204]
+WLB[203] WLB[202] WLB[201] WLB[200] WLB[199] WLB[198] WLB[197] WLB[196] WLB[195] WLB[194]
+WLB[193] WLB[192] WLB[191] WLB[190] WLB[189] WLB[188] WLB[187] WLB[186] WLB[185] WLB[184]
+WLB[183] WLB[182] WLB[181] WLB[180] WLB[179] WLB[178] WLB[177] WLB[176] WLB[175] WLB[174]
+WLB[173] WLB[172] WLB[171] WLB[170] WLB[169] WLB[168] WLB[167] WLB[166] WLB[165] WLB[164]
+WLB[163] WLB[162] WLB[161] WLB[160] WLB[159] WLB[158] WLB[157] WLB[156] WLB[155] WLB[154]
+WLB[153] WLB[152] WLB[151] WLB[150] WLB[149] WLB[148] WLB[147] WLB[146] WLB[145] WLB[144]
+WLB[143] WLB[142] WLB[141] WLB[140] WLB[139] WLB[138] WLB[137] WLB[136] WLB[135] WLB[134]
+WLB[133] WLB[132] WLB[131] WLB[130] WLB[129] WLB[128] WLB[127] WLB[126] WLB[125] WLB[124]
+WLB[123] WLB[122] WLB[121] WLB[120] WLB[119] WLB[118] WLB[117] WLB[116] WLB[115] WLB[114]
+WLB[113] WLB[112] WLB[111] WLB[110] WLB[109] WLB[108] WLB[107] WLB[106] WLB[105] WLB[104]
+WLB[103] WLB[102] WLB[101] WLB[100] WLB[99] WLB[98] WLB[97] WLB[96] WLB[95] WLB[94]
+WLB[93] WLB[92] WLB[91] WLB[90] WLB[89] WLB[88] WLB[87] WLB[86] WLB[85] WLB[84]
+WLB[83] WLB[82] WLB[81] WLB[80] WLB[79] WLB[78] WLB[77] WLB[76] WLB[75] WLB[74]
+WLB[73] WLB[72] WLB[71] WLB[70] WLB[69] WLB[68] WLB[67] WLB[66] WLB[65] WLB[64]
+WLB[63] WLB[62] WLB[61] WLB[60] WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54]
+WLB[53] WLB[52] WLB[51] WLB[50] WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44]
+WLB[43] WLB[42] WLB[41] WLB[40] WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34]
+WLB[33] WLB[32] WLB[31] WLB[30] WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24]
+WLB[23] WLB[22] WLB[21] WLB[20] WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14]
+WLB[13] WLB[12] WLB[11] WLB[10] WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4]
+WLB[3] WLB[2] WLB[1] WLB[0] YXA[7] YXA[6] YXA[5] YXA[4] YXA[3] YXA[2]
+YXA[1] YXA[0] YXB[7] YXB[6] YXB[5] YXB[4] YXB[3] YXB[2] YXB[1] YXB[0] S55NLLGDPH_X512Y8D16_BW_Y512X8CELL_BW
XI22 BWENA[6] BWENB[6] CLKA CLKB CLKXA CLKXB DATAA[6] DATAB[6] DOUTA[6] DOUTB[6]
+VSS VSS VSS VSS STWLB VSS VSS VSS RWLA[0] RWLA[1]
+RWLB[0] RWLB[1] SACK1A SACK1B SACK4A SACK4B VDD VSS WEA WEB
+WLA[511] WLA[510] WLA[509] WLA[508] WLA[507] WLA[506] WLA[505] WLA[504] WLA[503] WLA[502]
+WLA[501] WLA[500] WLA[499] WLA[498] WLA[497] WLA[496] WLA[495] WLA[494] WLA[493] WLA[492]
+WLA[491] WLA[490] WLA[489] WLA[488] WLA[487] WLA[486] WLA[485] WLA[484] WLA[483] WLA[482]
+WLA[481] WLA[480] WLA[479] WLA[478] WLA[477] WLA[476] WLA[475] WLA[474] WLA[473] WLA[472]
+WLA[471] WLA[470] WLA[469] WLA[468] WLA[467] WLA[466] WLA[465] WLA[464] WLA[463] WLA[462]
+WLA[461] WLA[460] WLA[459] WLA[458] WLA[457] WLA[456] WLA[455] WLA[454] WLA[453] WLA[452]
+WLA[451] WLA[450] WLA[449] WLA[448] WLA[447] WLA[446] WLA[445] WLA[444] WLA[443] WLA[442]
+WLA[441] WLA[440] WLA[439] WLA[438] WLA[437] WLA[436] WLA[435] WLA[434] WLA[433] WLA[432]
+WLA[431] WLA[430] WLA[429] WLA[428] WLA[427] WLA[426] WLA[425] WLA[424] WLA[423] WLA[422]
+WLA[421] WLA[420] WLA[419] WLA[418] WLA[417] WLA[416] WLA[415] WLA[414] WLA[413] WLA[412]
+WLA[411] WLA[410] WLA[409] WLA[408] WLA[407] WLA[406] WLA[405] WLA[404] WLA[403] WLA[402]
+WLA[401] WLA[400] WLA[399] WLA[398] WLA[397] WLA[396] WLA[395] WLA[394] WLA[393] WLA[392]
+WLA[391] WLA[390] WLA[389] WLA[388] WLA[387] WLA[386] WLA[385] WLA[384] WLA[383] WLA[382]
+WLA[381] WLA[380] WLA[379] WLA[378] WLA[377] WLA[376] WLA[375] WLA[374] WLA[373] WLA[372]
+WLA[371] WLA[370] WLA[369] WLA[368] WLA[367] WLA[366] WLA[365] WLA[364] WLA[363] WLA[362]
+WLA[361] WLA[360] WLA[359] WLA[358] WLA[357] WLA[356] WLA[355] WLA[354] WLA[353] WLA[352]
+WLA[351] WLA[350] WLA[349] WLA[348] WLA[347] WLA[346] WLA[345] WLA[344] WLA[343] WLA[342]
+WLA[341] WLA[340] WLA[339] WLA[338] WLA[337] WLA[336] WLA[335] WLA[334] WLA[333] WLA[332]
+WLA[331] WLA[330] WLA[329] WLA[328] WLA[327] WLA[326] WLA[325] WLA[324] WLA[323] WLA[322]
+WLA[321] WLA[320] WLA[319] WLA[318] WLA[317] WLA[316] WLA[315] WLA[314] WLA[313] WLA[312]
+WLA[311] WLA[310] WLA[309] WLA[308] WLA[307] WLA[306] WLA[305] WLA[304] WLA[303] WLA[302]
+WLA[301] WLA[300] WLA[299] WLA[298] WLA[297] WLA[296] WLA[295] WLA[294] WLA[293] WLA[292]
+WLA[291] WLA[290] WLA[289] WLA[288] WLA[287] WLA[286] WLA[285] WLA[284] WLA[283] WLA[282]
+WLA[281] WLA[280] WLA[279] WLA[278] WLA[277] WLA[276] WLA[275] WLA[274] WLA[273] WLA[272]
+WLA[271] WLA[270] WLA[269] WLA[268] WLA[267] WLA[266] WLA[265] WLA[264] WLA[263] WLA[262]
+WLA[261] WLA[260] WLA[259] WLA[258] WLA[257] WLA[256] WLA[255] WLA[254] WLA[253] WLA[252]
+WLA[251] WLA[250] WLA[249] WLA[248] WLA[247] WLA[246] WLA[245] WLA[244] WLA[243] WLA[242]
+WLA[241] WLA[240] WLA[239] WLA[238] WLA[237] WLA[236] WLA[235] WLA[234] WLA[233] WLA[232]
+WLA[231] WLA[230] WLA[229] WLA[228] WLA[227] WLA[226] WLA[225] WLA[224] WLA[223] WLA[222]
+WLA[221] WLA[220] WLA[219] WLA[218] WLA[217] WLA[216] WLA[215] WLA[214] WLA[213] WLA[212]
+WLA[211] WLA[210] WLA[209] WLA[208] WLA[207] WLA[206] WLA[205] WLA[204] WLA[203] WLA[202]
+WLA[201] WLA[200] WLA[199] WLA[198] WLA[197] WLA[196] WLA[195] WLA[194] WLA[193] WLA[192]
+WLA[191] WLA[190] WLA[189] WLA[188] WLA[187] WLA[186] WLA[185] WLA[184] WLA[183] WLA[182]
+WLA[181] WLA[180] WLA[179] WLA[178] WLA[177] WLA[176] WLA[175] WLA[174] WLA[173] WLA[172]
+WLA[171] WLA[170] WLA[169] WLA[168] WLA[167] WLA[166] WLA[165] WLA[164] WLA[163] WLA[162]
+WLA[161] WLA[160] WLA[159] WLA[158] WLA[157] WLA[156] WLA[155] WLA[154] WLA[153] WLA[152]
+WLA[151] WLA[150] WLA[149] WLA[148] WLA[147] WLA[146] WLA[145] WLA[144] WLA[143] WLA[142]
+WLA[141] WLA[140] WLA[139] WLA[138] WLA[137] WLA[136] WLA[135] WLA[134] WLA[133] WLA[132]
+WLA[131] WLA[130] WLA[129] WLA[128] WLA[127] WLA[126] WLA[125] WLA[124] WLA[123] WLA[122]
+WLA[121] WLA[120] WLA[119] WLA[118] WLA[117] WLA[116] WLA[115] WLA[114] WLA[113] WLA[112]
+WLA[111] WLA[110] WLA[109] WLA[108] WLA[107] WLA[106] WLA[105] WLA[104] WLA[103] WLA[102]
+WLA[101] WLA[100] WLA[99] WLA[98] WLA[97] WLA[96] WLA[95] WLA[94] WLA[93] WLA[92]
+WLA[91] WLA[90] WLA[89] WLA[88] WLA[87] WLA[86] WLA[85] WLA[84] WLA[83] WLA[82]
+WLA[81] WLA[80] WLA[79] WLA[78] WLA[77] WLA[76] WLA[75] WLA[74] WLA[73] WLA[72]
+WLA[71] WLA[70] WLA[69] WLA[68] WLA[67] WLA[66] WLA[65] WLA[64] WLA[63] WLA[62]
+WLA[61] WLA[60] WLA[59] WLA[58] WLA[57] WLA[56] WLA[55] WLA[54] WLA[53] WLA[52]
+WLA[51] WLA[50] WLA[49] WLA[48] WLA[47] WLA[46] WLA[45] WLA[44] WLA[43] WLA[42]
+WLA[41] WLA[40] WLA[39] WLA[38] WLA[37] WLA[36] WLA[35] WLA[34] WLA[33] WLA[32]
+WLA[31] WLA[30] WLA[29] WLA[28] WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22]
+WLA[21] WLA[20] WLA[19] WLA[18] WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12]
+WLA[11] WLA[10] WLA[9] WLA[8] WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2]
+WLA[1] WLA[0] WLB[511] WLB[510] WLB[509] WLB[508] WLB[507] WLB[506] WLB[505] WLB[504]
+WLB[503] WLB[502] WLB[501] WLB[500] WLB[499] WLB[498] WLB[497] WLB[496] WLB[495] WLB[494]
+WLB[493] WLB[492] WLB[491] WLB[490] WLB[489] WLB[488] WLB[487] WLB[486] WLB[485] WLB[484]
+WLB[483] WLB[482] WLB[481] WLB[480] WLB[479] WLB[478] WLB[477] WLB[476] WLB[475] WLB[474]
+WLB[473] WLB[472] WLB[471] WLB[470] WLB[469] WLB[468] WLB[467] WLB[466] WLB[465] WLB[464]
+WLB[463] WLB[462] WLB[461] WLB[460] WLB[459] WLB[458] WLB[457] WLB[456] WLB[455] WLB[454]
+WLB[453] WLB[452] WLB[451] WLB[450] WLB[449] WLB[448] WLB[447] WLB[446] WLB[445] WLB[444]
+WLB[443] WLB[442] WLB[441] WLB[440] WLB[439] WLB[438] WLB[437] WLB[436] WLB[435] WLB[434]
+WLB[433] WLB[432] WLB[431] WLB[430] WLB[429] WLB[428] WLB[427] WLB[426] WLB[425] WLB[424]
+WLB[423] WLB[422] WLB[421] WLB[420] WLB[419] WLB[418] WLB[417] WLB[416] WLB[415] WLB[414]
+WLB[413] WLB[412] WLB[411] WLB[410] WLB[409] WLB[408] WLB[407] WLB[406] WLB[405] WLB[404]
+WLB[403] WLB[402] WLB[401] WLB[400] WLB[399] WLB[398] WLB[397] WLB[396] WLB[395] WLB[394]
+WLB[393] WLB[392] WLB[391] WLB[390] WLB[389] WLB[388] WLB[387] WLB[386] WLB[385] WLB[384]
+WLB[383] WLB[382] WLB[381] WLB[380] WLB[379] WLB[378] WLB[377] WLB[376] WLB[375] WLB[374]
+WLB[373] WLB[372] WLB[371] WLB[370] WLB[369] WLB[368] WLB[367] WLB[366] WLB[365] WLB[364]
+WLB[363] WLB[362] WLB[361] WLB[360] WLB[359] WLB[358] WLB[357] WLB[356] WLB[355] WLB[354]
+WLB[353] WLB[352] WLB[351] WLB[350] WLB[349] WLB[348] WLB[347] WLB[346] WLB[345] WLB[344]
+WLB[343] WLB[342] WLB[341] WLB[340] WLB[339] WLB[338] WLB[337] WLB[336] WLB[335] WLB[334]
+WLB[333] WLB[332] WLB[331] WLB[330] WLB[329] WLB[328] WLB[327] WLB[326] WLB[325] WLB[324]
+WLB[323] WLB[322] WLB[321] WLB[320] WLB[319] WLB[318] WLB[317] WLB[316] WLB[315] WLB[314]
+WLB[313] WLB[312] WLB[311] WLB[310] WLB[309] WLB[308] WLB[307] WLB[306] WLB[305] WLB[304]
+WLB[303] WLB[302] WLB[301] WLB[300] WLB[299] WLB[298] WLB[297] WLB[296] WLB[295] WLB[294]
+WLB[293] WLB[292] WLB[291] WLB[290] WLB[289] WLB[288] WLB[287] WLB[286] WLB[285] WLB[284]
+WLB[283] WLB[282] WLB[281] WLB[280] WLB[279] WLB[278] WLB[277] WLB[276] WLB[275] WLB[274]
+WLB[273] WLB[272] WLB[271] WLB[270] WLB[269] WLB[268] WLB[267] WLB[266] WLB[265] WLB[264]
+WLB[263] WLB[262] WLB[261] WLB[260] WLB[259] WLB[258] WLB[257] WLB[256] WLB[255] WLB[254]
+WLB[253] WLB[252] WLB[251] WLB[250] WLB[249] WLB[248] WLB[247] WLB[246] WLB[245] WLB[244]
+WLB[243] WLB[242] WLB[241] WLB[240] WLB[239] WLB[238] WLB[237] WLB[236] WLB[235] WLB[234]
+WLB[233] WLB[232] WLB[231] WLB[230] WLB[229] WLB[228] WLB[227] WLB[226] WLB[225] WLB[224]
+WLB[223] WLB[222] WLB[221] WLB[220] WLB[219] WLB[218] WLB[217] WLB[216] WLB[215] WLB[214]
+WLB[213] WLB[212] WLB[211] WLB[210] WLB[209] WLB[208] WLB[207] WLB[206] WLB[205] WLB[204]
+WLB[203] WLB[202] WLB[201] WLB[200] WLB[199] WLB[198] WLB[197] WLB[196] WLB[195] WLB[194]
+WLB[193] WLB[192] WLB[191] WLB[190] WLB[189] WLB[188] WLB[187] WLB[186] WLB[185] WLB[184]
+WLB[183] WLB[182] WLB[181] WLB[180] WLB[179] WLB[178] WLB[177] WLB[176] WLB[175] WLB[174]
+WLB[173] WLB[172] WLB[171] WLB[170] WLB[169] WLB[168] WLB[167] WLB[166] WLB[165] WLB[164]
+WLB[163] WLB[162] WLB[161] WLB[160] WLB[159] WLB[158] WLB[157] WLB[156] WLB[155] WLB[154]
+WLB[153] WLB[152] WLB[151] WLB[150] WLB[149] WLB[148] WLB[147] WLB[146] WLB[145] WLB[144]
+WLB[143] WLB[142] WLB[141] WLB[140] WLB[139] WLB[138] WLB[137] WLB[136] WLB[135] WLB[134]
+WLB[133] WLB[132] WLB[131] WLB[130] WLB[129] WLB[128] WLB[127] WLB[126] WLB[125] WLB[124]
+WLB[123] WLB[122] WLB[121] WLB[120] WLB[119] WLB[118] WLB[117] WLB[116] WLB[115] WLB[114]
+WLB[113] WLB[112] WLB[111] WLB[110] WLB[109] WLB[108] WLB[107] WLB[106] WLB[105] WLB[104]
+WLB[103] WLB[102] WLB[101] WLB[100] WLB[99] WLB[98] WLB[97] WLB[96] WLB[95] WLB[94]
+WLB[93] WLB[92] WLB[91] WLB[90] WLB[89] WLB[88] WLB[87] WLB[86] WLB[85] WLB[84]
+WLB[83] WLB[82] WLB[81] WLB[80] WLB[79] WLB[78] WLB[77] WLB[76] WLB[75] WLB[74]
+WLB[73] WLB[72] WLB[71] WLB[70] WLB[69] WLB[68] WLB[67] WLB[66] WLB[65] WLB[64]
+WLB[63] WLB[62] WLB[61] WLB[60] WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54]
+WLB[53] WLB[52] WLB[51] WLB[50] WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44]
+WLB[43] WLB[42] WLB[41] WLB[40] WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34]
+WLB[33] WLB[32] WLB[31] WLB[30] WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24]
+WLB[23] WLB[22] WLB[21] WLB[20] WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14]
+WLB[13] WLB[12] WLB[11] WLB[10] WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4]
+WLB[3] WLB[2] WLB[1] WLB[0] YXA[7] YXA[6] YXA[5] YXA[4] YXA[3] YXA[2]
+YXA[1] YXA[0] YXB[7] YXB[6] YXB[5] YXB[4] YXB[3] YXB[2] YXB[1] YXB[0] S55NLLGDPH_X512Y8D16_BW_Y512X8CELL_BW
XI23 BWENA[7] BWENB[7] CLKA CLKB CLKXA CLKXB DATAA[7] DATAB[7] DOUTA[7] DOUTB[7]
+VSS VSS VSS VSS STWLB VSS VSS VSS RWLA[0] RWLA[1]
+RWLB[0] RWLB[1] SACK1A SACK1B SACK4A SACK4B VDD VSS WEA WEB
+WLA[511] WLA[510] WLA[509] WLA[508] WLA[507] WLA[506] WLA[505] WLA[504] WLA[503] WLA[502]
+WLA[501] WLA[500] WLA[499] WLA[498] WLA[497] WLA[496] WLA[495] WLA[494] WLA[493] WLA[492]
+WLA[491] WLA[490] WLA[489] WLA[488] WLA[487] WLA[486] WLA[485] WLA[484] WLA[483] WLA[482]
+WLA[481] WLA[480] WLA[479] WLA[478] WLA[477] WLA[476] WLA[475] WLA[474] WLA[473] WLA[472]
+WLA[471] WLA[470] WLA[469] WLA[468] WLA[467] WLA[466] WLA[465] WLA[464] WLA[463] WLA[462]
+WLA[461] WLA[460] WLA[459] WLA[458] WLA[457] WLA[456] WLA[455] WLA[454] WLA[453] WLA[452]
+WLA[451] WLA[450] WLA[449] WLA[448] WLA[447] WLA[446] WLA[445] WLA[444] WLA[443] WLA[442]
+WLA[441] WLA[440] WLA[439] WLA[438] WLA[437] WLA[436] WLA[435] WLA[434] WLA[433] WLA[432]
+WLA[431] WLA[430] WLA[429] WLA[428] WLA[427] WLA[426] WLA[425] WLA[424] WLA[423] WLA[422]
+WLA[421] WLA[420] WLA[419] WLA[418] WLA[417] WLA[416] WLA[415] WLA[414] WLA[413] WLA[412]
+WLA[411] WLA[410] WLA[409] WLA[408] WLA[407] WLA[406] WLA[405] WLA[404] WLA[403] WLA[402]
+WLA[401] WLA[400] WLA[399] WLA[398] WLA[397] WLA[396] WLA[395] WLA[394] WLA[393] WLA[392]
+WLA[391] WLA[390] WLA[389] WLA[388] WLA[387] WLA[386] WLA[385] WLA[384] WLA[383] WLA[382]
+WLA[381] WLA[380] WLA[379] WLA[378] WLA[377] WLA[376] WLA[375] WLA[374] WLA[373] WLA[372]
+WLA[371] WLA[370] WLA[369] WLA[368] WLA[367] WLA[366] WLA[365] WLA[364] WLA[363] WLA[362]
+WLA[361] WLA[360] WLA[359] WLA[358] WLA[357] WLA[356] WLA[355] WLA[354] WLA[353] WLA[352]
+WLA[351] WLA[350] WLA[349] WLA[348] WLA[347] WLA[346] WLA[345] WLA[344] WLA[343] WLA[342]
+WLA[341] WLA[340] WLA[339] WLA[338] WLA[337] WLA[336] WLA[335] WLA[334] WLA[333] WLA[332]
+WLA[331] WLA[330] WLA[329] WLA[328] WLA[327] WLA[326] WLA[325] WLA[324] WLA[323] WLA[322]
+WLA[321] WLA[320] WLA[319] WLA[318] WLA[317] WLA[316] WLA[315] WLA[314] WLA[313] WLA[312]
+WLA[311] WLA[310] WLA[309] WLA[308] WLA[307] WLA[306] WLA[305] WLA[304] WLA[303] WLA[302]
+WLA[301] WLA[300] WLA[299] WLA[298] WLA[297] WLA[296] WLA[295] WLA[294] WLA[293] WLA[292]
+WLA[291] WLA[290] WLA[289] WLA[288] WLA[287] WLA[286] WLA[285] WLA[284] WLA[283] WLA[282]
+WLA[281] WLA[280] WLA[279] WLA[278] WLA[277] WLA[276] WLA[275] WLA[274] WLA[273] WLA[272]
+WLA[271] WLA[270] WLA[269] WLA[268] WLA[267] WLA[266] WLA[265] WLA[264] WLA[263] WLA[262]
+WLA[261] WLA[260] WLA[259] WLA[258] WLA[257] WLA[256] WLA[255] WLA[254] WLA[253] WLA[252]
+WLA[251] WLA[250] WLA[249] WLA[248] WLA[247] WLA[246] WLA[245] WLA[244] WLA[243] WLA[242]
+WLA[241] WLA[240] WLA[239] WLA[238] WLA[237] WLA[236] WLA[235] WLA[234] WLA[233] WLA[232]
+WLA[231] WLA[230] WLA[229] WLA[228] WLA[227] WLA[226] WLA[225] WLA[224] WLA[223] WLA[222]
+WLA[221] WLA[220] WLA[219] WLA[218] WLA[217] WLA[216] WLA[215] WLA[214] WLA[213] WLA[212]
+WLA[211] WLA[210] WLA[209] WLA[208] WLA[207] WLA[206] WLA[205] WLA[204] WLA[203] WLA[202]
+WLA[201] WLA[200] WLA[199] WLA[198] WLA[197] WLA[196] WLA[195] WLA[194] WLA[193] WLA[192]
+WLA[191] WLA[190] WLA[189] WLA[188] WLA[187] WLA[186] WLA[185] WLA[184] WLA[183] WLA[182]
+WLA[181] WLA[180] WLA[179] WLA[178] WLA[177] WLA[176] WLA[175] WLA[174] WLA[173] WLA[172]
+WLA[171] WLA[170] WLA[169] WLA[168] WLA[167] WLA[166] WLA[165] WLA[164] WLA[163] WLA[162]
+WLA[161] WLA[160] WLA[159] WLA[158] WLA[157] WLA[156] WLA[155] WLA[154] WLA[153] WLA[152]
+WLA[151] WLA[150] WLA[149] WLA[148] WLA[147] WLA[146] WLA[145] WLA[144] WLA[143] WLA[142]
+WLA[141] WLA[140] WLA[139] WLA[138] WLA[137] WLA[136] WLA[135] WLA[134] WLA[133] WLA[132]
+WLA[131] WLA[130] WLA[129] WLA[128] WLA[127] WLA[126] WLA[125] WLA[124] WLA[123] WLA[122]
+WLA[121] WLA[120] WLA[119] WLA[118] WLA[117] WLA[116] WLA[115] WLA[114] WLA[113] WLA[112]
+WLA[111] WLA[110] WLA[109] WLA[108] WLA[107] WLA[106] WLA[105] WLA[104] WLA[103] WLA[102]
+WLA[101] WLA[100] WLA[99] WLA[98] WLA[97] WLA[96] WLA[95] WLA[94] WLA[93] WLA[92]
+WLA[91] WLA[90] WLA[89] WLA[88] WLA[87] WLA[86] WLA[85] WLA[84] WLA[83] WLA[82]
+WLA[81] WLA[80] WLA[79] WLA[78] WLA[77] WLA[76] WLA[75] WLA[74] WLA[73] WLA[72]
+WLA[71] WLA[70] WLA[69] WLA[68] WLA[67] WLA[66] WLA[65] WLA[64] WLA[63] WLA[62]
+WLA[61] WLA[60] WLA[59] WLA[58] WLA[57] WLA[56] WLA[55] WLA[54] WLA[53] WLA[52]
+WLA[51] WLA[50] WLA[49] WLA[48] WLA[47] WLA[46] WLA[45] WLA[44] WLA[43] WLA[42]
+WLA[41] WLA[40] WLA[39] WLA[38] WLA[37] WLA[36] WLA[35] WLA[34] WLA[33] WLA[32]
+WLA[31] WLA[30] WLA[29] WLA[28] WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22]
+WLA[21] WLA[20] WLA[19] WLA[18] WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12]
+WLA[11] WLA[10] WLA[9] WLA[8] WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2]
+WLA[1] WLA[0] WLB[511] WLB[510] WLB[509] WLB[508] WLB[507] WLB[506] WLB[505] WLB[504]
+WLB[503] WLB[502] WLB[501] WLB[500] WLB[499] WLB[498] WLB[497] WLB[496] WLB[495] WLB[494]
+WLB[493] WLB[492] WLB[491] WLB[490] WLB[489] WLB[488] WLB[487] WLB[486] WLB[485] WLB[484]
+WLB[483] WLB[482] WLB[481] WLB[480] WLB[479] WLB[478] WLB[477] WLB[476] WLB[475] WLB[474]
+WLB[473] WLB[472] WLB[471] WLB[470] WLB[469] WLB[468] WLB[467] WLB[466] WLB[465] WLB[464]
+WLB[463] WLB[462] WLB[461] WLB[460] WLB[459] WLB[458] WLB[457] WLB[456] WLB[455] WLB[454]
+WLB[453] WLB[452] WLB[451] WLB[450] WLB[449] WLB[448] WLB[447] WLB[446] WLB[445] WLB[444]
+WLB[443] WLB[442] WLB[441] WLB[440] WLB[439] WLB[438] WLB[437] WLB[436] WLB[435] WLB[434]
+WLB[433] WLB[432] WLB[431] WLB[430] WLB[429] WLB[428] WLB[427] WLB[426] WLB[425] WLB[424]
+WLB[423] WLB[422] WLB[421] WLB[420] WLB[419] WLB[418] WLB[417] WLB[416] WLB[415] WLB[414]
+WLB[413] WLB[412] WLB[411] WLB[410] WLB[409] WLB[408] WLB[407] WLB[406] WLB[405] WLB[404]
+WLB[403] WLB[402] WLB[401] WLB[400] WLB[399] WLB[398] WLB[397] WLB[396] WLB[395] WLB[394]
+WLB[393] WLB[392] WLB[391] WLB[390] WLB[389] WLB[388] WLB[387] WLB[386] WLB[385] WLB[384]
+WLB[383] WLB[382] WLB[381] WLB[380] WLB[379] WLB[378] WLB[377] WLB[376] WLB[375] WLB[374]
+WLB[373] WLB[372] WLB[371] WLB[370] WLB[369] WLB[368] WLB[367] WLB[366] WLB[365] WLB[364]
+WLB[363] WLB[362] WLB[361] WLB[360] WLB[359] WLB[358] WLB[357] WLB[356] WLB[355] WLB[354]
+WLB[353] WLB[352] WLB[351] WLB[350] WLB[349] WLB[348] WLB[347] WLB[346] WLB[345] WLB[344]
+WLB[343] WLB[342] WLB[341] WLB[340] WLB[339] WLB[338] WLB[337] WLB[336] WLB[335] WLB[334]
+WLB[333] WLB[332] WLB[331] WLB[330] WLB[329] WLB[328] WLB[327] WLB[326] WLB[325] WLB[324]
+WLB[323] WLB[322] WLB[321] WLB[320] WLB[319] WLB[318] WLB[317] WLB[316] WLB[315] WLB[314]
+WLB[313] WLB[312] WLB[311] WLB[310] WLB[309] WLB[308] WLB[307] WLB[306] WLB[305] WLB[304]
+WLB[303] WLB[302] WLB[301] WLB[300] WLB[299] WLB[298] WLB[297] WLB[296] WLB[295] WLB[294]
+WLB[293] WLB[292] WLB[291] WLB[290] WLB[289] WLB[288] WLB[287] WLB[286] WLB[285] WLB[284]
+WLB[283] WLB[282] WLB[281] WLB[280] WLB[279] WLB[278] WLB[277] WLB[276] WLB[275] WLB[274]
+WLB[273] WLB[272] WLB[271] WLB[270] WLB[269] WLB[268] WLB[267] WLB[266] WLB[265] WLB[264]
+WLB[263] WLB[262] WLB[261] WLB[260] WLB[259] WLB[258] WLB[257] WLB[256] WLB[255] WLB[254]
+WLB[253] WLB[252] WLB[251] WLB[250] WLB[249] WLB[248] WLB[247] WLB[246] WLB[245] WLB[244]
+WLB[243] WLB[242] WLB[241] WLB[240] WLB[239] WLB[238] WLB[237] WLB[236] WLB[235] WLB[234]
+WLB[233] WLB[232] WLB[231] WLB[230] WLB[229] WLB[228] WLB[227] WLB[226] WLB[225] WLB[224]
+WLB[223] WLB[222] WLB[221] WLB[220] WLB[219] WLB[218] WLB[217] WLB[216] WLB[215] WLB[214]
+WLB[213] WLB[212] WLB[211] WLB[210] WLB[209] WLB[208] WLB[207] WLB[206] WLB[205] WLB[204]
+WLB[203] WLB[202] WLB[201] WLB[200] WLB[199] WLB[198] WLB[197] WLB[196] WLB[195] WLB[194]
+WLB[193] WLB[192] WLB[191] WLB[190] WLB[189] WLB[188] WLB[187] WLB[186] WLB[185] WLB[184]
+WLB[183] WLB[182] WLB[181] WLB[180] WLB[179] WLB[178] WLB[177] WLB[176] WLB[175] WLB[174]
+WLB[173] WLB[172] WLB[171] WLB[170] WLB[169] WLB[168] WLB[167] WLB[166] WLB[165] WLB[164]
+WLB[163] WLB[162] WLB[161] WLB[160] WLB[159] WLB[158] WLB[157] WLB[156] WLB[155] WLB[154]
+WLB[153] WLB[152] WLB[151] WLB[150] WLB[149] WLB[148] WLB[147] WLB[146] WLB[145] WLB[144]
+WLB[143] WLB[142] WLB[141] WLB[140] WLB[139] WLB[138] WLB[137] WLB[136] WLB[135] WLB[134]
+WLB[133] WLB[132] WLB[131] WLB[130] WLB[129] WLB[128] WLB[127] WLB[126] WLB[125] WLB[124]
+WLB[123] WLB[122] WLB[121] WLB[120] WLB[119] WLB[118] WLB[117] WLB[116] WLB[115] WLB[114]
+WLB[113] WLB[112] WLB[111] WLB[110] WLB[109] WLB[108] WLB[107] WLB[106] WLB[105] WLB[104]
+WLB[103] WLB[102] WLB[101] WLB[100] WLB[99] WLB[98] WLB[97] WLB[96] WLB[95] WLB[94]
+WLB[93] WLB[92] WLB[91] WLB[90] WLB[89] WLB[88] WLB[87] WLB[86] WLB[85] WLB[84]
+WLB[83] WLB[82] WLB[81] WLB[80] WLB[79] WLB[78] WLB[77] WLB[76] WLB[75] WLB[74]
+WLB[73] WLB[72] WLB[71] WLB[70] WLB[69] WLB[68] WLB[67] WLB[66] WLB[65] WLB[64]
+WLB[63] WLB[62] WLB[61] WLB[60] WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54]
+WLB[53] WLB[52] WLB[51] WLB[50] WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44]
+WLB[43] WLB[42] WLB[41] WLB[40] WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34]
+WLB[33] WLB[32] WLB[31] WLB[30] WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24]
+WLB[23] WLB[22] WLB[21] WLB[20] WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14]
+WLB[13] WLB[12] WLB[11] WLB[10] WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4]
+WLB[3] WLB[2] WLB[1] WLB[0] YXA[7] YXA[6] YXA[5] YXA[4] YXA[3] YXA[2]
+YXA[1] YXA[0] YXB[7] YXB[6] YXB[5] YXB[4] YXB[3] YXB[2] YXB[1] YXB[0] S55NLLGDPH_X512Y8D16_BW_Y512X8CELL_BW
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    S55NLLGDPH_X512Y8D16_BW_EDGECELL66B_RED_RIGHT
* View Name:    schematic
************************************************************************

.SUBCKT S55NLLGDPH_X512Y8D16_BW_EDGECELL66B_RED_RIGHT RWL[0] RWL[1] VDD VSS WLA[63] WLA[62] WLA[61] WLA[60] WLA[59] WLA[58]
+WLA[57] WLA[56] WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48]
+WLA[47] WLA[46] WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38]
+WLA[37] WLA[36] WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28]
+WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18]
+WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8]
+WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0]
XI0 NET01 NET61 VDD VSS S55NLLGDPH_X512Y8D16_BW_BLSTRAP_B
XI1 NET01 NET31 NET61 NET91 VDD VSS RWL[0] S55NLLGDPH_X512Y8D16_BW_EDGECELL
XI2 NET02 NET31 NET62 NET91 VDD VSS RWL[1] S55NLLGDPH_X512Y8D16_BW_EDGECELL
XI3 NET02 NET32 NET62 NET92 VDD VSS WLA[7] WLA[6] WLA[5] WLA[4]
+WLA[3] WLA[2] WLA[1] WLA[0] S55NLLGDPH_X512Y8D16_BW_EDGECELL8B
XI4 NET03 NET32 NET63 NET92 VDD VSS WLA[15] WLA[14] WLA[13] WLA[12]
+WLA[11] WLA[10] WLA[9] WLA[8] S55NLLGDPH_X512Y8D16_BW_EDGECELL8B
XI5 NET03 NET33 NET63 NET93 VDD VSS WLA[23] WLA[22] WLA[21] WLA[20]
+WLA[19] WLA[18] WLA[17] WLA[16] S55NLLGDPH_X512Y8D16_BW_EDGECELL8B
XI6 NET04 NET33 NET64 NET93 VDD VSS WLA[31] WLA[30] WLA[29] WLA[28]
+WLA[27] WLA[26] WLA[25] WLA[24] S55NLLGDPH_X512Y8D16_BW_EDGECELL8B
XI7 NET04 NET34 NET64 NET94 VDD VSS WLA[39] WLA[38] WLA[37] WLA[36]
+WLA[35] WLA[34] WLA[33] WLA[32] S55NLLGDPH_X512Y8D16_BW_EDGECELL8B
XI8 NET05 NET34 NET65 NET94 VDD VSS WLA[47] WLA[46] WLA[45] WLA[44]
+WLA[43] WLA[42] WLA[41] WLA[40] S55NLLGDPH_X512Y8D16_BW_EDGECELL8B
XI9 NET05 NET35 NET65 NET95 VDD VSS WLA[55] WLA[54] WLA[53] WLA[52]
+WLA[51] WLA[50] WLA[49] WLA[48] S55NLLGDPH_X512Y8D16_BW_EDGECELL8B
XI10 NET06 NET35 NET66 NET95 VDD VSS WLA[63] WLA[62] WLA[61] WLA[60]
+WLA[59] WLA[58] WLA[57] WLA[56] S55NLLGDPH_X512Y8D16_BW_EDGECELL8B
XI11 NET06 NET66 VDD VSS S55NLLGDPH_X512Y8D16_BW_BLSTRAP_B
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    S55NLLGDPH_X512Y8D16_BW_EDGECELL64A_RIGHT
* View Name:    schematic
************************************************************************

.SUBCKT S55NLLGDPH_X512Y8D16_BW_EDGECELL64A_RIGHT VDD VSS WLA[63] WLA[62] WLA[61] WLA[60] WLA[59] WLA[58] WLA[57] WLA[56]
+WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48] WLA[47] WLA[46]
+WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38] WLA[37] WLA[36]
+WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28] WLA[27] WLA[26]
+WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18] WLA[17] WLA[16]
+WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8] WLA[7] WLA[6]
+WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0]
XI0 NET01 NET61 VDD VSS S55NLLGDPH_X512Y8D16_BW_BLSTRAP
XI1 NET01 NET31 NET61 NET91 VDD VSS WLA[7] WLA[6] WLA[5] WLA[4]
+WLA[3] WLA[2] WLA[1] WLA[0] S55NLLGDPH_X512Y8D16_BW_EDGECELL8A
XI2 NET02 NET31 NET62 NET91 VDD VSS WLA[15] WLA[14] WLA[13] WLA[12]
+WLA[11] WLA[10] WLA[9] WLA[8] S55NLLGDPH_X512Y8D16_BW_EDGECELL8A
XI3 NET02 NET32 NET62 NET92 VDD VSS WLA[23] WLA[22] WLA[21] WLA[20]
+WLA[19] WLA[18] WLA[17] WLA[16] S55NLLGDPH_X512Y8D16_BW_EDGECELL8A
XI4 NET03 NET32 NET63 NET92 VDD VSS WLA[31] WLA[30] WLA[29] WLA[28]
+WLA[27] WLA[26] WLA[25] WLA[24] S55NLLGDPH_X512Y8D16_BW_EDGECELL8A
XI5 NET03 NET33 NET63 NET93 VDD VSS WLA[39] WLA[38] WLA[37] WLA[36]
+WLA[35] WLA[34] WLA[33] WLA[32] S55NLLGDPH_X512Y8D16_BW_EDGECELL8A
XI6 NET04 NET33 NET64 NET93 VDD VSS WLA[47] WLA[46] WLA[45] WLA[44]
+WLA[43] WLA[42] WLA[41] WLA[40] S55NLLGDPH_X512Y8D16_BW_EDGECELL8A
XI7 NET04 NET34 NET64 NET94 VDD VSS WLA[55] WLA[54] WLA[53] WLA[52]
+WLA[51] WLA[50] WLA[49] WLA[48] S55NLLGDPH_X512Y8D16_BW_EDGECELL8A
XI8 NET05 NET34 NET65 NET94 VDD VSS WLA[63] WLA[62] WLA[61] WLA[60]
+WLA[59] WLA[58] WLA[57] WLA[56] S55NLLGDPH_X512Y8D16_BW_EDGECELL8A
XI9 NET05 NET65 VDD VSS S55NLLGDPH_X512Y8D16_BW_BLSTRAP
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    S55NLLGDPH_X512Y8D16_BW_EDGECELL64B_RIGHT
* View Name:    schematic
************************************************************************

.SUBCKT S55NLLGDPH_X512Y8D16_BW_EDGECELL64B_RIGHT VDD VSS WLA[63] WLA[62] WLA[61] WLA[60] WLA[59] WLA[58] WLA[57] WLA[56]
+WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48] WLA[47] WLA[46]
+WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38] WLA[37] WLA[36]
+WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28] WLA[27] WLA[26]
+WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18] WLA[17] WLA[16]
+WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8] WLA[7] WLA[6]
+WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0]
XI0 NET01 NET61 VDD VSS S55NLLGDPH_X512Y8D16_BW_BLSTRAP_B
XI1 NET01 NET31 NET61 NET91 VDD VSS WLA[7] WLA[6] WLA[5] WLA[4]
+WLA[3] WLA[2] WLA[1] WLA[0] S55NLLGDPH_X512Y8D16_BW_EDGECELL8B
XI2 NET02 NET31 NET62 NET91 VDD VSS WLA[15] WLA[14] WLA[13] WLA[12]
+WLA[11] WLA[10] WLA[9] WLA[8] S55NLLGDPH_X512Y8D16_BW_EDGECELL8B
XI3 NET02 NET32 NET62 NET92 VDD VSS WLA[23] WLA[22] WLA[21] WLA[20]
+WLA[19] WLA[18] WLA[17] WLA[16] S55NLLGDPH_X512Y8D16_BW_EDGECELL8B
XI4 NET03 NET32 NET63 NET92 VDD VSS WLA[31] WLA[30] WLA[29] WLA[28]
+WLA[27] WLA[26] WLA[25] WLA[24] S55NLLGDPH_X512Y8D16_BW_EDGECELL8B
XI5 NET03 NET33 NET63 NET93 VDD VSS WLA[39] WLA[38] WLA[37] WLA[36]
+WLA[35] WLA[34] WLA[33] WLA[32] S55NLLGDPH_X512Y8D16_BW_EDGECELL8B
XI6 NET04 NET33 NET64 NET93 VDD VSS WLA[47] WLA[46] WLA[45] WLA[44]
+WLA[43] WLA[42] WLA[41] WLA[40] S55NLLGDPH_X512Y8D16_BW_EDGECELL8B
XI7 NET04 NET34 NET64 NET94 VDD VSS WLA[55] WLA[54] WLA[53] WLA[52]
+WLA[51] WLA[50] WLA[49] WLA[48] S55NLLGDPH_X512Y8D16_BW_EDGECELL8B
XI8 NET05 NET34 NET65 NET94 VDD VSS WLA[63] WLA[62] WLA[61] WLA[60]
+WLA[59] WLA[58] WLA[57] WLA[56] S55NLLGDPH_X512Y8D16_BW_EDGECELL8B
XI9 NET05 NET65 VDD VSS S55NLLGDPH_X512Y8D16_BW_BLSTRAP_B
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    S55NLLGDPH_X512Y8D16_BW_EDGECELL68A_TOP_RIGHT
* View Name:    schematic
************************************************************************

.SUBCKT S55NLLGDPH_X512Y8D16_BW_EDGECELL68A_TOP_RIGHT STWLA VDD VSS WLA[63] WLA[62] WLA[61] WLA[60] WLA[59] WLA[58] WLA[57]
+WLA[56] WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48] WLA[47]
+WLA[46] WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38] WLA[37]
+WLA[36] WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28] WLA[27]
+WLA[26] WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18] WLA[17]
+WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8] WLA[7]
+WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0]
XI0 NET01 NET61 VDD VSS S55NLLGDPH_X512Y8D16_BW_BLSTRAP
XI1 NET01 NET31 NET61 NET91 VDD VSS WLA[7] WLA[6] WLA[5] WLA[4]
+WLA[3] WLA[2] WLA[1] WLA[0] S55NLLGDPH_X512Y8D16_BW_EDGECELL8A
XI2 NET02 NET31 NET62 NET91 VDD VSS WLA[15] WLA[14] WLA[13] WLA[12]
+WLA[11] WLA[10] WLA[9] WLA[8] S55NLLGDPH_X512Y8D16_BW_EDGECELL8A
XI3 NET02 NET32 NET62 NET92 VDD VSS WLA[23] WLA[22] WLA[21] WLA[20]
+WLA[19] WLA[18] WLA[17] WLA[16] S55NLLGDPH_X512Y8D16_BW_EDGECELL8A
XI4 NET03 NET32 NET63 NET92 VDD VSS WLA[31] WLA[30] WLA[29] WLA[28]
+WLA[27] WLA[26] WLA[25] WLA[24] S55NLLGDPH_X512Y8D16_BW_EDGECELL8A
XI5 NET03 NET33 NET63 NET93 VDD VSS WLA[39] WLA[38] WLA[37] WLA[36]
+WLA[35] WLA[34] WLA[33] WLA[32] S55NLLGDPH_X512Y8D16_BW_EDGECELL8A
XI6 NET04 NET33 NET64 NET93 VDD VSS WLA[47] WLA[46] WLA[45] WLA[44]
+WLA[43] WLA[42] WLA[41] WLA[40] S55NLLGDPH_X512Y8D16_BW_EDGECELL8A
XI7 NET04 NET34 NET64 NET94 VDD VSS WLA[55] WLA[54] WLA[53] WLA[52]
+WLA[51] WLA[50] WLA[49] WLA[48] S55NLLGDPH_X512Y8D16_BW_EDGECELL8A
XI8 NET05 NET34 NET65 NET94 VDD VSS WLA[63] WLA[62] WLA[61] WLA[60]
+WLA[59] WLA[58] WLA[57] WLA[56] S55NLLGDPH_X512Y8D16_BW_EDGECELL8A
XI9 NET05 NET35 NET65 NET95 VDD VSS STWLA VSS VSS VSS S55NLLGDPH_X512Y8D16_BW_EDGECELL4A
XI10 NET35 NET95 VDD VSS S55NLLGDPH_X512Y8D16_BW_BLSTRAP
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    S55NLLGDPH_X512Y8D16_BW_BITCELL_ST64B_TW_RIGHT
* View Name:    schematic
************************************************************************

.SUBCKT S55NLLGDPH_X512Y8D16_BW_BITCELL_ST64B_TW_RIGHT DUM_BL VDD VSS WLA[63] WLA[62] WLA[61] WLA[60] WLA[59] WLA[58] WLA[57]
+WLA[56] WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48] WLA[47]
+WLA[46] WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38] WLA[37]
+WLA[36] WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28] WLA[27]
+WLA[26] WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18] WLA[17]
+WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8] WLA[7]
+WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0]
XI0 NET01 NET61 VDD VSS S55NLLGDPH_X512Y8D16_BW_BLSTRAP_B
XI1 NET01 NET31 NET61 NET91 DUM_BL VDD VSS WLA[7] WLA[6] WLA[5]
+WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST8B_TW
XI2 NET02 NET31 NET62 NET91 DUM_BL VDD VSS WLA[15] WLA[14] WLA[13]
+WLA[12] WLA[11] WLA[10] WLA[9] WLA[8] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST8B_TW
XI3 NET02 NET32 NET62 NET92 DUM_BL VDD VSS WLA[23] WLA[22] WLA[21]
+WLA[20] WLA[19] WLA[18] WLA[17] WLA[16] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST8B_TW
XI4 NET03 NET32 NET63 NET92 DUM_BL VDD VSS WLA[31] WLA[30] WLA[29]
+WLA[28] WLA[27] WLA[26] WLA[25] WLA[24] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST8B_TW
XI5 NET03 NET33 NET63 NET93 DUM_BL VDD VSS WLA[39] WLA[38] WLA[37]
+WLA[36] WLA[35] WLA[34] WLA[33] WLA[32] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST8B_TW
XI6 NET04 NET33 NET64 NET93 DUM_BL VDD VSS WLA[47] WLA[46] WLA[45]
+WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST8B_TW
XI7 NET04 NET34 NET64 NET94 DUM_BL VDD VSS WLA[55] WLA[54] WLA[53]
+WLA[52] WLA[51] WLA[50] WLA[49] WLA[48] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST8B_TW
XI8 NET05 NET34 NET65 NET94 DUM_BL VDD VSS WLA[63] WLA[62] WLA[61]
+WLA[60] WLA[59] WLA[58] WLA[57] WLA[56] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST8B_TW
XI9 NET05 NET65 VDD VSS S55NLLGDPH_X512Y8D16_BW_BLSTRAP_B
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    S55NLLGDPH_X512Y8D16_BW_BITCELL_ST64A_TW_RIGHT
* View Name:    schematic
************************************************************************

.SUBCKT S55NLLGDPH_X512Y8D16_BW_BITCELL_ST64A_TW_RIGHT DUM_BL VDD VSS WLA[63] WLA[62] WLA[61] WLA[60] WLA[59] WLA[58] WLA[57]
+WLA[56] WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48] WLA[47]
+WLA[46] WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38] WLA[37]
+WLA[36] WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28] WLA[27]
+WLA[26] WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18] WLA[17]
+WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8] WLA[7]
+WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0]
XI0 NET01 DUM_BL VDD VSS S55NLLGDPH_X512Y8D16_BW_BLSTRAP
XI1 NET01 NET31 DUM_BL VDD VSS WLA[7] WLA[6] WLA[5] WLA[4] WLA[3]
+WLA[2] WLA[1] WLA[0] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST8A_TW
XI2 NET02 NET31 DUM_BL VDD VSS WLA[15] WLA[14] WLA[13] WLA[12] WLA[11]
+WLA[10] WLA[9] WLA[8] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST8A_TW
XI3 NET02 NET32 DUM_BL VDD VSS WLA[23] WLA[22] WLA[21] WLA[20] WLA[19]
+WLA[18] WLA[17] WLA[16] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST8A_TW
XI4 NET03 NET32 DUM_BL VDD VSS WLA[31] WLA[30] WLA[29] WLA[28] WLA[27]
+WLA[26] WLA[25] WLA[24] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST8A_TW
XI5 NET03 NET33 DUM_BL VDD VSS WLA[39] WLA[38] WLA[37] WLA[36] WLA[35]
+WLA[34] WLA[33] WLA[32] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST8A_TW
XI6 NET04 NET33 DUM_BL VDD VSS WLA[47] WLA[46] WLA[45] WLA[44] WLA[43]
+WLA[42] WLA[41] WLA[40] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST8A_TW
XI7 NET04 NET34 DUM_BL VDD VSS WLA[55] WLA[54] WLA[53] WLA[52] WLA[51]
+WLA[50] WLA[49] WLA[48] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST8A_TW
XI8 NET05 NET34 DUM_BL VDD VSS WLA[63] WLA[62] WLA[61] WLA[60] WLA[59]
+WLA[58] WLA[57] WLA[56] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST8A_TW
XI9 NET05 DUM_BL VDD VSS S55NLLGDPH_X512Y8D16_BW_BLSTRAP
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    S55NLLGDPH_X512Y8D16_BW_BITCELL_ST68A_TOP_TW_RIGHT
* View Name:    schematic
************************************************************************

.SUBCKT S55NLLGDPH_X512Y8D16_BW_BITCELL_ST68A_TOP_TW_RIGHT DUM_BL STWLA VDD VSS WLA[63] WLA[62] WLA[61] WLA[60] WLA[59] WLA[58]
+WLA[57] WLA[56] WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48]
+WLA[47] WLA[46] WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38]
+WLA[37] WLA[36] WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28]
+WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18]
+WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8]
+WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0]
XI0 NET01 DUM_BL VDD VSS S55NLLGDPH_X512Y8D16_BW_BLSTRAP
XI1 NET01 NET31 DUM_BL VDD VSS WLA[7] WLA[6] WLA[5] WLA[4] WLA[3]
+WLA[2] WLA[1] WLA[0] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST8A_TW
XI2 NET02 NET31 DUM_BL VDD VSS WLA[15] WLA[14] WLA[13] WLA[12] WLA[11]
+WLA[10] WLA[9] WLA[8] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST8A_TW
XI3 NET02 NET32 DUM_BL VDD VSS WLA[23] WLA[22] WLA[21] WLA[20] WLA[19]
+WLA[18] WLA[17] WLA[16] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST8A_TW
XI4 NET03 NET32 DUM_BL VDD VSS WLA[31] WLA[30] WLA[29] WLA[28] WLA[27]
+WLA[26] WLA[25] WLA[24] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST8A_TW
XI5 NET03 NET33 DUM_BL VDD VSS WLA[39] WLA[38] WLA[37] WLA[36] WLA[35]
+WLA[34] WLA[33] WLA[32] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST8A_TW
XI6 NET04 NET33 DUM_BL VDD VSS WLA[47] WLA[46] WLA[45] WLA[44] WLA[43]
+WLA[42] WLA[41] WLA[40] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST8A_TW
XI7 NET04 NET34 DUM_BL VDD VSS WLA[55] WLA[54] WLA[53] WLA[52] WLA[51]
+WLA[50] WLA[49] WLA[48] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST8A_TW
XI8 NET05 NET34 DUM_BL VDD VSS WLA[63] WLA[62] WLA[61] WLA[60] WLA[59]
+WLA[58] WLA[57] WLA[56] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST8A_TW
XI9 NET05 NET4 DUM_BL NET5 VDD VSS STWLA VSS VSS VSS S55NLLGDPH_X512Y8D16_BW_BITCELL_ST4A_TW
XI10 NET4 NET5 VDD VSS S55NLLGDPH_X512Y8D16_BW_BLSTRAP
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    S55NLLGDPH_X512Y8D16_BW_Y512X8CELLX8_BW_RIGHT
* View Name:    schematic
************************************************************************

.SUBCKT S55NLLGDPH_X512Y8D16_BW_Y512X8CELLX8_BW_RIGHT BWENA[7] BWENA[6] BWENA[5] BWENA[4] BWENA[3] BWENA[2] BWENA[1] BWENA[0] BWENB[7] BWENB[6]
+BWENB[5] BWENB[4] BWENB[3] BWENB[2] BWENB[1] BWENB[0] CLKA CLKB CLKXA CLKXB
+DATAA[7] DATAA[6] DATAA[5] DATAA[4] DATAA[3] DATAA[2] DATAA[1] DATAA[0] DATAB[7] DATAB[6]
+DATAB[5] DATAB[4] DATAB[3] DATAB[2] DATAB[1] DATAB[0] DBL DOUTA[7] DOUTA[6] DOUTA[5]
+DOUTA[4] DOUTA[3] DOUTA[2] DOUTA[1] DOUTA[0] DOUTB[7] DOUTB[6] DOUTB[5] DOUTB[4] DOUTB[3]
+DOUTB[2] DOUTB[1] DOUTB[0] RWLA[0] RWLA[1] RWLB[0] RWLB[1] SACK1A SACK1B SACK4A
+SACK4B STWLA STWLB VDD VSS WEA WEB WLA[511] WLA[510] WLA[509]
+WLA[508] WLA[507] WLA[506] WLA[505] WLA[504] WLA[503] WLA[502] WLA[501] WLA[500] WLA[499]
+WLA[498] WLA[497] WLA[496] WLA[495] WLA[494] WLA[493] WLA[492] WLA[491] WLA[490] WLA[489]
+WLA[488] WLA[487] WLA[486] WLA[485] WLA[484] WLA[483] WLA[482] WLA[481] WLA[480] WLA[479]
+WLA[478] WLA[477] WLA[476] WLA[475] WLA[474] WLA[473] WLA[472] WLA[471] WLA[470] WLA[469]
+WLA[468] WLA[467] WLA[466] WLA[465] WLA[464] WLA[463] WLA[462] WLA[461] WLA[460] WLA[459]
+WLA[458] WLA[457] WLA[456] WLA[455] WLA[454] WLA[453] WLA[452] WLA[451] WLA[450] WLA[449]
+WLA[448] WLA[447] WLA[446] WLA[445] WLA[444] WLA[443] WLA[442] WLA[441] WLA[440] WLA[439]
+WLA[438] WLA[437] WLA[436] WLA[435] WLA[434] WLA[433] WLA[432] WLA[431] WLA[430] WLA[429]
+WLA[428] WLA[427] WLA[426] WLA[425] WLA[424] WLA[423] WLA[422] WLA[421] WLA[420] WLA[419]
+WLA[418] WLA[417] WLA[416] WLA[415] WLA[414] WLA[413] WLA[412] WLA[411] WLA[410] WLA[409]
+WLA[408] WLA[407] WLA[406] WLA[405] WLA[404] WLA[403] WLA[402] WLA[401] WLA[400] WLA[399]
+WLA[398] WLA[397] WLA[396] WLA[395] WLA[394] WLA[393] WLA[392] WLA[391] WLA[390] WLA[389]
+WLA[388] WLA[387] WLA[386] WLA[385] WLA[384] WLA[383] WLA[382] WLA[381] WLA[380] WLA[379]
+WLA[378] WLA[377] WLA[376] WLA[375] WLA[374] WLA[373] WLA[372] WLA[371] WLA[370] WLA[369]
+WLA[368] WLA[367] WLA[366] WLA[365] WLA[364] WLA[363] WLA[362] WLA[361] WLA[360] WLA[359]
+WLA[358] WLA[357] WLA[356] WLA[355] WLA[354] WLA[353] WLA[352] WLA[351] WLA[350] WLA[349]
+WLA[348] WLA[347] WLA[346] WLA[345] WLA[344] WLA[343] WLA[342] WLA[341] WLA[340] WLA[339]
+WLA[338] WLA[337] WLA[336] WLA[335] WLA[334] WLA[333] WLA[332] WLA[331] WLA[330] WLA[329]
+WLA[328] WLA[327] WLA[326] WLA[325] WLA[324] WLA[323] WLA[322] WLA[321] WLA[320] WLA[319]
+WLA[318] WLA[317] WLA[316] WLA[315] WLA[314] WLA[313] WLA[312] WLA[311] WLA[310] WLA[309]
+WLA[308] WLA[307] WLA[306] WLA[305] WLA[304] WLA[303] WLA[302] WLA[301] WLA[300] WLA[299]
+WLA[298] WLA[297] WLA[296] WLA[295] WLA[294] WLA[293] WLA[292] WLA[291] WLA[290] WLA[289]
+WLA[288] WLA[287] WLA[286] WLA[285] WLA[284] WLA[283] WLA[282] WLA[281] WLA[280] WLA[279]
+WLA[278] WLA[277] WLA[276] WLA[275] WLA[274] WLA[273] WLA[272] WLA[271] WLA[270] WLA[269]
+WLA[268] WLA[267] WLA[266] WLA[265] WLA[264] WLA[263] WLA[262] WLA[261] WLA[260] WLA[259]
+WLA[258] WLA[257] WLA[256] WLA[255] WLA[254] WLA[253] WLA[252] WLA[251] WLA[250] WLA[249]
+WLA[248] WLA[247] WLA[246] WLA[245] WLA[244] WLA[243] WLA[242] WLA[241] WLA[240] WLA[239]
+WLA[238] WLA[237] WLA[236] WLA[235] WLA[234] WLA[233] WLA[232] WLA[231] WLA[230] WLA[229]
+WLA[228] WLA[227] WLA[226] WLA[225] WLA[224] WLA[223] WLA[222] WLA[221] WLA[220] WLA[219]
+WLA[218] WLA[217] WLA[216] WLA[215] WLA[214] WLA[213] WLA[212] WLA[211] WLA[210] WLA[209]
+WLA[208] WLA[207] WLA[206] WLA[205] WLA[204] WLA[203] WLA[202] WLA[201] WLA[200] WLA[199]
+WLA[198] WLA[197] WLA[196] WLA[195] WLA[194] WLA[193] WLA[192] WLA[191] WLA[190] WLA[189]
+WLA[188] WLA[187] WLA[186] WLA[185] WLA[184] WLA[183] WLA[182] WLA[181] WLA[180] WLA[179]
+WLA[178] WLA[177] WLA[176] WLA[175] WLA[174] WLA[173] WLA[172] WLA[171] WLA[170] WLA[169]
+WLA[168] WLA[167] WLA[166] WLA[165] WLA[164] WLA[163] WLA[162] WLA[161] WLA[160] WLA[159]
+WLA[158] WLA[157] WLA[156] WLA[155] WLA[154] WLA[153] WLA[152] WLA[151] WLA[150] WLA[149]
+WLA[148] WLA[147] WLA[146] WLA[145] WLA[144] WLA[143] WLA[142] WLA[141] WLA[140] WLA[139]
+WLA[138] WLA[137] WLA[136] WLA[135] WLA[134] WLA[133] WLA[132] WLA[131] WLA[130] WLA[129]
+WLA[128] WLA[127] WLA[126] WLA[125] WLA[124] WLA[123] WLA[122] WLA[121] WLA[120] WLA[119]
+WLA[118] WLA[117] WLA[116] WLA[115] WLA[114] WLA[113] WLA[112] WLA[111] WLA[110] WLA[109]
+WLA[108] WLA[107] WLA[106] WLA[105] WLA[104] WLA[103] WLA[102] WLA[101] WLA[100] WLA[99]
+WLA[98] WLA[97] WLA[96] WLA[95] WLA[94] WLA[93] WLA[92] WLA[91] WLA[90] WLA[89]
+WLA[88] WLA[87] WLA[86] WLA[85] WLA[84] WLA[83] WLA[82] WLA[81] WLA[80] WLA[79]
+WLA[78] WLA[77] WLA[76] WLA[75] WLA[74] WLA[73] WLA[72] WLA[71] WLA[70] WLA[69]
+WLA[68] WLA[67] WLA[66] WLA[65] WLA[64] WLA[63] WLA[62] WLA[61] WLA[60] WLA[59]
+WLA[58] WLA[57] WLA[56] WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50] WLA[49]
+WLA[48] WLA[47] WLA[46] WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39]
+WLA[38] WLA[37] WLA[36] WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29]
+WLA[28] WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19]
+WLA[18] WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9]
+WLA[8] WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] WLB[511]
+WLB[510] WLB[509] WLB[508] WLB[507] WLB[506] WLB[505] WLB[504] WLB[503] WLB[502] WLB[501]
+WLB[500] WLB[499] WLB[498] WLB[497] WLB[496] WLB[495] WLB[494] WLB[493] WLB[492] WLB[491]
+WLB[490] WLB[489] WLB[488] WLB[487] WLB[486] WLB[485] WLB[484] WLB[483] WLB[482] WLB[481]
+WLB[480] WLB[479] WLB[478] WLB[477] WLB[476] WLB[475] WLB[474] WLB[473] WLB[472] WLB[471]
+WLB[470] WLB[469] WLB[468] WLB[467] WLB[466] WLB[465] WLB[464] WLB[463] WLB[462] WLB[461]
+WLB[460] WLB[459] WLB[458] WLB[457] WLB[456] WLB[455] WLB[454] WLB[453] WLB[452] WLB[451]
+WLB[450] WLB[449] WLB[448] WLB[447] WLB[446] WLB[445] WLB[444] WLB[443] WLB[442] WLB[441]
+WLB[440] WLB[439] WLB[438] WLB[437] WLB[436] WLB[435] WLB[434] WLB[433] WLB[432] WLB[431]
+WLB[430] WLB[429] WLB[428] WLB[427] WLB[426] WLB[425] WLB[424] WLB[423] WLB[422] WLB[421]
+WLB[420] WLB[419] WLB[418] WLB[417] WLB[416] WLB[415] WLB[414] WLB[413] WLB[412] WLB[411]
+WLB[410] WLB[409] WLB[408] WLB[407] WLB[406] WLB[405] WLB[404] WLB[403] WLB[402] WLB[401]
+WLB[400] WLB[399] WLB[398] WLB[397] WLB[396] WLB[395] WLB[394] WLB[393] WLB[392] WLB[391]
+WLB[390] WLB[389] WLB[388] WLB[387] WLB[386] WLB[385] WLB[384] WLB[383] WLB[382] WLB[381]
+WLB[380] WLB[379] WLB[378] WLB[377] WLB[376] WLB[375] WLB[374] WLB[373] WLB[372] WLB[371]
+WLB[370] WLB[369] WLB[368] WLB[367] WLB[366] WLB[365] WLB[364] WLB[363] WLB[362] WLB[361]
+WLB[360] WLB[359] WLB[358] WLB[357] WLB[356] WLB[355] WLB[354] WLB[353] WLB[352] WLB[351]
+WLB[350] WLB[349] WLB[348] WLB[347] WLB[346] WLB[345] WLB[344] WLB[343] WLB[342] WLB[341]
+WLB[340] WLB[339] WLB[338] WLB[337] WLB[336] WLB[335] WLB[334] WLB[333] WLB[332] WLB[331]
+WLB[330] WLB[329] WLB[328] WLB[327] WLB[326] WLB[325] WLB[324] WLB[323] WLB[322] WLB[321]
+WLB[320] WLB[319] WLB[318] WLB[317] WLB[316] WLB[315] WLB[314] WLB[313] WLB[312] WLB[311]
+WLB[310] WLB[309] WLB[308] WLB[307] WLB[306] WLB[305] WLB[304] WLB[303] WLB[302] WLB[301]
+WLB[300] WLB[299] WLB[298] WLB[297] WLB[296] WLB[295] WLB[294] WLB[293] WLB[292] WLB[291]
+WLB[290] WLB[289] WLB[288] WLB[287] WLB[286] WLB[285] WLB[284] WLB[283] WLB[282] WLB[281]
+WLB[280] WLB[279] WLB[278] WLB[277] WLB[276] WLB[275] WLB[274] WLB[273] WLB[272] WLB[271]
+WLB[270] WLB[269] WLB[268] WLB[267] WLB[266] WLB[265] WLB[264] WLB[263] WLB[262] WLB[261]
+WLB[260] WLB[259] WLB[258] WLB[257] WLB[256] WLB[255] WLB[254] WLB[253] WLB[252] WLB[251]
+WLB[250] WLB[249] WLB[248] WLB[247] WLB[246] WLB[245] WLB[244] WLB[243] WLB[242] WLB[241]
+WLB[240] WLB[239] WLB[238] WLB[237] WLB[236] WLB[235] WLB[234] WLB[233] WLB[232] WLB[231]
+WLB[230] WLB[229] WLB[228] WLB[227] WLB[226] WLB[225] WLB[224] WLB[223] WLB[222] WLB[221]
+WLB[220] WLB[219] WLB[218] WLB[217] WLB[216] WLB[215] WLB[214] WLB[213] WLB[212] WLB[211]
+WLB[210] WLB[209] WLB[208] WLB[207] WLB[206] WLB[205] WLB[204] WLB[203] WLB[202] WLB[201]
+WLB[200] WLB[199] WLB[198] WLB[197] WLB[196] WLB[195] WLB[194] WLB[193] WLB[192] WLB[191]
+WLB[190] WLB[189] WLB[188] WLB[187] WLB[186] WLB[185] WLB[184] WLB[183] WLB[182] WLB[181]
+WLB[180] WLB[179] WLB[178] WLB[177] WLB[176] WLB[175] WLB[174] WLB[173] WLB[172] WLB[171]
+WLB[170] WLB[169] WLB[168] WLB[167] WLB[166] WLB[165] WLB[164] WLB[163] WLB[162] WLB[161]
+WLB[160] WLB[159] WLB[158] WLB[157] WLB[156] WLB[155] WLB[154] WLB[153] WLB[152] WLB[151]
+WLB[150] WLB[149] WLB[148] WLB[147] WLB[146] WLB[145] WLB[144] WLB[143] WLB[142] WLB[141]
+WLB[140] WLB[139] WLB[138] WLB[137] WLB[136] WLB[135] WLB[134] WLB[133] WLB[132] WLB[131]
+WLB[130] WLB[129] WLB[128] WLB[127] WLB[126] WLB[125] WLB[124] WLB[123] WLB[122] WLB[121]
+WLB[120] WLB[119] WLB[118] WLB[117] WLB[116] WLB[115] WLB[114] WLB[113] WLB[112] WLB[111]
+WLB[110] WLB[109] WLB[108] WLB[107] WLB[106] WLB[105] WLB[104] WLB[103] WLB[102] WLB[101]
+WLB[100] WLB[99] WLB[98] WLB[97] WLB[96] WLB[95] WLB[94] WLB[93] WLB[92] WLB[91]
+WLB[90] WLB[89] WLB[88] WLB[87] WLB[86] WLB[85] WLB[84] WLB[83] WLB[82] WLB[81]
+WLB[80] WLB[79] WLB[78] WLB[77] WLB[76] WLB[75] WLB[74] WLB[73] WLB[72] WLB[71]
+WLB[70] WLB[69] WLB[68] WLB[67] WLB[66] WLB[65] WLB[64] WLB[63] WLB[62] WLB[61]
+WLB[60] WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54] WLB[53] WLB[52] WLB[51]
+WLB[50] WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44] WLB[43] WLB[42] WLB[41]
+WLB[40] WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34] WLB[33] WLB[32] WLB[31]
+WLB[30] WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24] WLB[23] WLB[22] WLB[21]
+WLB[20] WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14] WLB[13] WLB[12] WLB[11]
+WLB[10] WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4] WLB[3] WLB[2] WLB[1]
+WLB[0] YXA[7] YXA[6] YXA[5] YXA[4] YXA[3] YXA[2] YXA[1] YXA[0] YXB[7]
+YXB[6] YXB[5] YXB[4] YXB[3] YXB[2] YXB[1] YXB[0]
XI0 RWLA[0] RWLA[1] VDD VSS WLA[63] WLA[62] WLA[61] WLA[60] WLA[59] WLA[58]
+WLA[57] WLA[56] WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48]
+WLA[47] WLA[46] WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38]
+WLA[37] WLA[36] WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28]
+WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18]
+WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8]
+WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] S55NLLGDPH_X512Y8D16_BW_EDGECELL66B_RED_RIGHT
XI1 VDD VSS WLA[127] WLA[126] WLA[125] WLA[124] WLA[123] WLA[122] WLA[121] WLA[120]
+WLA[119] WLA[118] WLA[117] WLA[116] WLA[115] WLA[114] WLA[113] WLA[112] WLA[111] WLA[110]
+WLA[109] WLA[108] WLA[107] WLA[106] WLA[105] WLA[104] WLA[103] WLA[102] WLA[101] WLA[100]
+WLA[99] WLA[98] WLA[97] WLA[96] WLA[95] WLA[94] WLA[93] WLA[92] WLA[91] WLA[90]
+WLA[89] WLA[88] WLA[87] WLA[86] WLA[85] WLA[84] WLA[83] WLA[82] WLA[81] WLA[80]
+WLA[79] WLA[78] WLA[77] WLA[76] WLA[75] WLA[74] WLA[73] WLA[72] WLA[71] WLA[70]
+WLA[69] WLA[68] WLA[67] WLA[66] WLA[65] WLA[64] S55NLLGDPH_X512Y8D16_BW_EDGECELL64A_RIGHT
XI2 VDD VSS WLA[191] WLA[190] WLA[189] WLA[188] WLA[187] WLA[186] WLA[185] WLA[184]
+WLA[183] WLA[182] WLA[181] WLA[180] WLA[179] WLA[178] WLA[177] WLA[176] WLA[175] WLA[174]
+WLA[173] WLA[172] WLA[171] WLA[170] WLA[169] WLA[168] WLA[167] WLA[166] WLA[165] WLA[164]
+WLA[163] WLA[162] WLA[161] WLA[160] WLA[159] WLA[158] WLA[157] WLA[156] WLA[155] WLA[154]
+WLA[153] WLA[152] WLA[151] WLA[150] WLA[149] WLA[148] WLA[147] WLA[146] WLA[145] WLA[144]
+WLA[143] WLA[142] WLA[141] WLA[140] WLA[139] WLA[138] WLA[137] WLA[136] WLA[135] WLA[134]
+WLA[133] WLA[132] WLA[131] WLA[130] WLA[129] WLA[128] S55NLLGDPH_X512Y8D16_BW_EDGECELL64B_RIGHT
XI3 VDD VSS WLA[255] WLA[254] WLA[253] WLA[252] WLA[251] WLA[250] WLA[249] WLA[248]
+WLA[247] WLA[246] WLA[245] WLA[244] WLA[243] WLA[242] WLA[241] WLA[240] WLA[239] WLA[238]
+WLA[237] WLA[236] WLA[235] WLA[234] WLA[233] WLA[232] WLA[231] WLA[230] WLA[229] WLA[228]
+WLA[227] WLA[226] WLA[225] WLA[224] WLA[223] WLA[222] WLA[221] WLA[220] WLA[219] WLA[218]
+WLA[217] WLA[216] WLA[215] WLA[214] WLA[213] WLA[212] WLA[211] WLA[210] WLA[209] WLA[208]
+WLA[207] WLA[206] WLA[205] WLA[204] WLA[203] WLA[202] WLA[201] WLA[200] WLA[199] WLA[198]
+WLA[197] WLA[196] WLA[195] WLA[194] WLA[193] WLA[192] S55NLLGDPH_X512Y8D16_BW_EDGECELL64A_RIGHT
XI4 VDD VSS WLA[319] WLA[318] WLA[317] WLA[316] WLA[315] WLA[314] WLA[313] WLA[312]
+WLA[311] WLA[310] WLA[309] WLA[308] WLA[307] WLA[306] WLA[305] WLA[304] WLA[303] WLA[302]
+WLA[301] WLA[300] WLA[299] WLA[298] WLA[297] WLA[296] WLA[295] WLA[294] WLA[293] WLA[292]
+WLA[291] WLA[290] WLA[289] WLA[288] WLA[287] WLA[286] WLA[285] WLA[284] WLA[283] WLA[282]
+WLA[281] WLA[280] WLA[279] WLA[278] WLA[277] WLA[276] WLA[275] WLA[274] WLA[273] WLA[272]
+WLA[271] WLA[270] WLA[269] WLA[268] WLA[267] WLA[266] WLA[265] WLA[264] WLA[263] WLA[262]
+WLA[261] WLA[260] WLA[259] WLA[258] WLA[257] WLA[256] S55NLLGDPH_X512Y8D16_BW_EDGECELL64B_RIGHT
XI5 VDD VSS WLA[383] WLA[382] WLA[381] WLA[380] WLA[379] WLA[378] WLA[377] WLA[376]
+WLA[375] WLA[374] WLA[373] WLA[372] WLA[371] WLA[370] WLA[369] WLA[368] WLA[367] WLA[366]
+WLA[365] WLA[364] WLA[363] WLA[362] WLA[361] WLA[360] WLA[359] WLA[358] WLA[357] WLA[356]
+WLA[355] WLA[354] WLA[353] WLA[352] WLA[351] WLA[350] WLA[349] WLA[348] WLA[347] WLA[346]
+WLA[345] WLA[344] WLA[343] WLA[342] WLA[341] WLA[340] WLA[339] WLA[338] WLA[337] WLA[336]
+WLA[335] WLA[334] WLA[333] WLA[332] WLA[331] WLA[330] WLA[329] WLA[328] WLA[327] WLA[326]
+WLA[325] WLA[324] WLA[323] WLA[322] WLA[321] WLA[320] S55NLLGDPH_X512Y8D16_BW_EDGECELL64A_RIGHT
XI6 VDD VSS WLA[447] WLA[446] WLA[445] WLA[444] WLA[443] WLA[442] WLA[441] WLA[440]
+WLA[439] WLA[438] WLA[437] WLA[436] WLA[435] WLA[434] WLA[433] WLA[432] WLA[431] WLA[430]
+WLA[429] WLA[428] WLA[427] WLA[426] WLA[425] WLA[424] WLA[423] WLA[422] WLA[421] WLA[420]
+WLA[419] WLA[418] WLA[417] WLA[416] WLA[415] WLA[414] WLA[413] WLA[412] WLA[411] WLA[410]
+WLA[409] WLA[408] WLA[407] WLA[406] WLA[405] WLA[404] WLA[403] WLA[402] WLA[401] WLA[400]
+WLA[399] WLA[398] WLA[397] WLA[396] WLA[395] WLA[394] WLA[393] WLA[392] WLA[391] WLA[390]
+WLA[389] WLA[388] WLA[387] WLA[386] WLA[385] WLA[384] S55NLLGDPH_X512Y8D16_BW_EDGECELL64B_RIGHT
XI7 STWLA VDD VSS WLA[511] WLA[510] WLA[509] WLA[508] WLA[507] WLA[506] WLA[505]
+WLA[504] WLA[503] WLA[502] WLA[501] WLA[500] WLA[499] WLA[498] WLA[497] WLA[496] WLA[495]
+WLA[494] WLA[493] WLA[492] WLA[491] WLA[490] WLA[489] WLA[488] WLA[487] WLA[486] WLA[485]
+WLA[484] WLA[483] WLA[482] WLA[481] WLA[480] WLA[479] WLA[478] WLA[477] WLA[476] WLA[475]
+WLA[474] WLA[473] WLA[472] WLA[471] WLA[470] WLA[469] WLA[468] WLA[467] WLA[466] WLA[465]
+WLA[464] WLA[463] WLA[462] WLA[461] WLA[460] WLA[459] WLA[458] WLA[457] WLA[456] WLA[455]
+WLA[454] WLA[453] WLA[452] WLA[451] WLA[450] WLA[449] WLA[448] S55NLLGDPH_X512Y8D16_BW_EDGECELL68A_TOP_RIGHT
XI8 DBL RWLA[0] RWLA[1] VDD VSS WLA[63] WLA[62] WLA[61] WLA[60] WLA[59]
+WLA[58] WLA[57] WLA[56] WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50] WLA[49]
+WLA[48] WLA[47] WLA[46] WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39]
+WLA[38] WLA[37] WLA[36] WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29]
+WLA[28] WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19]
+WLA[18] WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9]
+WLA[8] WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST66B
XI9 DBL VDD VSS WLA[127] WLA[126] WLA[125] WLA[124] WLA[123] WLA[122] WLA[121]
+WLA[120] WLA[119] WLA[118] WLA[117] WLA[116] WLA[115] WLA[114] WLA[113] WLA[112] WLA[111]
+WLA[110] WLA[109] WLA[108] WLA[107] WLA[106] WLA[105] WLA[104] WLA[103] WLA[102] WLA[101]
+WLA[100] WLA[99] WLA[98] WLA[97] WLA[96] WLA[95] WLA[94] WLA[93] WLA[92] WLA[91]
+WLA[90] WLA[89] WLA[88] WLA[87] WLA[86] WLA[85] WLA[84] WLA[83] WLA[82] WLA[81]
+WLA[80] WLA[79] WLA[78] WLA[77] WLA[76] WLA[75] WLA[74] WLA[73] WLA[72] WLA[71]
+WLA[70] WLA[69] WLA[68] WLA[67] WLA[66] WLA[65] WLA[64] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST64A
XI10 DBL VDD VSS WLA[191] WLA[190] WLA[189] WLA[188] WLA[187] WLA[186] WLA[185]
+WLA[184] WLA[183] WLA[182] WLA[181] WLA[180] WLA[179] WLA[178] WLA[177] WLA[176] WLA[175]
+WLA[174] WLA[173] WLA[172] WLA[171] WLA[170] WLA[169] WLA[168] WLA[167] WLA[166] WLA[165]
+WLA[164] WLA[163] WLA[162] WLA[161] WLA[160] WLA[159] WLA[158] WLA[157] WLA[156] WLA[155]
+WLA[154] WLA[153] WLA[152] WLA[151] WLA[150] WLA[149] WLA[148] WLA[147] WLA[146] WLA[145]
+WLA[144] WLA[143] WLA[142] WLA[141] WLA[140] WLA[139] WLA[138] WLA[137] WLA[136] WLA[135]
+WLA[134] WLA[133] WLA[132] WLA[131] WLA[130] WLA[129] WLA[128] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST64B
XI11 DBL VDD VSS WLA[255] WLA[254] WLA[253] WLA[252] WLA[251] WLA[250] WLA[249]
+WLA[248] WLA[247] WLA[246] WLA[245] WLA[244] WLA[243] WLA[242] WLA[241] WLA[240] WLA[239]
+WLA[238] WLA[237] WLA[236] WLA[235] WLA[234] WLA[233] WLA[232] WLA[231] WLA[230] WLA[229]
+WLA[228] WLA[227] WLA[226] WLA[225] WLA[224] WLA[223] WLA[222] WLA[221] WLA[220] WLA[219]
+WLA[218] WLA[217] WLA[216] WLA[215] WLA[214] WLA[213] WLA[212] WLA[211] WLA[210] WLA[209]
+WLA[208] WLA[207] WLA[206] WLA[205] WLA[204] WLA[203] WLA[202] WLA[201] WLA[200] WLA[199]
+WLA[198] WLA[197] WLA[196] WLA[195] WLA[194] WLA[193] WLA[192] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST64A
XI12 DBL VDD VSS WLA[319] WLA[318] WLA[317] WLA[316] WLA[315] WLA[314] WLA[313]
+WLA[312] WLA[311] WLA[310] WLA[309] WLA[308] WLA[307] WLA[306] WLA[305] WLA[304] WLA[303]
+WLA[302] WLA[301] WLA[300] WLA[299] WLA[298] WLA[297] WLA[296] WLA[295] WLA[294] WLA[293]
+WLA[292] WLA[291] WLA[290] WLA[289] WLA[288] WLA[287] WLA[286] WLA[285] WLA[284] WLA[283]
+WLA[282] WLA[281] WLA[280] WLA[279] WLA[278] WLA[277] WLA[276] WLA[275] WLA[274] WLA[273]
+WLA[272] WLA[271] WLA[270] WLA[269] WLA[268] WLA[267] WLA[266] WLA[265] WLA[264] WLA[263]
+WLA[262] WLA[261] WLA[260] WLA[259] WLA[258] WLA[257] WLA[256] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST64B_TW_RIGHT
XI13 DBL VDD VSS WLA[383] WLA[382] WLA[381] WLA[380] WLA[379] WLA[378] WLA[377]
+WLA[376] WLA[375] WLA[374] WLA[373] WLA[372] WLA[371] WLA[370] WLA[369] WLA[368] WLA[367]
+WLA[366] WLA[365] WLA[364] WLA[363] WLA[362] WLA[361] WLA[360] WLA[359] WLA[358] WLA[357]
+WLA[356] WLA[355] WLA[354] WLA[353] WLA[352] WLA[351] WLA[350] WLA[349] WLA[348] WLA[347]
+WLA[346] WLA[345] WLA[344] WLA[343] WLA[342] WLA[341] WLA[340] WLA[339] WLA[338] WLA[337]
+WLA[336] WLA[335] WLA[334] WLA[333] WLA[332] WLA[331] WLA[330] WLA[329] WLA[328] WLA[327]
+WLA[326] WLA[325] WLA[324] WLA[323] WLA[322] WLA[321] WLA[320] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST64A_TW_RIGHT
XI14 DBL VDD VSS WLA[447] WLA[446] WLA[445] WLA[444] WLA[443] WLA[442] WLA[441]
+WLA[440] WLA[439] WLA[438] WLA[437] WLA[436] WLA[435] WLA[434] WLA[433] WLA[432] WLA[431]
+WLA[430] WLA[429] WLA[428] WLA[427] WLA[426] WLA[425] WLA[424] WLA[423] WLA[422] WLA[421]
+WLA[420] WLA[419] WLA[418] WLA[417] WLA[416] WLA[415] WLA[414] WLA[413] WLA[412] WLA[411]
+WLA[410] WLA[409] WLA[408] WLA[407] WLA[406] WLA[405] WLA[404] WLA[403] WLA[402] WLA[401]
+WLA[400] WLA[399] WLA[398] WLA[397] WLA[396] WLA[395] WLA[394] WLA[393] WLA[392] WLA[391]
+WLA[390] WLA[389] WLA[388] WLA[387] WLA[386] WLA[385] WLA[384] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST64B_TW_RIGHT
XI15 DBL STWLA VDD VSS WLA[511] WLA[510] WLA[509] WLA[508] WLA[507] WLA[506]
+WLA[505] WLA[504] WLA[503] WLA[502] WLA[501] WLA[500] WLA[499] WLA[498] WLA[497] WLA[496]
+WLA[495] WLA[494] WLA[493] WLA[492] WLA[491] WLA[490] WLA[489] WLA[488] WLA[487] WLA[486]
+WLA[485] WLA[484] WLA[483] WLA[482] WLA[481] WLA[480] WLA[479] WLA[478] WLA[477] WLA[476]
+WLA[475] WLA[474] WLA[473] WLA[472] WLA[471] WLA[470] WLA[469] WLA[468] WLA[467] WLA[466]
+WLA[465] WLA[464] WLA[463] WLA[462] WLA[461] WLA[460] WLA[459] WLA[458] WLA[457] WLA[456]
+WLA[455] WLA[454] WLA[453] WLA[452] WLA[451] WLA[450] WLA[449] WLA[448] S55NLLGDPH_X512Y8D16_BW_BITCELL_ST68A_TOP_TW_RIGHT
XI16 BWENA[0] BWENB[0] CLKA CLKB CLKXA CLKXB DATAA[0] DATAB[0] DOUTA[0] DOUTB[0]
+STWLA VSS VSS VSS STWLB STWLB VSS VSS RWLA[0] RWLA[1]
+RWLB[0] RWLB[1] SACK1A SACK1B SACK4A SACK4B VDD VSS WEA WEB
+WLA[511] WLA[510] WLA[509] WLA[508] WLA[507] WLA[506] WLA[505] WLA[504] WLA[503] WLA[502]
+WLA[501] WLA[500] WLA[499] WLA[498] WLA[497] WLA[496] WLA[495] WLA[494] WLA[493] WLA[492]
+WLA[491] WLA[490] WLA[489] WLA[488] WLA[487] WLA[486] WLA[485] WLA[484] WLA[483] WLA[482]
+WLA[481] WLA[480] WLA[479] WLA[478] WLA[477] WLA[476] WLA[475] WLA[474] WLA[473] WLA[472]
+WLA[471] WLA[470] WLA[469] WLA[468] WLA[467] WLA[466] WLA[465] WLA[464] WLA[463] WLA[462]
+WLA[461] WLA[460] WLA[459] WLA[458] WLA[457] WLA[456] WLA[455] WLA[454] WLA[453] WLA[452]
+WLA[451] WLA[450] WLA[449] WLA[448] WLA[447] WLA[446] WLA[445] WLA[444] WLA[443] WLA[442]
+WLA[441] WLA[440] WLA[439] WLA[438] WLA[437] WLA[436] WLA[435] WLA[434] WLA[433] WLA[432]
+WLA[431] WLA[430] WLA[429] WLA[428] WLA[427] WLA[426] WLA[425] WLA[424] WLA[423] WLA[422]
+WLA[421] WLA[420] WLA[419] WLA[418] WLA[417] WLA[416] WLA[415] WLA[414] WLA[413] WLA[412]
+WLA[411] WLA[410] WLA[409] WLA[408] WLA[407] WLA[406] WLA[405] WLA[404] WLA[403] WLA[402]
+WLA[401] WLA[400] WLA[399] WLA[398] WLA[397] WLA[396] WLA[395] WLA[394] WLA[393] WLA[392]
+WLA[391] WLA[390] WLA[389] WLA[388] WLA[387] WLA[386] WLA[385] WLA[384] WLA[383] WLA[382]
+WLA[381] WLA[380] WLA[379] WLA[378] WLA[377] WLA[376] WLA[375] WLA[374] WLA[373] WLA[372]
+WLA[371] WLA[370] WLA[369] WLA[368] WLA[367] WLA[366] WLA[365] WLA[364] WLA[363] WLA[362]
+WLA[361] WLA[360] WLA[359] WLA[358] WLA[357] WLA[356] WLA[355] WLA[354] WLA[353] WLA[352]
+WLA[351] WLA[350] WLA[349] WLA[348] WLA[347] WLA[346] WLA[345] WLA[344] WLA[343] WLA[342]
+WLA[341] WLA[340] WLA[339] WLA[338] WLA[337] WLA[336] WLA[335] WLA[334] WLA[333] WLA[332]
+WLA[331] WLA[330] WLA[329] WLA[328] WLA[327] WLA[326] WLA[325] WLA[324] WLA[323] WLA[322]
+WLA[321] WLA[320] WLA[319] WLA[318] WLA[317] WLA[316] WLA[315] WLA[314] WLA[313] WLA[312]
+WLA[311] WLA[310] WLA[309] WLA[308] WLA[307] WLA[306] WLA[305] WLA[304] WLA[303] WLA[302]
+WLA[301] WLA[300] WLA[299] WLA[298] WLA[297] WLA[296] WLA[295] WLA[294] WLA[293] WLA[292]
+WLA[291] WLA[290] WLA[289] WLA[288] WLA[287] WLA[286] WLA[285] WLA[284] WLA[283] WLA[282]
+WLA[281] WLA[280] WLA[279] WLA[278] WLA[277] WLA[276] WLA[275] WLA[274] WLA[273] WLA[272]
+WLA[271] WLA[270] WLA[269] WLA[268] WLA[267] WLA[266] WLA[265] WLA[264] WLA[263] WLA[262]
+WLA[261] WLA[260] WLA[259] WLA[258] WLA[257] WLA[256] WLA[255] WLA[254] WLA[253] WLA[252]
+WLA[251] WLA[250] WLA[249] WLA[248] WLA[247] WLA[246] WLA[245] WLA[244] WLA[243] WLA[242]
+WLA[241] WLA[240] WLA[239] WLA[238] WLA[237] WLA[236] WLA[235] WLA[234] WLA[233] WLA[232]
+WLA[231] WLA[230] WLA[229] WLA[228] WLA[227] WLA[226] WLA[225] WLA[224] WLA[223] WLA[222]
+WLA[221] WLA[220] WLA[219] WLA[218] WLA[217] WLA[216] WLA[215] WLA[214] WLA[213] WLA[212]
+WLA[211] WLA[210] WLA[209] WLA[208] WLA[207] WLA[206] WLA[205] WLA[204] WLA[203] WLA[202]
+WLA[201] WLA[200] WLA[199] WLA[198] WLA[197] WLA[196] WLA[195] WLA[194] WLA[193] WLA[192]
+WLA[191] WLA[190] WLA[189] WLA[188] WLA[187] WLA[186] WLA[185] WLA[184] WLA[183] WLA[182]
+WLA[181] WLA[180] WLA[179] WLA[178] WLA[177] WLA[176] WLA[175] WLA[174] WLA[173] WLA[172]
+WLA[171] WLA[170] WLA[169] WLA[168] WLA[167] WLA[166] WLA[165] WLA[164] WLA[163] WLA[162]
+WLA[161] WLA[160] WLA[159] WLA[158] WLA[157] WLA[156] WLA[155] WLA[154] WLA[153] WLA[152]
+WLA[151] WLA[150] WLA[149] WLA[148] WLA[147] WLA[146] WLA[145] WLA[144] WLA[143] WLA[142]
+WLA[141] WLA[140] WLA[139] WLA[138] WLA[137] WLA[136] WLA[135] WLA[134] WLA[133] WLA[132]
+WLA[131] WLA[130] WLA[129] WLA[128] WLA[127] WLA[126] WLA[125] WLA[124] WLA[123] WLA[122]
+WLA[121] WLA[120] WLA[119] WLA[118] WLA[117] WLA[116] WLA[115] WLA[114] WLA[113] WLA[112]
+WLA[111] WLA[110] WLA[109] WLA[108] WLA[107] WLA[106] WLA[105] WLA[104] WLA[103] WLA[102]
+WLA[101] WLA[100] WLA[99] WLA[98] WLA[97] WLA[96] WLA[95] WLA[94] WLA[93] WLA[92]
+WLA[91] WLA[90] WLA[89] WLA[88] WLA[87] WLA[86] WLA[85] WLA[84] WLA[83] WLA[82]
+WLA[81] WLA[80] WLA[79] WLA[78] WLA[77] WLA[76] WLA[75] WLA[74] WLA[73] WLA[72]
+WLA[71] WLA[70] WLA[69] WLA[68] WLA[67] WLA[66] WLA[65] WLA[64] WLA[63] WLA[62]
+WLA[61] WLA[60] WLA[59] WLA[58] WLA[57] WLA[56] WLA[55] WLA[54] WLA[53] WLA[52]
+WLA[51] WLA[50] WLA[49] WLA[48] WLA[47] WLA[46] WLA[45] WLA[44] WLA[43] WLA[42]
+WLA[41] WLA[40] WLA[39] WLA[38] WLA[37] WLA[36] WLA[35] WLA[34] WLA[33] WLA[32]
+WLA[31] WLA[30] WLA[29] WLA[28] WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22]
+WLA[21] WLA[20] WLA[19] WLA[18] WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12]
+WLA[11] WLA[10] WLA[9] WLA[8] WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2]
+WLA[1] WLA[0] WLB[511] WLB[510] WLB[509] WLB[508] WLB[507] WLB[506] WLB[505] WLB[504]
+WLB[503] WLB[502] WLB[501] WLB[500] WLB[499] WLB[498] WLB[497] WLB[496] WLB[495] WLB[494]
+WLB[493] WLB[492] WLB[491] WLB[490] WLB[489] WLB[488] WLB[487] WLB[486] WLB[485] WLB[484]
+WLB[483] WLB[482] WLB[481] WLB[480] WLB[479] WLB[478] WLB[477] WLB[476] WLB[475] WLB[474]
+WLB[473] WLB[472] WLB[471] WLB[470] WLB[469] WLB[468] WLB[467] WLB[466] WLB[465] WLB[464]
+WLB[463] WLB[462] WLB[461] WLB[460] WLB[459] WLB[458] WLB[457] WLB[456] WLB[455] WLB[454]
+WLB[453] WLB[452] WLB[451] WLB[450] WLB[449] WLB[448] WLB[447] WLB[446] WLB[445] WLB[444]
+WLB[443] WLB[442] WLB[441] WLB[440] WLB[439] WLB[438] WLB[437] WLB[436] WLB[435] WLB[434]
+WLB[433] WLB[432] WLB[431] WLB[430] WLB[429] WLB[428] WLB[427] WLB[426] WLB[425] WLB[424]
+WLB[423] WLB[422] WLB[421] WLB[420] WLB[419] WLB[418] WLB[417] WLB[416] WLB[415] WLB[414]
+WLB[413] WLB[412] WLB[411] WLB[410] WLB[409] WLB[408] WLB[407] WLB[406] WLB[405] WLB[404]
+WLB[403] WLB[402] WLB[401] WLB[400] WLB[399] WLB[398] WLB[397] WLB[396] WLB[395] WLB[394]
+WLB[393] WLB[392] WLB[391] WLB[390] WLB[389] WLB[388] WLB[387] WLB[386] WLB[385] WLB[384]
+WLB[383] WLB[382] WLB[381] WLB[380] WLB[379] WLB[378] WLB[377] WLB[376] WLB[375] WLB[374]
+WLB[373] WLB[372] WLB[371] WLB[370] WLB[369] WLB[368] WLB[367] WLB[366] WLB[365] WLB[364]
+WLB[363] WLB[362] WLB[361] WLB[360] WLB[359] WLB[358] WLB[357] WLB[356] WLB[355] WLB[354]
+WLB[353] WLB[352] WLB[351] WLB[350] WLB[349] WLB[348] WLB[347] WLB[346] WLB[345] WLB[344]
+WLB[343] WLB[342] WLB[341] WLB[340] WLB[339] WLB[338] WLB[337] WLB[336] WLB[335] WLB[334]
+WLB[333] WLB[332] WLB[331] WLB[330] WLB[329] WLB[328] WLB[327] WLB[326] WLB[325] WLB[324]
+WLB[323] WLB[322] WLB[321] WLB[320] WLB[319] WLB[318] WLB[317] WLB[316] WLB[315] WLB[314]
+WLB[313] WLB[312] WLB[311] WLB[310] WLB[309] WLB[308] WLB[307] WLB[306] WLB[305] WLB[304]
+WLB[303] WLB[302] WLB[301] WLB[300] WLB[299] WLB[298] WLB[297] WLB[296] WLB[295] WLB[294]
+WLB[293] WLB[292] WLB[291] WLB[290] WLB[289] WLB[288] WLB[287] WLB[286] WLB[285] WLB[284]
+WLB[283] WLB[282] WLB[281] WLB[280] WLB[279] WLB[278] WLB[277] WLB[276] WLB[275] WLB[274]
+WLB[273] WLB[272] WLB[271] WLB[270] WLB[269] WLB[268] WLB[267] WLB[266] WLB[265] WLB[264]
+WLB[263] WLB[262] WLB[261] WLB[260] WLB[259] WLB[258] WLB[257] WLB[256] WLB[255] WLB[254]
+WLB[253] WLB[252] WLB[251] WLB[250] WLB[249] WLB[248] WLB[247] WLB[246] WLB[245] WLB[244]
+WLB[243] WLB[242] WLB[241] WLB[240] WLB[239] WLB[238] WLB[237] WLB[236] WLB[235] WLB[234]
+WLB[233] WLB[232] WLB[231] WLB[230] WLB[229] WLB[228] WLB[227] WLB[226] WLB[225] WLB[224]
+WLB[223] WLB[222] WLB[221] WLB[220] WLB[219] WLB[218] WLB[217] WLB[216] WLB[215] WLB[214]
+WLB[213] WLB[212] WLB[211] WLB[210] WLB[209] WLB[208] WLB[207] WLB[206] WLB[205] WLB[204]
+WLB[203] WLB[202] WLB[201] WLB[200] WLB[199] WLB[198] WLB[197] WLB[196] WLB[195] WLB[194]
+WLB[193] WLB[192] WLB[191] WLB[190] WLB[189] WLB[188] WLB[187] WLB[186] WLB[185] WLB[184]
+WLB[183] WLB[182] WLB[181] WLB[180] WLB[179] WLB[178] WLB[177] WLB[176] WLB[175] WLB[174]
+WLB[173] WLB[172] WLB[171] WLB[170] WLB[169] WLB[168] WLB[167] WLB[166] WLB[165] WLB[164]
+WLB[163] WLB[162] WLB[161] WLB[160] WLB[159] WLB[158] WLB[157] WLB[156] WLB[155] WLB[154]
+WLB[153] WLB[152] WLB[151] WLB[150] WLB[149] WLB[148] WLB[147] WLB[146] WLB[145] WLB[144]
+WLB[143] WLB[142] WLB[141] WLB[140] WLB[139] WLB[138] WLB[137] WLB[136] WLB[135] WLB[134]
+WLB[133] WLB[132] WLB[131] WLB[130] WLB[129] WLB[128] WLB[127] WLB[126] WLB[125] WLB[124]
+WLB[123] WLB[122] WLB[121] WLB[120] WLB[119] WLB[118] WLB[117] WLB[116] WLB[115] WLB[114]
+WLB[113] WLB[112] WLB[111] WLB[110] WLB[109] WLB[108] WLB[107] WLB[106] WLB[105] WLB[104]
+WLB[103] WLB[102] WLB[101] WLB[100] WLB[99] WLB[98] WLB[97] WLB[96] WLB[95] WLB[94]
+WLB[93] WLB[92] WLB[91] WLB[90] WLB[89] WLB[88] WLB[87] WLB[86] WLB[85] WLB[84]
+WLB[83] WLB[82] WLB[81] WLB[80] WLB[79] WLB[78] WLB[77] WLB[76] WLB[75] WLB[74]
+WLB[73] WLB[72] WLB[71] WLB[70] WLB[69] WLB[68] WLB[67] WLB[66] WLB[65] WLB[64]
+WLB[63] WLB[62] WLB[61] WLB[60] WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54]
+WLB[53] WLB[52] WLB[51] WLB[50] WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44]
+WLB[43] WLB[42] WLB[41] WLB[40] WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34]
+WLB[33] WLB[32] WLB[31] WLB[30] WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24]
+WLB[23] WLB[22] WLB[21] WLB[20] WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14]
+WLB[13] WLB[12] WLB[11] WLB[10] WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4]
+WLB[3] WLB[2] WLB[1] WLB[0] YXA[7] YXA[6] YXA[5] YXA[4] YXA[3] YXA[2]
+YXA[1] YXA[0] YXB[7] YXB[6] YXB[5] YXB[4] YXB[3] YXB[2] YXB[1] YXB[0] S55NLLGDPH_X512Y8D16_BW_Y512X8CELL_BW
XI17 BWENA[1] BWENB[1] CLKA CLKB CLKXA CLKXB DATAA[1] DATAB[1] DOUTA[1] DOUTB[1]
+STWLA VSS VSS VSS STWLB STWLB VSS VSS RWLA[0] RWLA[1]
+RWLB[0] RWLB[1] SACK1A SACK1B SACK4A SACK4B VDD VSS WEA WEB
+WLA[511] WLA[510] WLA[509] WLA[508] WLA[507] WLA[506] WLA[505] WLA[504] WLA[503] WLA[502]
+WLA[501] WLA[500] WLA[499] WLA[498] WLA[497] WLA[496] WLA[495] WLA[494] WLA[493] WLA[492]
+WLA[491] WLA[490] WLA[489] WLA[488] WLA[487] WLA[486] WLA[485] WLA[484] WLA[483] WLA[482]
+WLA[481] WLA[480] WLA[479] WLA[478] WLA[477] WLA[476] WLA[475] WLA[474] WLA[473] WLA[472]
+WLA[471] WLA[470] WLA[469] WLA[468] WLA[467] WLA[466] WLA[465] WLA[464] WLA[463] WLA[462]
+WLA[461] WLA[460] WLA[459] WLA[458] WLA[457] WLA[456] WLA[455] WLA[454] WLA[453] WLA[452]
+WLA[451] WLA[450] WLA[449] WLA[448] WLA[447] WLA[446] WLA[445] WLA[444] WLA[443] WLA[442]
+WLA[441] WLA[440] WLA[439] WLA[438] WLA[437] WLA[436] WLA[435] WLA[434] WLA[433] WLA[432]
+WLA[431] WLA[430] WLA[429] WLA[428] WLA[427] WLA[426] WLA[425] WLA[424] WLA[423] WLA[422]
+WLA[421] WLA[420] WLA[419] WLA[418] WLA[417] WLA[416] WLA[415] WLA[414] WLA[413] WLA[412]
+WLA[411] WLA[410] WLA[409] WLA[408] WLA[407] WLA[406] WLA[405] WLA[404] WLA[403] WLA[402]
+WLA[401] WLA[400] WLA[399] WLA[398] WLA[397] WLA[396] WLA[395] WLA[394] WLA[393] WLA[392]
+WLA[391] WLA[390] WLA[389] WLA[388] WLA[387] WLA[386] WLA[385] WLA[384] WLA[383] WLA[382]
+WLA[381] WLA[380] WLA[379] WLA[378] WLA[377] WLA[376] WLA[375] WLA[374] WLA[373] WLA[372]
+WLA[371] WLA[370] WLA[369] WLA[368] WLA[367] WLA[366] WLA[365] WLA[364] WLA[363] WLA[362]
+WLA[361] WLA[360] WLA[359] WLA[358] WLA[357] WLA[356] WLA[355] WLA[354] WLA[353] WLA[352]
+WLA[351] WLA[350] WLA[349] WLA[348] WLA[347] WLA[346] WLA[345] WLA[344] WLA[343] WLA[342]
+WLA[341] WLA[340] WLA[339] WLA[338] WLA[337] WLA[336] WLA[335] WLA[334] WLA[333] WLA[332]
+WLA[331] WLA[330] WLA[329] WLA[328] WLA[327] WLA[326] WLA[325] WLA[324] WLA[323] WLA[322]
+WLA[321] WLA[320] WLA[319] WLA[318] WLA[317] WLA[316] WLA[315] WLA[314] WLA[313] WLA[312]
+WLA[311] WLA[310] WLA[309] WLA[308] WLA[307] WLA[306] WLA[305] WLA[304] WLA[303] WLA[302]
+WLA[301] WLA[300] WLA[299] WLA[298] WLA[297] WLA[296] WLA[295] WLA[294] WLA[293] WLA[292]
+WLA[291] WLA[290] WLA[289] WLA[288] WLA[287] WLA[286] WLA[285] WLA[284] WLA[283] WLA[282]
+WLA[281] WLA[280] WLA[279] WLA[278] WLA[277] WLA[276] WLA[275] WLA[274] WLA[273] WLA[272]
+WLA[271] WLA[270] WLA[269] WLA[268] WLA[267] WLA[266] WLA[265] WLA[264] WLA[263] WLA[262]
+WLA[261] WLA[260] WLA[259] WLA[258] WLA[257] WLA[256] WLA[255] WLA[254] WLA[253] WLA[252]
+WLA[251] WLA[250] WLA[249] WLA[248] WLA[247] WLA[246] WLA[245] WLA[244] WLA[243] WLA[242]
+WLA[241] WLA[240] WLA[239] WLA[238] WLA[237] WLA[236] WLA[235] WLA[234] WLA[233] WLA[232]
+WLA[231] WLA[230] WLA[229] WLA[228] WLA[227] WLA[226] WLA[225] WLA[224] WLA[223] WLA[222]
+WLA[221] WLA[220] WLA[219] WLA[218] WLA[217] WLA[216] WLA[215] WLA[214] WLA[213] WLA[212]
+WLA[211] WLA[210] WLA[209] WLA[208] WLA[207] WLA[206] WLA[205] WLA[204] WLA[203] WLA[202]
+WLA[201] WLA[200] WLA[199] WLA[198] WLA[197] WLA[196] WLA[195] WLA[194] WLA[193] WLA[192]
+WLA[191] WLA[190] WLA[189] WLA[188] WLA[187] WLA[186] WLA[185] WLA[184] WLA[183] WLA[182]
+WLA[181] WLA[180] WLA[179] WLA[178] WLA[177] WLA[176] WLA[175] WLA[174] WLA[173] WLA[172]
+WLA[171] WLA[170] WLA[169] WLA[168] WLA[167] WLA[166] WLA[165] WLA[164] WLA[163] WLA[162]
+WLA[161] WLA[160] WLA[159] WLA[158] WLA[157] WLA[156] WLA[155] WLA[154] WLA[153] WLA[152]
+WLA[151] WLA[150] WLA[149] WLA[148] WLA[147] WLA[146] WLA[145] WLA[144] WLA[143] WLA[142]
+WLA[141] WLA[140] WLA[139] WLA[138] WLA[137] WLA[136] WLA[135] WLA[134] WLA[133] WLA[132]
+WLA[131] WLA[130] WLA[129] WLA[128] WLA[127] WLA[126] WLA[125] WLA[124] WLA[123] WLA[122]
+WLA[121] WLA[120] WLA[119] WLA[118] WLA[117] WLA[116] WLA[115] WLA[114] WLA[113] WLA[112]
+WLA[111] WLA[110] WLA[109] WLA[108] WLA[107] WLA[106] WLA[105] WLA[104] WLA[103] WLA[102]
+WLA[101] WLA[100] WLA[99] WLA[98] WLA[97] WLA[96] WLA[95] WLA[94] WLA[93] WLA[92]
+WLA[91] WLA[90] WLA[89] WLA[88] WLA[87] WLA[86] WLA[85] WLA[84] WLA[83] WLA[82]
+WLA[81] WLA[80] WLA[79] WLA[78] WLA[77] WLA[76] WLA[75] WLA[74] WLA[73] WLA[72]
+WLA[71] WLA[70] WLA[69] WLA[68] WLA[67] WLA[66] WLA[65] WLA[64] WLA[63] WLA[62]
+WLA[61] WLA[60] WLA[59] WLA[58] WLA[57] WLA[56] WLA[55] WLA[54] WLA[53] WLA[52]
+WLA[51] WLA[50] WLA[49] WLA[48] WLA[47] WLA[46] WLA[45] WLA[44] WLA[43] WLA[42]
+WLA[41] WLA[40] WLA[39] WLA[38] WLA[37] WLA[36] WLA[35] WLA[34] WLA[33] WLA[32]
+WLA[31] WLA[30] WLA[29] WLA[28] WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22]
+WLA[21] WLA[20] WLA[19] WLA[18] WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12]
+WLA[11] WLA[10] WLA[9] WLA[8] WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2]
+WLA[1] WLA[0] WLB[511] WLB[510] WLB[509] WLB[508] WLB[507] WLB[506] WLB[505] WLB[504]
+WLB[503] WLB[502] WLB[501] WLB[500] WLB[499] WLB[498] WLB[497] WLB[496] WLB[495] WLB[494]
+WLB[493] WLB[492] WLB[491] WLB[490] WLB[489] WLB[488] WLB[487] WLB[486] WLB[485] WLB[484]
+WLB[483] WLB[482] WLB[481] WLB[480] WLB[479] WLB[478] WLB[477] WLB[476] WLB[475] WLB[474]
+WLB[473] WLB[472] WLB[471] WLB[470] WLB[469] WLB[468] WLB[467] WLB[466] WLB[465] WLB[464]
+WLB[463] WLB[462] WLB[461] WLB[460] WLB[459] WLB[458] WLB[457] WLB[456] WLB[455] WLB[454]
+WLB[453] WLB[452] WLB[451] WLB[450] WLB[449] WLB[448] WLB[447] WLB[446] WLB[445] WLB[444]
+WLB[443] WLB[442] WLB[441] WLB[440] WLB[439] WLB[438] WLB[437] WLB[436] WLB[435] WLB[434]
+WLB[433] WLB[432] WLB[431] WLB[430] WLB[429] WLB[428] WLB[427] WLB[426] WLB[425] WLB[424]
+WLB[423] WLB[422] WLB[421] WLB[420] WLB[419] WLB[418] WLB[417] WLB[416] WLB[415] WLB[414]
+WLB[413] WLB[412] WLB[411] WLB[410] WLB[409] WLB[408] WLB[407] WLB[406] WLB[405] WLB[404]
+WLB[403] WLB[402] WLB[401] WLB[400] WLB[399] WLB[398] WLB[397] WLB[396] WLB[395] WLB[394]
+WLB[393] WLB[392] WLB[391] WLB[390] WLB[389] WLB[388] WLB[387] WLB[386] WLB[385] WLB[384]
+WLB[383] WLB[382] WLB[381] WLB[380] WLB[379] WLB[378] WLB[377] WLB[376] WLB[375] WLB[374]
+WLB[373] WLB[372] WLB[371] WLB[370] WLB[369] WLB[368] WLB[367] WLB[366] WLB[365] WLB[364]
+WLB[363] WLB[362] WLB[361] WLB[360] WLB[359] WLB[358] WLB[357] WLB[356] WLB[355] WLB[354]
+WLB[353] WLB[352] WLB[351] WLB[350] WLB[349] WLB[348] WLB[347] WLB[346] WLB[345] WLB[344]
+WLB[343] WLB[342] WLB[341] WLB[340] WLB[339] WLB[338] WLB[337] WLB[336] WLB[335] WLB[334]
+WLB[333] WLB[332] WLB[331] WLB[330] WLB[329] WLB[328] WLB[327] WLB[326] WLB[325] WLB[324]
+WLB[323] WLB[322] WLB[321] WLB[320] WLB[319] WLB[318] WLB[317] WLB[316] WLB[315] WLB[314]
+WLB[313] WLB[312] WLB[311] WLB[310] WLB[309] WLB[308] WLB[307] WLB[306] WLB[305] WLB[304]
+WLB[303] WLB[302] WLB[301] WLB[300] WLB[299] WLB[298] WLB[297] WLB[296] WLB[295] WLB[294]
+WLB[293] WLB[292] WLB[291] WLB[290] WLB[289] WLB[288] WLB[287] WLB[286] WLB[285] WLB[284]
+WLB[283] WLB[282] WLB[281] WLB[280] WLB[279] WLB[278] WLB[277] WLB[276] WLB[275] WLB[274]
+WLB[273] WLB[272] WLB[271] WLB[270] WLB[269] WLB[268] WLB[267] WLB[266] WLB[265] WLB[264]
+WLB[263] WLB[262] WLB[261] WLB[260] WLB[259] WLB[258] WLB[257] WLB[256] WLB[255] WLB[254]
+WLB[253] WLB[252] WLB[251] WLB[250] WLB[249] WLB[248] WLB[247] WLB[246] WLB[245] WLB[244]
+WLB[243] WLB[242] WLB[241] WLB[240] WLB[239] WLB[238] WLB[237] WLB[236] WLB[235] WLB[234]
+WLB[233] WLB[232] WLB[231] WLB[230] WLB[229] WLB[228] WLB[227] WLB[226] WLB[225] WLB[224]
+WLB[223] WLB[222] WLB[221] WLB[220] WLB[219] WLB[218] WLB[217] WLB[216] WLB[215] WLB[214]
+WLB[213] WLB[212] WLB[211] WLB[210] WLB[209] WLB[208] WLB[207] WLB[206] WLB[205] WLB[204]
+WLB[203] WLB[202] WLB[201] WLB[200] WLB[199] WLB[198] WLB[197] WLB[196] WLB[195] WLB[194]
+WLB[193] WLB[192] WLB[191] WLB[190] WLB[189] WLB[188] WLB[187] WLB[186] WLB[185] WLB[184]
+WLB[183] WLB[182] WLB[181] WLB[180] WLB[179] WLB[178] WLB[177] WLB[176] WLB[175] WLB[174]
+WLB[173] WLB[172] WLB[171] WLB[170] WLB[169] WLB[168] WLB[167] WLB[166] WLB[165] WLB[164]
+WLB[163] WLB[162] WLB[161] WLB[160] WLB[159] WLB[158] WLB[157] WLB[156] WLB[155] WLB[154]
+WLB[153] WLB[152] WLB[151] WLB[150] WLB[149] WLB[148] WLB[147] WLB[146] WLB[145] WLB[144]
+WLB[143] WLB[142] WLB[141] WLB[140] WLB[139] WLB[138] WLB[137] WLB[136] WLB[135] WLB[134]
+WLB[133] WLB[132] WLB[131] WLB[130] WLB[129] WLB[128] WLB[127] WLB[126] WLB[125] WLB[124]
+WLB[123] WLB[122] WLB[121] WLB[120] WLB[119] WLB[118] WLB[117] WLB[116] WLB[115] WLB[114]
+WLB[113] WLB[112] WLB[111] WLB[110] WLB[109] WLB[108] WLB[107] WLB[106] WLB[105] WLB[104]
+WLB[103] WLB[102] WLB[101] WLB[100] WLB[99] WLB[98] WLB[97] WLB[96] WLB[95] WLB[94]
+WLB[93] WLB[92] WLB[91] WLB[90] WLB[89] WLB[88] WLB[87] WLB[86] WLB[85] WLB[84]
+WLB[83] WLB[82] WLB[81] WLB[80] WLB[79] WLB[78] WLB[77] WLB[76] WLB[75] WLB[74]
+WLB[73] WLB[72] WLB[71] WLB[70] WLB[69] WLB[68] WLB[67] WLB[66] WLB[65] WLB[64]
+WLB[63] WLB[62] WLB[61] WLB[60] WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54]
+WLB[53] WLB[52] WLB[51] WLB[50] WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44]
+WLB[43] WLB[42] WLB[41] WLB[40] WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34]
+WLB[33] WLB[32] WLB[31] WLB[30] WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24]
+WLB[23] WLB[22] WLB[21] WLB[20] WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14]
+WLB[13] WLB[12] WLB[11] WLB[10] WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4]
+WLB[3] WLB[2] WLB[1] WLB[0] YXA[7] YXA[6] YXA[5] YXA[4] YXA[3] YXA[2]
+YXA[1] YXA[0] YXB[7] YXB[6] YXB[5] YXB[4] YXB[3] YXB[2] YXB[1] YXB[0] S55NLLGDPH_X512Y8D16_BW_Y512X8CELL_BW
XI18 BWENA[2] BWENB[2] CLKA CLKB CLKXA CLKXB DATAA[2] DATAB[2] DOUTA[2] DOUTB[2]
+STWLA VSS VSS VSS STWLB STWLB VSS VSS RWLA[0] RWLA[1]
+RWLB[0] RWLB[1] SACK1A SACK1B SACK4A SACK4B VDD VSS WEA WEB
+WLA[511] WLA[510] WLA[509] WLA[508] WLA[507] WLA[506] WLA[505] WLA[504] WLA[503] WLA[502]
+WLA[501] WLA[500] WLA[499] WLA[498] WLA[497] WLA[496] WLA[495] WLA[494] WLA[493] WLA[492]
+WLA[491] WLA[490] WLA[489] WLA[488] WLA[487] WLA[486] WLA[485] WLA[484] WLA[483] WLA[482]
+WLA[481] WLA[480] WLA[479] WLA[478] WLA[477] WLA[476] WLA[475] WLA[474] WLA[473] WLA[472]
+WLA[471] WLA[470] WLA[469] WLA[468] WLA[467] WLA[466] WLA[465] WLA[464] WLA[463] WLA[462]
+WLA[461] WLA[460] WLA[459] WLA[458] WLA[457] WLA[456] WLA[455] WLA[454] WLA[453] WLA[452]
+WLA[451] WLA[450] WLA[449] WLA[448] WLA[447] WLA[446] WLA[445] WLA[444] WLA[443] WLA[442]
+WLA[441] WLA[440] WLA[439] WLA[438] WLA[437] WLA[436] WLA[435] WLA[434] WLA[433] WLA[432]
+WLA[431] WLA[430] WLA[429] WLA[428] WLA[427] WLA[426] WLA[425] WLA[424] WLA[423] WLA[422]
+WLA[421] WLA[420] WLA[419] WLA[418] WLA[417] WLA[416] WLA[415] WLA[414] WLA[413] WLA[412]
+WLA[411] WLA[410] WLA[409] WLA[408] WLA[407] WLA[406] WLA[405] WLA[404] WLA[403] WLA[402]
+WLA[401] WLA[400] WLA[399] WLA[398] WLA[397] WLA[396] WLA[395] WLA[394] WLA[393] WLA[392]
+WLA[391] WLA[390] WLA[389] WLA[388] WLA[387] WLA[386] WLA[385] WLA[384] WLA[383] WLA[382]
+WLA[381] WLA[380] WLA[379] WLA[378] WLA[377] WLA[376] WLA[375] WLA[374] WLA[373] WLA[372]
+WLA[371] WLA[370] WLA[369] WLA[368] WLA[367] WLA[366] WLA[365] WLA[364] WLA[363] WLA[362]
+WLA[361] WLA[360] WLA[359] WLA[358] WLA[357] WLA[356] WLA[355] WLA[354] WLA[353] WLA[352]
+WLA[351] WLA[350] WLA[349] WLA[348] WLA[347] WLA[346] WLA[345] WLA[344] WLA[343] WLA[342]
+WLA[341] WLA[340] WLA[339] WLA[338] WLA[337] WLA[336] WLA[335] WLA[334] WLA[333] WLA[332]
+WLA[331] WLA[330] WLA[329] WLA[328] WLA[327] WLA[326] WLA[325] WLA[324] WLA[323] WLA[322]
+WLA[321] WLA[320] WLA[319] WLA[318] WLA[317] WLA[316] WLA[315] WLA[314] WLA[313] WLA[312]
+WLA[311] WLA[310] WLA[309] WLA[308] WLA[307] WLA[306] WLA[305] WLA[304] WLA[303] WLA[302]
+WLA[301] WLA[300] WLA[299] WLA[298] WLA[297] WLA[296] WLA[295] WLA[294] WLA[293] WLA[292]
+WLA[291] WLA[290] WLA[289] WLA[288] WLA[287] WLA[286] WLA[285] WLA[284] WLA[283] WLA[282]
+WLA[281] WLA[280] WLA[279] WLA[278] WLA[277] WLA[276] WLA[275] WLA[274] WLA[273] WLA[272]
+WLA[271] WLA[270] WLA[269] WLA[268] WLA[267] WLA[266] WLA[265] WLA[264] WLA[263] WLA[262]
+WLA[261] WLA[260] WLA[259] WLA[258] WLA[257] WLA[256] WLA[255] WLA[254] WLA[253] WLA[252]
+WLA[251] WLA[250] WLA[249] WLA[248] WLA[247] WLA[246] WLA[245] WLA[244] WLA[243] WLA[242]
+WLA[241] WLA[240] WLA[239] WLA[238] WLA[237] WLA[236] WLA[235] WLA[234] WLA[233] WLA[232]
+WLA[231] WLA[230] WLA[229] WLA[228] WLA[227] WLA[226] WLA[225] WLA[224] WLA[223] WLA[222]
+WLA[221] WLA[220] WLA[219] WLA[218] WLA[217] WLA[216] WLA[215] WLA[214] WLA[213] WLA[212]
+WLA[211] WLA[210] WLA[209] WLA[208] WLA[207] WLA[206] WLA[205] WLA[204] WLA[203] WLA[202]
+WLA[201] WLA[200] WLA[199] WLA[198] WLA[197] WLA[196] WLA[195] WLA[194] WLA[193] WLA[192]
+WLA[191] WLA[190] WLA[189] WLA[188] WLA[187] WLA[186] WLA[185] WLA[184] WLA[183] WLA[182]
+WLA[181] WLA[180] WLA[179] WLA[178] WLA[177] WLA[176] WLA[175] WLA[174] WLA[173] WLA[172]
+WLA[171] WLA[170] WLA[169] WLA[168] WLA[167] WLA[166] WLA[165] WLA[164] WLA[163] WLA[162]
+WLA[161] WLA[160] WLA[159] WLA[158] WLA[157] WLA[156] WLA[155] WLA[154] WLA[153] WLA[152]
+WLA[151] WLA[150] WLA[149] WLA[148] WLA[147] WLA[146] WLA[145] WLA[144] WLA[143] WLA[142]
+WLA[141] WLA[140] WLA[139] WLA[138] WLA[137] WLA[136] WLA[135] WLA[134] WLA[133] WLA[132]
+WLA[131] WLA[130] WLA[129] WLA[128] WLA[127] WLA[126] WLA[125] WLA[124] WLA[123] WLA[122]
+WLA[121] WLA[120] WLA[119] WLA[118] WLA[117] WLA[116] WLA[115] WLA[114] WLA[113] WLA[112]
+WLA[111] WLA[110] WLA[109] WLA[108] WLA[107] WLA[106] WLA[105] WLA[104] WLA[103] WLA[102]
+WLA[101] WLA[100] WLA[99] WLA[98] WLA[97] WLA[96] WLA[95] WLA[94] WLA[93] WLA[92]
+WLA[91] WLA[90] WLA[89] WLA[88] WLA[87] WLA[86] WLA[85] WLA[84] WLA[83] WLA[82]
+WLA[81] WLA[80] WLA[79] WLA[78] WLA[77] WLA[76] WLA[75] WLA[74] WLA[73] WLA[72]
+WLA[71] WLA[70] WLA[69] WLA[68] WLA[67] WLA[66] WLA[65] WLA[64] WLA[63] WLA[62]
+WLA[61] WLA[60] WLA[59] WLA[58] WLA[57] WLA[56] WLA[55] WLA[54] WLA[53] WLA[52]
+WLA[51] WLA[50] WLA[49] WLA[48] WLA[47] WLA[46] WLA[45] WLA[44] WLA[43] WLA[42]
+WLA[41] WLA[40] WLA[39] WLA[38] WLA[37] WLA[36] WLA[35] WLA[34] WLA[33] WLA[32]
+WLA[31] WLA[30] WLA[29] WLA[28] WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22]
+WLA[21] WLA[20] WLA[19] WLA[18] WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12]
+WLA[11] WLA[10] WLA[9] WLA[8] WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2]
+WLA[1] WLA[0] WLB[511] WLB[510] WLB[509] WLB[508] WLB[507] WLB[506] WLB[505] WLB[504]
+WLB[503] WLB[502] WLB[501] WLB[500] WLB[499] WLB[498] WLB[497] WLB[496] WLB[495] WLB[494]
+WLB[493] WLB[492] WLB[491] WLB[490] WLB[489] WLB[488] WLB[487] WLB[486] WLB[485] WLB[484]
+WLB[483] WLB[482] WLB[481] WLB[480] WLB[479] WLB[478] WLB[477] WLB[476] WLB[475] WLB[474]
+WLB[473] WLB[472] WLB[471] WLB[470] WLB[469] WLB[468] WLB[467] WLB[466] WLB[465] WLB[464]
+WLB[463] WLB[462] WLB[461] WLB[460] WLB[459] WLB[458] WLB[457] WLB[456] WLB[455] WLB[454]
+WLB[453] WLB[452] WLB[451] WLB[450] WLB[449] WLB[448] WLB[447] WLB[446] WLB[445] WLB[444]
+WLB[443] WLB[442] WLB[441] WLB[440] WLB[439] WLB[438] WLB[437] WLB[436] WLB[435] WLB[434]
+WLB[433] WLB[432] WLB[431] WLB[430] WLB[429] WLB[428] WLB[427] WLB[426] WLB[425] WLB[424]
+WLB[423] WLB[422] WLB[421] WLB[420] WLB[419] WLB[418] WLB[417] WLB[416] WLB[415] WLB[414]
+WLB[413] WLB[412] WLB[411] WLB[410] WLB[409] WLB[408] WLB[407] WLB[406] WLB[405] WLB[404]
+WLB[403] WLB[402] WLB[401] WLB[400] WLB[399] WLB[398] WLB[397] WLB[396] WLB[395] WLB[394]
+WLB[393] WLB[392] WLB[391] WLB[390] WLB[389] WLB[388] WLB[387] WLB[386] WLB[385] WLB[384]
+WLB[383] WLB[382] WLB[381] WLB[380] WLB[379] WLB[378] WLB[377] WLB[376] WLB[375] WLB[374]
+WLB[373] WLB[372] WLB[371] WLB[370] WLB[369] WLB[368] WLB[367] WLB[366] WLB[365] WLB[364]
+WLB[363] WLB[362] WLB[361] WLB[360] WLB[359] WLB[358] WLB[357] WLB[356] WLB[355] WLB[354]
+WLB[353] WLB[352] WLB[351] WLB[350] WLB[349] WLB[348] WLB[347] WLB[346] WLB[345] WLB[344]
+WLB[343] WLB[342] WLB[341] WLB[340] WLB[339] WLB[338] WLB[337] WLB[336] WLB[335] WLB[334]
+WLB[333] WLB[332] WLB[331] WLB[330] WLB[329] WLB[328] WLB[327] WLB[326] WLB[325] WLB[324]
+WLB[323] WLB[322] WLB[321] WLB[320] WLB[319] WLB[318] WLB[317] WLB[316] WLB[315] WLB[314]
+WLB[313] WLB[312] WLB[311] WLB[310] WLB[309] WLB[308] WLB[307] WLB[306] WLB[305] WLB[304]
+WLB[303] WLB[302] WLB[301] WLB[300] WLB[299] WLB[298] WLB[297] WLB[296] WLB[295] WLB[294]
+WLB[293] WLB[292] WLB[291] WLB[290] WLB[289] WLB[288] WLB[287] WLB[286] WLB[285] WLB[284]
+WLB[283] WLB[282] WLB[281] WLB[280] WLB[279] WLB[278] WLB[277] WLB[276] WLB[275] WLB[274]
+WLB[273] WLB[272] WLB[271] WLB[270] WLB[269] WLB[268] WLB[267] WLB[266] WLB[265] WLB[264]
+WLB[263] WLB[262] WLB[261] WLB[260] WLB[259] WLB[258] WLB[257] WLB[256] WLB[255] WLB[254]
+WLB[253] WLB[252] WLB[251] WLB[250] WLB[249] WLB[248] WLB[247] WLB[246] WLB[245] WLB[244]
+WLB[243] WLB[242] WLB[241] WLB[240] WLB[239] WLB[238] WLB[237] WLB[236] WLB[235] WLB[234]
+WLB[233] WLB[232] WLB[231] WLB[230] WLB[229] WLB[228] WLB[227] WLB[226] WLB[225] WLB[224]
+WLB[223] WLB[222] WLB[221] WLB[220] WLB[219] WLB[218] WLB[217] WLB[216] WLB[215] WLB[214]
+WLB[213] WLB[212] WLB[211] WLB[210] WLB[209] WLB[208] WLB[207] WLB[206] WLB[205] WLB[204]
+WLB[203] WLB[202] WLB[201] WLB[200] WLB[199] WLB[198] WLB[197] WLB[196] WLB[195] WLB[194]
+WLB[193] WLB[192] WLB[191] WLB[190] WLB[189] WLB[188] WLB[187] WLB[186] WLB[185] WLB[184]
+WLB[183] WLB[182] WLB[181] WLB[180] WLB[179] WLB[178] WLB[177] WLB[176] WLB[175] WLB[174]
+WLB[173] WLB[172] WLB[171] WLB[170] WLB[169] WLB[168] WLB[167] WLB[166] WLB[165] WLB[164]
+WLB[163] WLB[162] WLB[161] WLB[160] WLB[159] WLB[158] WLB[157] WLB[156] WLB[155] WLB[154]
+WLB[153] WLB[152] WLB[151] WLB[150] WLB[149] WLB[148] WLB[147] WLB[146] WLB[145] WLB[144]
+WLB[143] WLB[142] WLB[141] WLB[140] WLB[139] WLB[138] WLB[137] WLB[136] WLB[135] WLB[134]
+WLB[133] WLB[132] WLB[131] WLB[130] WLB[129] WLB[128] WLB[127] WLB[126] WLB[125] WLB[124]
+WLB[123] WLB[122] WLB[121] WLB[120] WLB[119] WLB[118] WLB[117] WLB[116] WLB[115] WLB[114]
+WLB[113] WLB[112] WLB[111] WLB[110] WLB[109] WLB[108] WLB[107] WLB[106] WLB[105] WLB[104]
+WLB[103] WLB[102] WLB[101] WLB[100] WLB[99] WLB[98] WLB[97] WLB[96] WLB[95] WLB[94]
+WLB[93] WLB[92] WLB[91] WLB[90] WLB[89] WLB[88] WLB[87] WLB[86] WLB[85] WLB[84]
+WLB[83] WLB[82] WLB[81] WLB[80] WLB[79] WLB[78] WLB[77] WLB[76] WLB[75] WLB[74]
+WLB[73] WLB[72] WLB[71] WLB[70] WLB[69] WLB[68] WLB[67] WLB[66] WLB[65] WLB[64]
+WLB[63] WLB[62] WLB[61] WLB[60] WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54]
+WLB[53] WLB[52] WLB[51] WLB[50] WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44]
+WLB[43] WLB[42] WLB[41] WLB[40] WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34]
+WLB[33] WLB[32] WLB[31] WLB[30] WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24]
+WLB[23] WLB[22] WLB[21] WLB[20] WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14]
+WLB[13] WLB[12] WLB[11] WLB[10] WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4]
+WLB[3] WLB[2] WLB[1] WLB[0] YXA[7] YXA[6] YXA[5] YXA[4] YXA[3] YXA[2]
+YXA[1] YXA[0] YXB[7] YXB[6] YXB[5] YXB[4] YXB[3] YXB[2] YXB[1] YXB[0] S55NLLGDPH_X512Y8D16_BW_Y512X8CELL_BW
XI19 BWENA[3] BWENB[3] CLKA CLKB CLKXA CLKXB DATAA[3] DATAB[3] DOUTA[3] DOUTB[3]
+STWLA VSS VSS VSS STWLB STWLB VSS VSS RWLA[0] RWLA[1]
+RWLB[0] RWLB[1] SACK1A SACK1B SACK4A SACK4B VDD VSS WEA WEB
+WLA[511] WLA[510] WLA[509] WLA[508] WLA[507] WLA[506] WLA[505] WLA[504] WLA[503] WLA[502]
+WLA[501] WLA[500] WLA[499] WLA[498] WLA[497] WLA[496] WLA[495] WLA[494] WLA[493] WLA[492]
+WLA[491] WLA[490] WLA[489] WLA[488] WLA[487] WLA[486] WLA[485] WLA[484] WLA[483] WLA[482]
+WLA[481] WLA[480] WLA[479] WLA[478] WLA[477] WLA[476] WLA[475] WLA[474] WLA[473] WLA[472]
+WLA[471] WLA[470] WLA[469] WLA[468] WLA[467] WLA[466] WLA[465] WLA[464] WLA[463] WLA[462]
+WLA[461] WLA[460] WLA[459] WLA[458] WLA[457] WLA[456] WLA[455] WLA[454] WLA[453] WLA[452]
+WLA[451] WLA[450] WLA[449] WLA[448] WLA[447] WLA[446] WLA[445] WLA[444] WLA[443] WLA[442]
+WLA[441] WLA[440] WLA[439] WLA[438] WLA[437] WLA[436] WLA[435] WLA[434] WLA[433] WLA[432]
+WLA[431] WLA[430] WLA[429] WLA[428] WLA[427] WLA[426] WLA[425] WLA[424] WLA[423] WLA[422]
+WLA[421] WLA[420] WLA[419] WLA[418] WLA[417] WLA[416] WLA[415] WLA[414] WLA[413] WLA[412]
+WLA[411] WLA[410] WLA[409] WLA[408] WLA[407] WLA[406] WLA[405] WLA[404] WLA[403] WLA[402]
+WLA[401] WLA[400] WLA[399] WLA[398] WLA[397] WLA[396] WLA[395] WLA[394] WLA[393] WLA[392]
+WLA[391] WLA[390] WLA[389] WLA[388] WLA[387] WLA[386] WLA[385] WLA[384] WLA[383] WLA[382]
+WLA[381] WLA[380] WLA[379] WLA[378] WLA[377] WLA[376] WLA[375] WLA[374] WLA[373] WLA[372]
+WLA[371] WLA[370] WLA[369] WLA[368] WLA[367] WLA[366] WLA[365] WLA[364] WLA[363] WLA[362]
+WLA[361] WLA[360] WLA[359] WLA[358] WLA[357] WLA[356] WLA[355] WLA[354] WLA[353] WLA[352]
+WLA[351] WLA[350] WLA[349] WLA[348] WLA[347] WLA[346] WLA[345] WLA[344] WLA[343] WLA[342]
+WLA[341] WLA[340] WLA[339] WLA[338] WLA[337] WLA[336] WLA[335] WLA[334] WLA[333] WLA[332]
+WLA[331] WLA[330] WLA[329] WLA[328] WLA[327] WLA[326] WLA[325] WLA[324] WLA[323] WLA[322]
+WLA[321] WLA[320] WLA[319] WLA[318] WLA[317] WLA[316] WLA[315] WLA[314] WLA[313] WLA[312]
+WLA[311] WLA[310] WLA[309] WLA[308] WLA[307] WLA[306] WLA[305] WLA[304] WLA[303] WLA[302]
+WLA[301] WLA[300] WLA[299] WLA[298] WLA[297] WLA[296] WLA[295] WLA[294] WLA[293] WLA[292]
+WLA[291] WLA[290] WLA[289] WLA[288] WLA[287] WLA[286] WLA[285] WLA[284] WLA[283] WLA[282]
+WLA[281] WLA[280] WLA[279] WLA[278] WLA[277] WLA[276] WLA[275] WLA[274] WLA[273] WLA[272]
+WLA[271] WLA[270] WLA[269] WLA[268] WLA[267] WLA[266] WLA[265] WLA[264] WLA[263] WLA[262]
+WLA[261] WLA[260] WLA[259] WLA[258] WLA[257] WLA[256] WLA[255] WLA[254] WLA[253] WLA[252]
+WLA[251] WLA[250] WLA[249] WLA[248] WLA[247] WLA[246] WLA[245] WLA[244] WLA[243] WLA[242]
+WLA[241] WLA[240] WLA[239] WLA[238] WLA[237] WLA[236] WLA[235] WLA[234] WLA[233] WLA[232]
+WLA[231] WLA[230] WLA[229] WLA[228] WLA[227] WLA[226] WLA[225] WLA[224] WLA[223] WLA[222]
+WLA[221] WLA[220] WLA[219] WLA[218] WLA[217] WLA[216] WLA[215] WLA[214] WLA[213] WLA[212]
+WLA[211] WLA[210] WLA[209] WLA[208] WLA[207] WLA[206] WLA[205] WLA[204] WLA[203] WLA[202]
+WLA[201] WLA[200] WLA[199] WLA[198] WLA[197] WLA[196] WLA[195] WLA[194] WLA[193] WLA[192]
+WLA[191] WLA[190] WLA[189] WLA[188] WLA[187] WLA[186] WLA[185] WLA[184] WLA[183] WLA[182]
+WLA[181] WLA[180] WLA[179] WLA[178] WLA[177] WLA[176] WLA[175] WLA[174] WLA[173] WLA[172]
+WLA[171] WLA[170] WLA[169] WLA[168] WLA[167] WLA[166] WLA[165] WLA[164] WLA[163] WLA[162]
+WLA[161] WLA[160] WLA[159] WLA[158] WLA[157] WLA[156] WLA[155] WLA[154] WLA[153] WLA[152]
+WLA[151] WLA[150] WLA[149] WLA[148] WLA[147] WLA[146] WLA[145] WLA[144] WLA[143] WLA[142]
+WLA[141] WLA[140] WLA[139] WLA[138] WLA[137] WLA[136] WLA[135] WLA[134] WLA[133] WLA[132]
+WLA[131] WLA[130] WLA[129] WLA[128] WLA[127] WLA[126] WLA[125] WLA[124] WLA[123] WLA[122]
+WLA[121] WLA[120] WLA[119] WLA[118] WLA[117] WLA[116] WLA[115] WLA[114] WLA[113] WLA[112]
+WLA[111] WLA[110] WLA[109] WLA[108] WLA[107] WLA[106] WLA[105] WLA[104] WLA[103] WLA[102]
+WLA[101] WLA[100] WLA[99] WLA[98] WLA[97] WLA[96] WLA[95] WLA[94] WLA[93] WLA[92]
+WLA[91] WLA[90] WLA[89] WLA[88] WLA[87] WLA[86] WLA[85] WLA[84] WLA[83] WLA[82]
+WLA[81] WLA[80] WLA[79] WLA[78] WLA[77] WLA[76] WLA[75] WLA[74] WLA[73] WLA[72]
+WLA[71] WLA[70] WLA[69] WLA[68] WLA[67] WLA[66] WLA[65] WLA[64] WLA[63] WLA[62]
+WLA[61] WLA[60] WLA[59] WLA[58] WLA[57] WLA[56] WLA[55] WLA[54] WLA[53] WLA[52]
+WLA[51] WLA[50] WLA[49] WLA[48] WLA[47] WLA[46] WLA[45] WLA[44] WLA[43] WLA[42]
+WLA[41] WLA[40] WLA[39] WLA[38] WLA[37] WLA[36] WLA[35] WLA[34] WLA[33] WLA[32]
+WLA[31] WLA[30] WLA[29] WLA[28] WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22]
+WLA[21] WLA[20] WLA[19] WLA[18] WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12]
+WLA[11] WLA[10] WLA[9] WLA[8] WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2]
+WLA[1] WLA[0] WLB[511] WLB[510] WLB[509] WLB[508] WLB[507] WLB[506] WLB[505] WLB[504]
+WLB[503] WLB[502] WLB[501] WLB[500] WLB[499] WLB[498] WLB[497] WLB[496] WLB[495] WLB[494]
+WLB[493] WLB[492] WLB[491] WLB[490] WLB[489] WLB[488] WLB[487] WLB[486] WLB[485] WLB[484]
+WLB[483] WLB[482] WLB[481] WLB[480] WLB[479] WLB[478] WLB[477] WLB[476] WLB[475] WLB[474]
+WLB[473] WLB[472] WLB[471] WLB[470] WLB[469] WLB[468] WLB[467] WLB[466] WLB[465] WLB[464]
+WLB[463] WLB[462] WLB[461] WLB[460] WLB[459] WLB[458] WLB[457] WLB[456] WLB[455] WLB[454]
+WLB[453] WLB[452] WLB[451] WLB[450] WLB[449] WLB[448] WLB[447] WLB[446] WLB[445] WLB[444]
+WLB[443] WLB[442] WLB[441] WLB[440] WLB[439] WLB[438] WLB[437] WLB[436] WLB[435] WLB[434]
+WLB[433] WLB[432] WLB[431] WLB[430] WLB[429] WLB[428] WLB[427] WLB[426] WLB[425] WLB[424]
+WLB[423] WLB[422] WLB[421] WLB[420] WLB[419] WLB[418] WLB[417] WLB[416] WLB[415] WLB[414]
+WLB[413] WLB[412] WLB[411] WLB[410] WLB[409] WLB[408] WLB[407] WLB[406] WLB[405] WLB[404]
+WLB[403] WLB[402] WLB[401] WLB[400] WLB[399] WLB[398] WLB[397] WLB[396] WLB[395] WLB[394]
+WLB[393] WLB[392] WLB[391] WLB[390] WLB[389] WLB[388] WLB[387] WLB[386] WLB[385] WLB[384]
+WLB[383] WLB[382] WLB[381] WLB[380] WLB[379] WLB[378] WLB[377] WLB[376] WLB[375] WLB[374]
+WLB[373] WLB[372] WLB[371] WLB[370] WLB[369] WLB[368] WLB[367] WLB[366] WLB[365] WLB[364]
+WLB[363] WLB[362] WLB[361] WLB[360] WLB[359] WLB[358] WLB[357] WLB[356] WLB[355] WLB[354]
+WLB[353] WLB[352] WLB[351] WLB[350] WLB[349] WLB[348] WLB[347] WLB[346] WLB[345] WLB[344]
+WLB[343] WLB[342] WLB[341] WLB[340] WLB[339] WLB[338] WLB[337] WLB[336] WLB[335] WLB[334]
+WLB[333] WLB[332] WLB[331] WLB[330] WLB[329] WLB[328] WLB[327] WLB[326] WLB[325] WLB[324]
+WLB[323] WLB[322] WLB[321] WLB[320] WLB[319] WLB[318] WLB[317] WLB[316] WLB[315] WLB[314]
+WLB[313] WLB[312] WLB[311] WLB[310] WLB[309] WLB[308] WLB[307] WLB[306] WLB[305] WLB[304]
+WLB[303] WLB[302] WLB[301] WLB[300] WLB[299] WLB[298] WLB[297] WLB[296] WLB[295] WLB[294]
+WLB[293] WLB[292] WLB[291] WLB[290] WLB[289] WLB[288] WLB[287] WLB[286] WLB[285] WLB[284]
+WLB[283] WLB[282] WLB[281] WLB[280] WLB[279] WLB[278] WLB[277] WLB[276] WLB[275] WLB[274]
+WLB[273] WLB[272] WLB[271] WLB[270] WLB[269] WLB[268] WLB[267] WLB[266] WLB[265] WLB[264]
+WLB[263] WLB[262] WLB[261] WLB[260] WLB[259] WLB[258] WLB[257] WLB[256] WLB[255] WLB[254]
+WLB[253] WLB[252] WLB[251] WLB[250] WLB[249] WLB[248] WLB[247] WLB[246] WLB[245] WLB[244]
+WLB[243] WLB[242] WLB[241] WLB[240] WLB[239] WLB[238] WLB[237] WLB[236] WLB[235] WLB[234]
+WLB[233] WLB[232] WLB[231] WLB[230] WLB[229] WLB[228] WLB[227] WLB[226] WLB[225] WLB[224]
+WLB[223] WLB[222] WLB[221] WLB[220] WLB[219] WLB[218] WLB[217] WLB[216] WLB[215] WLB[214]
+WLB[213] WLB[212] WLB[211] WLB[210] WLB[209] WLB[208] WLB[207] WLB[206] WLB[205] WLB[204]
+WLB[203] WLB[202] WLB[201] WLB[200] WLB[199] WLB[198] WLB[197] WLB[196] WLB[195] WLB[194]
+WLB[193] WLB[192] WLB[191] WLB[190] WLB[189] WLB[188] WLB[187] WLB[186] WLB[185] WLB[184]
+WLB[183] WLB[182] WLB[181] WLB[180] WLB[179] WLB[178] WLB[177] WLB[176] WLB[175] WLB[174]
+WLB[173] WLB[172] WLB[171] WLB[170] WLB[169] WLB[168] WLB[167] WLB[166] WLB[165] WLB[164]
+WLB[163] WLB[162] WLB[161] WLB[160] WLB[159] WLB[158] WLB[157] WLB[156] WLB[155] WLB[154]
+WLB[153] WLB[152] WLB[151] WLB[150] WLB[149] WLB[148] WLB[147] WLB[146] WLB[145] WLB[144]
+WLB[143] WLB[142] WLB[141] WLB[140] WLB[139] WLB[138] WLB[137] WLB[136] WLB[135] WLB[134]
+WLB[133] WLB[132] WLB[131] WLB[130] WLB[129] WLB[128] WLB[127] WLB[126] WLB[125] WLB[124]
+WLB[123] WLB[122] WLB[121] WLB[120] WLB[119] WLB[118] WLB[117] WLB[116] WLB[115] WLB[114]
+WLB[113] WLB[112] WLB[111] WLB[110] WLB[109] WLB[108] WLB[107] WLB[106] WLB[105] WLB[104]
+WLB[103] WLB[102] WLB[101] WLB[100] WLB[99] WLB[98] WLB[97] WLB[96] WLB[95] WLB[94]
+WLB[93] WLB[92] WLB[91] WLB[90] WLB[89] WLB[88] WLB[87] WLB[86] WLB[85] WLB[84]
+WLB[83] WLB[82] WLB[81] WLB[80] WLB[79] WLB[78] WLB[77] WLB[76] WLB[75] WLB[74]
+WLB[73] WLB[72] WLB[71] WLB[70] WLB[69] WLB[68] WLB[67] WLB[66] WLB[65] WLB[64]
+WLB[63] WLB[62] WLB[61] WLB[60] WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54]
+WLB[53] WLB[52] WLB[51] WLB[50] WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44]
+WLB[43] WLB[42] WLB[41] WLB[40] WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34]
+WLB[33] WLB[32] WLB[31] WLB[30] WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24]
+WLB[23] WLB[22] WLB[21] WLB[20] WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14]
+WLB[13] WLB[12] WLB[11] WLB[10] WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4]
+WLB[3] WLB[2] WLB[1] WLB[0] YXA[7] YXA[6] YXA[5] YXA[4] YXA[3] YXA[2]
+YXA[1] YXA[0] YXB[7] YXB[6] YXB[5] YXB[4] YXB[3] YXB[2] YXB[1] YXB[0] S55NLLGDPH_X512Y8D16_BW_Y512X8CELL_BW
XI20 BWENA[4] BWENB[4] CLKA CLKB CLKXA CLKXB DATAA[4] DATAB[4] DOUTA[4] DOUTB[4]
+STWLA VSS VSS VSS VSS VSS VSS VSS RWLA[0] RWLA[1]
+RWLB[0] RWLB[1] SACK1A SACK1B SACK4A SACK4B VDD VSS WEA WEB
+WLA[511] WLA[510] WLA[509] WLA[508] WLA[507] WLA[506] WLA[505] WLA[504] WLA[503] WLA[502]
+WLA[501] WLA[500] WLA[499] WLA[498] WLA[497] WLA[496] WLA[495] WLA[494] WLA[493] WLA[492]
+WLA[491] WLA[490] WLA[489] WLA[488] WLA[487] WLA[486] WLA[485] WLA[484] WLA[483] WLA[482]
+WLA[481] WLA[480] WLA[479] WLA[478] WLA[477] WLA[476] WLA[475] WLA[474] WLA[473] WLA[472]
+WLA[471] WLA[470] WLA[469] WLA[468] WLA[467] WLA[466] WLA[465] WLA[464] WLA[463] WLA[462]
+WLA[461] WLA[460] WLA[459] WLA[458] WLA[457] WLA[456] WLA[455] WLA[454] WLA[453] WLA[452]
+WLA[451] WLA[450] WLA[449] WLA[448] WLA[447] WLA[446] WLA[445] WLA[444] WLA[443] WLA[442]
+WLA[441] WLA[440] WLA[439] WLA[438] WLA[437] WLA[436] WLA[435] WLA[434] WLA[433] WLA[432]
+WLA[431] WLA[430] WLA[429] WLA[428] WLA[427] WLA[426] WLA[425] WLA[424] WLA[423] WLA[422]
+WLA[421] WLA[420] WLA[419] WLA[418] WLA[417] WLA[416] WLA[415] WLA[414] WLA[413] WLA[412]
+WLA[411] WLA[410] WLA[409] WLA[408] WLA[407] WLA[406] WLA[405] WLA[404] WLA[403] WLA[402]
+WLA[401] WLA[400] WLA[399] WLA[398] WLA[397] WLA[396] WLA[395] WLA[394] WLA[393] WLA[392]
+WLA[391] WLA[390] WLA[389] WLA[388] WLA[387] WLA[386] WLA[385] WLA[384] WLA[383] WLA[382]
+WLA[381] WLA[380] WLA[379] WLA[378] WLA[377] WLA[376] WLA[375] WLA[374] WLA[373] WLA[372]
+WLA[371] WLA[370] WLA[369] WLA[368] WLA[367] WLA[366] WLA[365] WLA[364] WLA[363] WLA[362]
+WLA[361] WLA[360] WLA[359] WLA[358] WLA[357] WLA[356] WLA[355] WLA[354] WLA[353] WLA[352]
+WLA[351] WLA[350] WLA[349] WLA[348] WLA[347] WLA[346] WLA[345] WLA[344] WLA[343] WLA[342]
+WLA[341] WLA[340] WLA[339] WLA[338] WLA[337] WLA[336] WLA[335] WLA[334] WLA[333] WLA[332]
+WLA[331] WLA[330] WLA[329] WLA[328] WLA[327] WLA[326] WLA[325] WLA[324] WLA[323] WLA[322]
+WLA[321] WLA[320] WLA[319] WLA[318] WLA[317] WLA[316] WLA[315] WLA[314] WLA[313] WLA[312]
+WLA[311] WLA[310] WLA[309] WLA[308] WLA[307] WLA[306] WLA[305] WLA[304] WLA[303] WLA[302]
+WLA[301] WLA[300] WLA[299] WLA[298] WLA[297] WLA[296] WLA[295] WLA[294] WLA[293] WLA[292]
+WLA[291] WLA[290] WLA[289] WLA[288] WLA[287] WLA[286] WLA[285] WLA[284] WLA[283] WLA[282]
+WLA[281] WLA[280] WLA[279] WLA[278] WLA[277] WLA[276] WLA[275] WLA[274] WLA[273] WLA[272]
+WLA[271] WLA[270] WLA[269] WLA[268] WLA[267] WLA[266] WLA[265] WLA[264] WLA[263] WLA[262]
+WLA[261] WLA[260] WLA[259] WLA[258] WLA[257] WLA[256] WLA[255] WLA[254] WLA[253] WLA[252]
+WLA[251] WLA[250] WLA[249] WLA[248] WLA[247] WLA[246] WLA[245] WLA[244] WLA[243] WLA[242]
+WLA[241] WLA[240] WLA[239] WLA[238] WLA[237] WLA[236] WLA[235] WLA[234] WLA[233] WLA[232]
+WLA[231] WLA[230] WLA[229] WLA[228] WLA[227] WLA[226] WLA[225] WLA[224] WLA[223] WLA[222]
+WLA[221] WLA[220] WLA[219] WLA[218] WLA[217] WLA[216] WLA[215] WLA[214] WLA[213] WLA[212]
+WLA[211] WLA[210] WLA[209] WLA[208] WLA[207] WLA[206] WLA[205] WLA[204] WLA[203] WLA[202]
+WLA[201] WLA[200] WLA[199] WLA[198] WLA[197] WLA[196] WLA[195] WLA[194] WLA[193] WLA[192]
+WLA[191] WLA[190] WLA[189] WLA[188] WLA[187] WLA[186] WLA[185] WLA[184] WLA[183] WLA[182]
+WLA[181] WLA[180] WLA[179] WLA[178] WLA[177] WLA[176] WLA[175] WLA[174] WLA[173] WLA[172]
+WLA[171] WLA[170] WLA[169] WLA[168] WLA[167] WLA[166] WLA[165] WLA[164] WLA[163] WLA[162]
+WLA[161] WLA[160] WLA[159] WLA[158] WLA[157] WLA[156] WLA[155] WLA[154] WLA[153] WLA[152]
+WLA[151] WLA[150] WLA[149] WLA[148] WLA[147] WLA[146] WLA[145] WLA[144] WLA[143] WLA[142]
+WLA[141] WLA[140] WLA[139] WLA[138] WLA[137] WLA[136] WLA[135] WLA[134] WLA[133] WLA[132]
+WLA[131] WLA[130] WLA[129] WLA[128] WLA[127] WLA[126] WLA[125] WLA[124] WLA[123] WLA[122]
+WLA[121] WLA[120] WLA[119] WLA[118] WLA[117] WLA[116] WLA[115] WLA[114] WLA[113] WLA[112]
+WLA[111] WLA[110] WLA[109] WLA[108] WLA[107] WLA[106] WLA[105] WLA[104] WLA[103] WLA[102]
+WLA[101] WLA[100] WLA[99] WLA[98] WLA[97] WLA[96] WLA[95] WLA[94] WLA[93] WLA[92]
+WLA[91] WLA[90] WLA[89] WLA[88] WLA[87] WLA[86] WLA[85] WLA[84] WLA[83] WLA[82]
+WLA[81] WLA[80] WLA[79] WLA[78] WLA[77] WLA[76] WLA[75] WLA[74] WLA[73] WLA[72]
+WLA[71] WLA[70] WLA[69] WLA[68] WLA[67] WLA[66] WLA[65] WLA[64] WLA[63] WLA[62]
+WLA[61] WLA[60] WLA[59] WLA[58] WLA[57] WLA[56] WLA[55] WLA[54] WLA[53] WLA[52]
+WLA[51] WLA[50] WLA[49] WLA[48] WLA[47] WLA[46] WLA[45] WLA[44] WLA[43] WLA[42]
+WLA[41] WLA[40] WLA[39] WLA[38] WLA[37] WLA[36] WLA[35] WLA[34] WLA[33] WLA[32]
+WLA[31] WLA[30] WLA[29] WLA[28] WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22]
+WLA[21] WLA[20] WLA[19] WLA[18] WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12]
+WLA[11] WLA[10] WLA[9] WLA[8] WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2]
+WLA[1] WLA[0] WLB[511] WLB[510] WLB[509] WLB[508] WLB[507] WLB[506] WLB[505] WLB[504]
+WLB[503] WLB[502] WLB[501] WLB[500] WLB[499] WLB[498] WLB[497] WLB[496] WLB[495] WLB[494]
+WLB[493] WLB[492] WLB[491] WLB[490] WLB[489] WLB[488] WLB[487] WLB[486] WLB[485] WLB[484]
+WLB[483] WLB[482] WLB[481] WLB[480] WLB[479] WLB[478] WLB[477] WLB[476] WLB[475] WLB[474]
+WLB[473] WLB[472] WLB[471] WLB[470] WLB[469] WLB[468] WLB[467] WLB[466] WLB[465] WLB[464]
+WLB[463] WLB[462] WLB[461] WLB[460] WLB[459] WLB[458] WLB[457] WLB[456] WLB[455] WLB[454]
+WLB[453] WLB[452] WLB[451] WLB[450] WLB[449] WLB[448] WLB[447] WLB[446] WLB[445] WLB[444]
+WLB[443] WLB[442] WLB[441] WLB[440] WLB[439] WLB[438] WLB[437] WLB[436] WLB[435] WLB[434]
+WLB[433] WLB[432] WLB[431] WLB[430] WLB[429] WLB[428] WLB[427] WLB[426] WLB[425] WLB[424]
+WLB[423] WLB[422] WLB[421] WLB[420] WLB[419] WLB[418] WLB[417] WLB[416] WLB[415] WLB[414]
+WLB[413] WLB[412] WLB[411] WLB[410] WLB[409] WLB[408] WLB[407] WLB[406] WLB[405] WLB[404]
+WLB[403] WLB[402] WLB[401] WLB[400] WLB[399] WLB[398] WLB[397] WLB[396] WLB[395] WLB[394]
+WLB[393] WLB[392] WLB[391] WLB[390] WLB[389] WLB[388] WLB[387] WLB[386] WLB[385] WLB[384]
+WLB[383] WLB[382] WLB[381] WLB[380] WLB[379] WLB[378] WLB[377] WLB[376] WLB[375] WLB[374]
+WLB[373] WLB[372] WLB[371] WLB[370] WLB[369] WLB[368] WLB[367] WLB[366] WLB[365] WLB[364]
+WLB[363] WLB[362] WLB[361] WLB[360] WLB[359] WLB[358] WLB[357] WLB[356] WLB[355] WLB[354]
+WLB[353] WLB[352] WLB[351] WLB[350] WLB[349] WLB[348] WLB[347] WLB[346] WLB[345] WLB[344]
+WLB[343] WLB[342] WLB[341] WLB[340] WLB[339] WLB[338] WLB[337] WLB[336] WLB[335] WLB[334]
+WLB[333] WLB[332] WLB[331] WLB[330] WLB[329] WLB[328] WLB[327] WLB[326] WLB[325] WLB[324]
+WLB[323] WLB[322] WLB[321] WLB[320] WLB[319] WLB[318] WLB[317] WLB[316] WLB[315] WLB[314]
+WLB[313] WLB[312] WLB[311] WLB[310] WLB[309] WLB[308] WLB[307] WLB[306] WLB[305] WLB[304]
+WLB[303] WLB[302] WLB[301] WLB[300] WLB[299] WLB[298] WLB[297] WLB[296] WLB[295] WLB[294]
+WLB[293] WLB[292] WLB[291] WLB[290] WLB[289] WLB[288] WLB[287] WLB[286] WLB[285] WLB[284]
+WLB[283] WLB[282] WLB[281] WLB[280] WLB[279] WLB[278] WLB[277] WLB[276] WLB[275] WLB[274]
+WLB[273] WLB[272] WLB[271] WLB[270] WLB[269] WLB[268] WLB[267] WLB[266] WLB[265] WLB[264]
+WLB[263] WLB[262] WLB[261] WLB[260] WLB[259] WLB[258] WLB[257] WLB[256] WLB[255] WLB[254]
+WLB[253] WLB[252] WLB[251] WLB[250] WLB[249] WLB[248] WLB[247] WLB[246] WLB[245] WLB[244]
+WLB[243] WLB[242] WLB[241] WLB[240] WLB[239] WLB[238] WLB[237] WLB[236] WLB[235] WLB[234]
+WLB[233] WLB[232] WLB[231] WLB[230] WLB[229] WLB[228] WLB[227] WLB[226] WLB[225] WLB[224]
+WLB[223] WLB[222] WLB[221] WLB[220] WLB[219] WLB[218] WLB[217] WLB[216] WLB[215] WLB[214]
+WLB[213] WLB[212] WLB[211] WLB[210] WLB[209] WLB[208] WLB[207] WLB[206] WLB[205] WLB[204]
+WLB[203] WLB[202] WLB[201] WLB[200] WLB[199] WLB[198] WLB[197] WLB[196] WLB[195] WLB[194]
+WLB[193] WLB[192] WLB[191] WLB[190] WLB[189] WLB[188] WLB[187] WLB[186] WLB[185] WLB[184]
+WLB[183] WLB[182] WLB[181] WLB[180] WLB[179] WLB[178] WLB[177] WLB[176] WLB[175] WLB[174]
+WLB[173] WLB[172] WLB[171] WLB[170] WLB[169] WLB[168] WLB[167] WLB[166] WLB[165] WLB[164]
+WLB[163] WLB[162] WLB[161] WLB[160] WLB[159] WLB[158] WLB[157] WLB[156] WLB[155] WLB[154]
+WLB[153] WLB[152] WLB[151] WLB[150] WLB[149] WLB[148] WLB[147] WLB[146] WLB[145] WLB[144]
+WLB[143] WLB[142] WLB[141] WLB[140] WLB[139] WLB[138] WLB[137] WLB[136] WLB[135] WLB[134]
+WLB[133] WLB[132] WLB[131] WLB[130] WLB[129] WLB[128] WLB[127] WLB[126] WLB[125] WLB[124]
+WLB[123] WLB[122] WLB[121] WLB[120] WLB[119] WLB[118] WLB[117] WLB[116] WLB[115] WLB[114]
+WLB[113] WLB[112] WLB[111] WLB[110] WLB[109] WLB[108] WLB[107] WLB[106] WLB[105] WLB[104]
+WLB[103] WLB[102] WLB[101] WLB[100] WLB[99] WLB[98] WLB[97] WLB[96] WLB[95] WLB[94]
+WLB[93] WLB[92] WLB[91] WLB[90] WLB[89] WLB[88] WLB[87] WLB[86] WLB[85] WLB[84]
+WLB[83] WLB[82] WLB[81] WLB[80] WLB[79] WLB[78] WLB[77] WLB[76] WLB[75] WLB[74]
+WLB[73] WLB[72] WLB[71] WLB[70] WLB[69] WLB[68] WLB[67] WLB[66] WLB[65] WLB[64]
+WLB[63] WLB[62] WLB[61] WLB[60] WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54]
+WLB[53] WLB[52] WLB[51] WLB[50] WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44]
+WLB[43] WLB[42] WLB[41] WLB[40] WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34]
+WLB[33] WLB[32] WLB[31] WLB[30] WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24]
+WLB[23] WLB[22] WLB[21] WLB[20] WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14]
+WLB[13] WLB[12] WLB[11] WLB[10] WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4]
+WLB[3] WLB[2] WLB[1] WLB[0] YXA[7] YXA[6] YXA[5] YXA[4] YXA[3] YXA[2]
+YXA[1] YXA[0] YXB[7] YXB[6] YXB[5] YXB[4] YXB[3] YXB[2] YXB[1] YXB[0] S55NLLGDPH_X512Y8D16_BW_Y512X8CELL_BW
XI21 BWENA[5] BWENB[5] CLKA CLKB CLKXA CLKXB DATAA[5] DATAB[5] DOUTA[5] DOUTB[5]
+STWLA VSS VSS VSS VSS VSS VSS VSS RWLA[0] RWLA[1]
+RWLB[0] RWLB[1] SACK1A SACK1B SACK4A SACK4B VDD VSS WEA WEB
+WLA[511] WLA[510] WLA[509] WLA[508] WLA[507] WLA[506] WLA[505] WLA[504] WLA[503] WLA[502]
+WLA[501] WLA[500] WLA[499] WLA[498] WLA[497] WLA[496] WLA[495] WLA[494] WLA[493] WLA[492]
+WLA[491] WLA[490] WLA[489] WLA[488] WLA[487] WLA[486] WLA[485] WLA[484] WLA[483] WLA[482]
+WLA[481] WLA[480] WLA[479] WLA[478] WLA[477] WLA[476] WLA[475] WLA[474] WLA[473] WLA[472]
+WLA[471] WLA[470] WLA[469] WLA[468] WLA[467] WLA[466] WLA[465] WLA[464] WLA[463] WLA[462]
+WLA[461] WLA[460] WLA[459] WLA[458] WLA[457] WLA[456] WLA[455] WLA[454] WLA[453] WLA[452]
+WLA[451] WLA[450] WLA[449] WLA[448] WLA[447] WLA[446] WLA[445] WLA[444] WLA[443] WLA[442]
+WLA[441] WLA[440] WLA[439] WLA[438] WLA[437] WLA[436] WLA[435] WLA[434] WLA[433] WLA[432]
+WLA[431] WLA[430] WLA[429] WLA[428] WLA[427] WLA[426] WLA[425] WLA[424] WLA[423] WLA[422]
+WLA[421] WLA[420] WLA[419] WLA[418] WLA[417] WLA[416] WLA[415] WLA[414] WLA[413] WLA[412]
+WLA[411] WLA[410] WLA[409] WLA[408] WLA[407] WLA[406] WLA[405] WLA[404] WLA[403] WLA[402]
+WLA[401] WLA[400] WLA[399] WLA[398] WLA[397] WLA[396] WLA[395] WLA[394] WLA[393] WLA[392]
+WLA[391] WLA[390] WLA[389] WLA[388] WLA[387] WLA[386] WLA[385] WLA[384] WLA[383] WLA[382]
+WLA[381] WLA[380] WLA[379] WLA[378] WLA[377] WLA[376] WLA[375] WLA[374] WLA[373] WLA[372]
+WLA[371] WLA[370] WLA[369] WLA[368] WLA[367] WLA[366] WLA[365] WLA[364] WLA[363] WLA[362]
+WLA[361] WLA[360] WLA[359] WLA[358] WLA[357] WLA[356] WLA[355] WLA[354] WLA[353] WLA[352]
+WLA[351] WLA[350] WLA[349] WLA[348] WLA[347] WLA[346] WLA[345] WLA[344] WLA[343] WLA[342]
+WLA[341] WLA[340] WLA[339] WLA[338] WLA[337] WLA[336] WLA[335] WLA[334] WLA[333] WLA[332]
+WLA[331] WLA[330] WLA[329] WLA[328] WLA[327] WLA[326] WLA[325] WLA[324] WLA[323] WLA[322]
+WLA[321] WLA[320] WLA[319] WLA[318] WLA[317] WLA[316] WLA[315] WLA[314] WLA[313] WLA[312]
+WLA[311] WLA[310] WLA[309] WLA[308] WLA[307] WLA[306] WLA[305] WLA[304] WLA[303] WLA[302]
+WLA[301] WLA[300] WLA[299] WLA[298] WLA[297] WLA[296] WLA[295] WLA[294] WLA[293] WLA[292]
+WLA[291] WLA[290] WLA[289] WLA[288] WLA[287] WLA[286] WLA[285] WLA[284] WLA[283] WLA[282]
+WLA[281] WLA[280] WLA[279] WLA[278] WLA[277] WLA[276] WLA[275] WLA[274] WLA[273] WLA[272]
+WLA[271] WLA[270] WLA[269] WLA[268] WLA[267] WLA[266] WLA[265] WLA[264] WLA[263] WLA[262]
+WLA[261] WLA[260] WLA[259] WLA[258] WLA[257] WLA[256] WLA[255] WLA[254] WLA[253] WLA[252]
+WLA[251] WLA[250] WLA[249] WLA[248] WLA[247] WLA[246] WLA[245] WLA[244] WLA[243] WLA[242]
+WLA[241] WLA[240] WLA[239] WLA[238] WLA[237] WLA[236] WLA[235] WLA[234] WLA[233] WLA[232]
+WLA[231] WLA[230] WLA[229] WLA[228] WLA[227] WLA[226] WLA[225] WLA[224] WLA[223] WLA[222]
+WLA[221] WLA[220] WLA[219] WLA[218] WLA[217] WLA[216] WLA[215] WLA[214] WLA[213] WLA[212]
+WLA[211] WLA[210] WLA[209] WLA[208] WLA[207] WLA[206] WLA[205] WLA[204] WLA[203] WLA[202]
+WLA[201] WLA[200] WLA[199] WLA[198] WLA[197] WLA[196] WLA[195] WLA[194] WLA[193] WLA[192]
+WLA[191] WLA[190] WLA[189] WLA[188] WLA[187] WLA[186] WLA[185] WLA[184] WLA[183] WLA[182]
+WLA[181] WLA[180] WLA[179] WLA[178] WLA[177] WLA[176] WLA[175] WLA[174] WLA[173] WLA[172]
+WLA[171] WLA[170] WLA[169] WLA[168] WLA[167] WLA[166] WLA[165] WLA[164] WLA[163] WLA[162]
+WLA[161] WLA[160] WLA[159] WLA[158] WLA[157] WLA[156] WLA[155] WLA[154] WLA[153] WLA[152]
+WLA[151] WLA[150] WLA[149] WLA[148] WLA[147] WLA[146] WLA[145] WLA[144] WLA[143] WLA[142]
+WLA[141] WLA[140] WLA[139] WLA[138] WLA[137] WLA[136] WLA[135] WLA[134] WLA[133] WLA[132]
+WLA[131] WLA[130] WLA[129] WLA[128] WLA[127] WLA[126] WLA[125] WLA[124] WLA[123] WLA[122]
+WLA[121] WLA[120] WLA[119] WLA[118] WLA[117] WLA[116] WLA[115] WLA[114] WLA[113] WLA[112]
+WLA[111] WLA[110] WLA[109] WLA[108] WLA[107] WLA[106] WLA[105] WLA[104] WLA[103] WLA[102]
+WLA[101] WLA[100] WLA[99] WLA[98] WLA[97] WLA[96] WLA[95] WLA[94] WLA[93] WLA[92]
+WLA[91] WLA[90] WLA[89] WLA[88] WLA[87] WLA[86] WLA[85] WLA[84] WLA[83] WLA[82]
+WLA[81] WLA[80] WLA[79] WLA[78] WLA[77] WLA[76] WLA[75] WLA[74] WLA[73] WLA[72]
+WLA[71] WLA[70] WLA[69] WLA[68] WLA[67] WLA[66] WLA[65] WLA[64] WLA[63] WLA[62]
+WLA[61] WLA[60] WLA[59] WLA[58] WLA[57] WLA[56] WLA[55] WLA[54] WLA[53] WLA[52]
+WLA[51] WLA[50] WLA[49] WLA[48] WLA[47] WLA[46] WLA[45] WLA[44] WLA[43] WLA[42]
+WLA[41] WLA[40] WLA[39] WLA[38] WLA[37] WLA[36] WLA[35] WLA[34] WLA[33] WLA[32]
+WLA[31] WLA[30] WLA[29] WLA[28] WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22]
+WLA[21] WLA[20] WLA[19] WLA[18] WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12]
+WLA[11] WLA[10] WLA[9] WLA[8] WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2]
+WLA[1] WLA[0] WLB[511] WLB[510] WLB[509] WLB[508] WLB[507] WLB[506] WLB[505] WLB[504]
+WLB[503] WLB[502] WLB[501] WLB[500] WLB[499] WLB[498] WLB[497] WLB[496] WLB[495] WLB[494]
+WLB[493] WLB[492] WLB[491] WLB[490] WLB[489] WLB[488] WLB[487] WLB[486] WLB[485] WLB[484]
+WLB[483] WLB[482] WLB[481] WLB[480] WLB[479] WLB[478] WLB[477] WLB[476] WLB[475] WLB[474]
+WLB[473] WLB[472] WLB[471] WLB[470] WLB[469] WLB[468] WLB[467] WLB[466] WLB[465] WLB[464]
+WLB[463] WLB[462] WLB[461] WLB[460] WLB[459] WLB[458] WLB[457] WLB[456] WLB[455] WLB[454]
+WLB[453] WLB[452] WLB[451] WLB[450] WLB[449] WLB[448] WLB[447] WLB[446] WLB[445] WLB[444]
+WLB[443] WLB[442] WLB[441] WLB[440] WLB[439] WLB[438] WLB[437] WLB[436] WLB[435] WLB[434]
+WLB[433] WLB[432] WLB[431] WLB[430] WLB[429] WLB[428] WLB[427] WLB[426] WLB[425] WLB[424]
+WLB[423] WLB[422] WLB[421] WLB[420] WLB[419] WLB[418] WLB[417] WLB[416] WLB[415] WLB[414]
+WLB[413] WLB[412] WLB[411] WLB[410] WLB[409] WLB[408] WLB[407] WLB[406] WLB[405] WLB[404]
+WLB[403] WLB[402] WLB[401] WLB[400] WLB[399] WLB[398] WLB[397] WLB[396] WLB[395] WLB[394]
+WLB[393] WLB[392] WLB[391] WLB[390] WLB[389] WLB[388] WLB[387] WLB[386] WLB[385] WLB[384]
+WLB[383] WLB[382] WLB[381] WLB[380] WLB[379] WLB[378] WLB[377] WLB[376] WLB[375] WLB[374]
+WLB[373] WLB[372] WLB[371] WLB[370] WLB[369] WLB[368] WLB[367] WLB[366] WLB[365] WLB[364]
+WLB[363] WLB[362] WLB[361] WLB[360] WLB[359] WLB[358] WLB[357] WLB[356] WLB[355] WLB[354]
+WLB[353] WLB[352] WLB[351] WLB[350] WLB[349] WLB[348] WLB[347] WLB[346] WLB[345] WLB[344]
+WLB[343] WLB[342] WLB[341] WLB[340] WLB[339] WLB[338] WLB[337] WLB[336] WLB[335] WLB[334]
+WLB[333] WLB[332] WLB[331] WLB[330] WLB[329] WLB[328] WLB[327] WLB[326] WLB[325] WLB[324]
+WLB[323] WLB[322] WLB[321] WLB[320] WLB[319] WLB[318] WLB[317] WLB[316] WLB[315] WLB[314]
+WLB[313] WLB[312] WLB[311] WLB[310] WLB[309] WLB[308] WLB[307] WLB[306] WLB[305] WLB[304]
+WLB[303] WLB[302] WLB[301] WLB[300] WLB[299] WLB[298] WLB[297] WLB[296] WLB[295] WLB[294]
+WLB[293] WLB[292] WLB[291] WLB[290] WLB[289] WLB[288] WLB[287] WLB[286] WLB[285] WLB[284]
+WLB[283] WLB[282] WLB[281] WLB[280] WLB[279] WLB[278] WLB[277] WLB[276] WLB[275] WLB[274]
+WLB[273] WLB[272] WLB[271] WLB[270] WLB[269] WLB[268] WLB[267] WLB[266] WLB[265] WLB[264]
+WLB[263] WLB[262] WLB[261] WLB[260] WLB[259] WLB[258] WLB[257] WLB[256] WLB[255] WLB[254]
+WLB[253] WLB[252] WLB[251] WLB[250] WLB[249] WLB[248] WLB[247] WLB[246] WLB[245] WLB[244]
+WLB[243] WLB[242] WLB[241] WLB[240] WLB[239] WLB[238] WLB[237] WLB[236] WLB[235] WLB[234]
+WLB[233] WLB[232] WLB[231] WLB[230] WLB[229] WLB[228] WLB[227] WLB[226] WLB[225] WLB[224]
+WLB[223] WLB[222] WLB[221] WLB[220] WLB[219] WLB[218] WLB[217] WLB[216] WLB[215] WLB[214]
+WLB[213] WLB[212] WLB[211] WLB[210] WLB[209] WLB[208] WLB[207] WLB[206] WLB[205] WLB[204]
+WLB[203] WLB[202] WLB[201] WLB[200] WLB[199] WLB[198] WLB[197] WLB[196] WLB[195] WLB[194]
+WLB[193] WLB[192] WLB[191] WLB[190] WLB[189] WLB[188] WLB[187] WLB[186] WLB[185] WLB[184]
+WLB[183] WLB[182] WLB[181] WLB[180] WLB[179] WLB[178] WLB[177] WLB[176] WLB[175] WLB[174]
+WLB[173] WLB[172] WLB[171] WLB[170] WLB[169] WLB[168] WLB[167] WLB[166] WLB[165] WLB[164]
+WLB[163] WLB[162] WLB[161] WLB[160] WLB[159] WLB[158] WLB[157] WLB[156] WLB[155] WLB[154]
+WLB[153] WLB[152] WLB[151] WLB[150] WLB[149] WLB[148] WLB[147] WLB[146] WLB[145] WLB[144]
+WLB[143] WLB[142] WLB[141] WLB[140] WLB[139] WLB[138] WLB[137] WLB[136] WLB[135] WLB[134]
+WLB[133] WLB[132] WLB[131] WLB[130] WLB[129] WLB[128] WLB[127] WLB[126] WLB[125] WLB[124]
+WLB[123] WLB[122] WLB[121] WLB[120] WLB[119] WLB[118] WLB[117] WLB[116] WLB[115] WLB[114]
+WLB[113] WLB[112] WLB[111] WLB[110] WLB[109] WLB[108] WLB[107] WLB[106] WLB[105] WLB[104]
+WLB[103] WLB[102] WLB[101] WLB[100] WLB[99] WLB[98] WLB[97] WLB[96] WLB[95] WLB[94]
+WLB[93] WLB[92] WLB[91] WLB[90] WLB[89] WLB[88] WLB[87] WLB[86] WLB[85] WLB[84]
+WLB[83] WLB[82] WLB[81] WLB[80] WLB[79] WLB[78] WLB[77] WLB[76] WLB[75] WLB[74]
+WLB[73] WLB[72] WLB[71] WLB[70] WLB[69] WLB[68] WLB[67] WLB[66] WLB[65] WLB[64]
+WLB[63] WLB[62] WLB[61] WLB[60] WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54]
+WLB[53] WLB[52] WLB[51] WLB[50] WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44]
+WLB[43] WLB[42] WLB[41] WLB[40] WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34]
+WLB[33] WLB[32] WLB[31] WLB[30] WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24]
+WLB[23] WLB[22] WLB[21] WLB[20] WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14]
+WLB[13] WLB[12] WLB[11] WLB[10] WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4]
+WLB[3] WLB[2] WLB[1] WLB[0] YXA[7] YXA[6] YXA[5] YXA[4] YXA[3] YXA[2]
+YXA[1] YXA[0] YXB[7] YXB[6] YXB[5] YXB[4] YXB[3] YXB[2] YXB[1] YXB[0] S55NLLGDPH_X512Y8D16_BW_Y512X8CELL_BW
XI22 BWENA[6] BWENB[6] CLKA CLKB CLKXA CLKXB DATAA[6] DATAB[6] DOUTA[6] DOUTB[6]
+STWLA VSS VSS VSS VSS VSS VSS VSS RWLA[0] RWLA[1]
+RWLB[0] RWLB[1] SACK1A SACK1B SACK4A SACK4B VDD VSS WEA WEB
+WLA[511] WLA[510] WLA[509] WLA[508] WLA[507] WLA[506] WLA[505] WLA[504] WLA[503] WLA[502]
+WLA[501] WLA[500] WLA[499] WLA[498] WLA[497] WLA[496] WLA[495] WLA[494] WLA[493] WLA[492]
+WLA[491] WLA[490] WLA[489] WLA[488] WLA[487] WLA[486] WLA[485] WLA[484] WLA[483] WLA[482]
+WLA[481] WLA[480] WLA[479] WLA[478] WLA[477] WLA[476] WLA[475] WLA[474] WLA[473] WLA[472]
+WLA[471] WLA[470] WLA[469] WLA[468] WLA[467] WLA[466] WLA[465] WLA[464] WLA[463] WLA[462]
+WLA[461] WLA[460] WLA[459] WLA[458] WLA[457] WLA[456] WLA[455] WLA[454] WLA[453] WLA[452]
+WLA[451] WLA[450] WLA[449] WLA[448] WLA[447] WLA[446] WLA[445] WLA[444] WLA[443] WLA[442]
+WLA[441] WLA[440] WLA[439] WLA[438] WLA[437] WLA[436] WLA[435] WLA[434] WLA[433] WLA[432]
+WLA[431] WLA[430] WLA[429] WLA[428] WLA[427] WLA[426] WLA[425] WLA[424] WLA[423] WLA[422]
+WLA[421] WLA[420] WLA[419] WLA[418] WLA[417] WLA[416] WLA[415] WLA[414] WLA[413] WLA[412]
+WLA[411] WLA[410] WLA[409] WLA[408] WLA[407] WLA[406] WLA[405] WLA[404] WLA[403] WLA[402]
+WLA[401] WLA[400] WLA[399] WLA[398] WLA[397] WLA[396] WLA[395] WLA[394] WLA[393] WLA[392]
+WLA[391] WLA[390] WLA[389] WLA[388] WLA[387] WLA[386] WLA[385] WLA[384] WLA[383] WLA[382]
+WLA[381] WLA[380] WLA[379] WLA[378] WLA[377] WLA[376] WLA[375] WLA[374] WLA[373] WLA[372]
+WLA[371] WLA[370] WLA[369] WLA[368] WLA[367] WLA[366] WLA[365] WLA[364] WLA[363] WLA[362]
+WLA[361] WLA[360] WLA[359] WLA[358] WLA[357] WLA[356] WLA[355] WLA[354] WLA[353] WLA[352]
+WLA[351] WLA[350] WLA[349] WLA[348] WLA[347] WLA[346] WLA[345] WLA[344] WLA[343] WLA[342]
+WLA[341] WLA[340] WLA[339] WLA[338] WLA[337] WLA[336] WLA[335] WLA[334] WLA[333] WLA[332]
+WLA[331] WLA[330] WLA[329] WLA[328] WLA[327] WLA[326] WLA[325] WLA[324] WLA[323] WLA[322]
+WLA[321] WLA[320] WLA[319] WLA[318] WLA[317] WLA[316] WLA[315] WLA[314] WLA[313] WLA[312]
+WLA[311] WLA[310] WLA[309] WLA[308] WLA[307] WLA[306] WLA[305] WLA[304] WLA[303] WLA[302]
+WLA[301] WLA[300] WLA[299] WLA[298] WLA[297] WLA[296] WLA[295] WLA[294] WLA[293] WLA[292]
+WLA[291] WLA[290] WLA[289] WLA[288] WLA[287] WLA[286] WLA[285] WLA[284] WLA[283] WLA[282]
+WLA[281] WLA[280] WLA[279] WLA[278] WLA[277] WLA[276] WLA[275] WLA[274] WLA[273] WLA[272]
+WLA[271] WLA[270] WLA[269] WLA[268] WLA[267] WLA[266] WLA[265] WLA[264] WLA[263] WLA[262]
+WLA[261] WLA[260] WLA[259] WLA[258] WLA[257] WLA[256] WLA[255] WLA[254] WLA[253] WLA[252]
+WLA[251] WLA[250] WLA[249] WLA[248] WLA[247] WLA[246] WLA[245] WLA[244] WLA[243] WLA[242]
+WLA[241] WLA[240] WLA[239] WLA[238] WLA[237] WLA[236] WLA[235] WLA[234] WLA[233] WLA[232]
+WLA[231] WLA[230] WLA[229] WLA[228] WLA[227] WLA[226] WLA[225] WLA[224] WLA[223] WLA[222]
+WLA[221] WLA[220] WLA[219] WLA[218] WLA[217] WLA[216] WLA[215] WLA[214] WLA[213] WLA[212]
+WLA[211] WLA[210] WLA[209] WLA[208] WLA[207] WLA[206] WLA[205] WLA[204] WLA[203] WLA[202]
+WLA[201] WLA[200] WLA[199] WLA[198] WLA[197] WLA[196] WLA[195] WLA[194] WLA[193] WLA[192]
+WLA[191] WLA[190] WLA[189] WLA[188] WLA[187] WLA[186] WLA[185] WLA[184] WLA[183] WLA[182]
+WLA[181] WLA[180] WLA[179] WLA[178] WLA[177] WLA[176] WLA[175] WLA[174] WLA[173] WLA[172]
+WLA[171] WLA[170] WLA[169] WLA[168] WLA[167] WLA[166] WLA[165] WLA[164] WLA[163] WLA[162]
+WLA[161] WLA[160] WLA[159] WLA[158] WLA[157] WLA[156] WLA[155] WLA[154] WLA[153] WLA[152]
+WLA[151] WLA[150] WLA[149] WLA[148] WLA[147] WLA[146] WLA[145] WLA[144] WLA[143] WLA[142]
+WLA[141] WLA[140] WLA[139] WLA[138] WLA[137] WLA[136] WLA[135] WLA[134] WLA[133] WLA[132]
+WLA[131] WLA[130] WLA[129] WLA[128] WLA[127] WLA[126] WLA[125] WLA[124] WLA[123] WLA[122]
+WLA[121] WLA[120] WLA[119] WLA[118] WLA[117] WLA[116] WLA[115] WLA[114] WLA[113] WLA[112]
+WLA[111] WLA[110] WLA[109] WLA[108] WLA[107] WLA[106] WLA[105] WLA[104] WLA[103] WLA[102]
+WLA[101] WLA[100] WLA[99] WLA[98] WLA[97] WLA[96] WLA[95] WLA[94] WLA[93] WLA[92]
+WLA[91] WLA[90] WLA[89] WLA[88] WLA[87] WLA[86] WLA[85] WLA[84] WLA[83] WLA[82]
+WLA[81] WLA[80] WLA[79] WLA[78] WLA[77] WLA[76] WLA[75] WLA[74] WLA[73] WLA[72]
+WLA[71] WLA[70] WLA[69] WLA[68] WLA[67] WLA[66] WLA[65] WLA[64] WLA[63] WLA[62]
+WLA[61] WLA[60] WLA[59] WLA[58] WLA[57] WLA[56] WLA[55] WLA[54] WLA[53] WLA[52]
+WLA[51] WLA[50] WLA[49] WLA[48] WLA[47] WLA[46] WLA[45] WLA[44] WLA[43] WLA[42]
+WLA[41] WLA[40] WLA[39] WLA[38] WLA[37] WLA[36] WLA[35] WLA[34] WLA[33] WLA[32]
+WLA[31] WLA[30] WLA[29] WLA[28] WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22]
+WLA[21] WLA[20] WLA[19] WLA[18] WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12]
+WLA[11] WLA[10] WLA[9] WLA[8] WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2]
+WLA[1] WLA[0] WLB[511] WLB[510] WLB[509] WLB[508] WLB[507] WLB[506] WLB[505] WLB[504]
+WLB[503] WLB[502] WLB[501] WLB[500] WLB[499] WLB[498] WLB[497] WLB[496] WLB[495] WLB[494]
+WLB[493] WLB[492] WLB[491] WLB[490] WLB[489] WLB[488] WLB[487] WLB[486] WLB[485] WLB[484]
+WLB[483] WLB[482] WLB[481] WLB[480] WLB[479] WLB[478] WLB[477] WLB[476] WLB[475] WLB[474]
+WLB[473] WLB[472] WLB[471] WLB[470] WLB[469] WLB[468] WLB[467] WLB[466] WLB[465] WLB[464]
+WLB[463] WLB[462] WLB[461] WLB[460] WLB[459] WLB[458] WLB[457] WLB[456] WLB[455] WLB[454]
+WLB[453] WLB[452] WLB[451] WLB[450] WLB[449] WLB[448] WLB[447] WLB[446] WLB[445] WLB[444]
+WLB[443] WLB[442] WLB[441] WLB[440] WLB[439] WLB[438] WLB[437] WLB[436] WLB[435] WLB[434]
+WLB[433] WLB[432] WLB[431] WLB[430] WLB[429] WLB[428] WLB[427] WLB[426] WLB[425] WLB[424]
+WLB[423] WLB[422] WLB[421] WLB[420] WLB[419] WLB[418] WLB[417] WLB[416] WLB[415] WLB[414]
+WLB[413] WLB[412] WLB[411] WLB[410] WLB[409] WLB[408] WLB[407] WLB[406] WLB[405] WLB[404]
+WLB[403] WLB[402] WLB[401] WLB[400] WLB[399] WLB[398] WLB[397] WLB[396] WLB[395] WLB[394]
+WLB[393] WLB[392] WLB[391] WLB[390] WLB[389] WLB[388] WLB[387] WLB[386] WLB[385] WLB[384]
+WLB[383] WLB[382] WLB[381] WLB[380] WLB[379] WLB[378] WLB[377] WLB[376] WLB[375] WLB[374]
+WLB[373] WLB[372] WLB[371] WLB[370] WLB[369] WLB[368] WLB[367] WLB[366] WLB[365] WLB[364]
+WLB[363] WLB[362] WLB[361] WLB[360] WLB[359] WLB[358] WLB[357] WLB[356] WLB[355] WLB[354]
+WLB[353] WLB[352] WLB[351] WLB[350] WLB[349] WLB[348] WLB[347] WLB[346] WLB[345] WLB[344]
+WLB[343] WLB[342] WLB[341] WLB[340] WLB[339] WLB[338] WLB[337] WLB[336] WLB[335] WLB[334]
+WLB[333] WLB[332] WLB[331] WLB[330] WLB[329] WLB[328] WLB[327] WLB[326] WLB[325] WLB[324]
+WLB[323] WLB[322] WLB[321] WLB[320] WLB[319] WLB[318] WLB[317] WLB[316] WLB[315] WLB[314]
+WLB[313] WLB[312] WLB[311] WLB[310] WLB[309] WLB[308] WLB[307] WLB[306] WLB[305] WLB[304]
+WLB[303] WLB[302] WLB[301] WLB[300] WLB[299] WLB[298] WLB[297] WLB[296] WLB[295] WLB[294]
+WLB[293] WLB[292] WLB[291] WLB[290] WLB[289] WLB[288] WLB[287] WLB[286] WLB[285] WLB[284]
+WLB[283] WLB[282] WLB[281] WLB[280] WLB[279] WLB[278] WLB[277] WLB[276] WLB[275] WLB[274]
+WLB[273] WLB[272] WLB[271] WLB[270] WLB[269] WLB[268] WLB[267] WLB[266] WLB[265] WLB[264]
+WLB[263] WLB[262] WLB[261] WLB[260] WLB[259] WLB[258] WLB[257] WLB[256] WLB[255] WLB[254]
+WLB[253] WLB[252] WLB[251] WLB[250] WLB[249] WLB[248] WLB[247] WLB[246] WLB[245] WLB[244]
+WLB[243] WLB[242] WLB[241] WLB[240] WLB[239] WLB[238] WLB[237] WLB[236] WLB[235] WLB[234]
+WLB[233] WLB[232] WLB[231] WLB[230] WLB[229] WLB[228] WLB[227] WLB[226] WLB[225] WLB[224]
+WLB[223] WLB[222] WLB[221] WLB[220] WLB[219] WLB[218] WLB[217] WLB[216] WLB[215] WLB[214]
+WLB[213] WLB[212] WLB[211] WLB[210] WLB[209] WLB[208] WLB[207] WLB[206] WLB[205] WLB[204]
+WLB[203] WLB[202] WLB[201] WLB[200] WLB[199] WLB[198] WLB[197] WLB[196] WLB[195] WLB[194]
+WLB[193] WLB[192] WLB[191] WLB[190] WLB[189] WLB[188] WLB[187] WLB[186] WLB[185] WLB[184]
+WLB[183] WLB[182] WLB[181] WLB[180] WLB[179] WLB[178] WLB[177] WLB[176] WLB[175] WLB[174]
+WLB[173] WLB[172] WLB[171] WLB[170] WLB[169] WLB[168] WLB[167] WLB[166] WLB[165] WLB[164]
+WLB[163] WLB[162] WLB[161] WLB[160] WLB[159] WLB[158] WLB[157] WLB[156] WLB[155] WLB[154]
+WLB[153] WLB[152] WLB[151] WLB[150] WLB[149] WLB[148] WLB[147] WLB[146] WLB[145] WLB[144]
+WLB[143] WLB[142] WLB[141] WLB[140] WLB[139] WLB[138] WLB[137] WLB[136] WLB[135] WLB[134]
+WLB[133] WLB[132] WLB[131] WLB[130] WLB[129] WLB[128] WLB[127] WLB[126] WLB[125] WLB[124]
+WLB[123] WLB[122] WLB[121] WLB[120] WLB[119] WLB[118] WLB[117] WLB[116] WLB[115] WLB[114]
+WLB[113] WLB[112] WLB[111] WLB[110] WLB[109] WLB[108] WLB[107] WLB[106] WLB[105] WLB[104]
+WLB[103] WLB[102] WLB[101] WLB[100] WLB[99] WLB[98] WLB[97] WLB[96] WLB[95] WLB[94]
+WLB[93] WLB[92] WLB[91] WLB[90] WLB[89] WLB[88] WLB[87] WLB[86] WLB[85] WLB[84]
+WLB[83] WLB[82] WLB[81] WLB[80] WLB[79] WLB[78] WLB[77] WLB[76] WLB[75] WLB[74]
+WLB[73] WLB[72] WLB[71] WLB[70] WLB[69] WLB[68] WLB[67] WLB[66] WLB[65] WLB[64]
+WLB[63] WLB[62] WLB[61] WLB[60] WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54]
+WLB[53] WLB[52] WLB[51] WLB[50] WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44]
+WLB[43] WLB[42] WLB[41] WLB[40] WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34]
+WLB[33] WLB[32] WLB[31] WLB[30] WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24]
+WLB[23] WLB[22] WLB[21] WLB[20] WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14]
+WLB[13] WLB[12] WLB[11] WLB[10] WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4]
+WLB[3] WLB[2] WLB[1] WLB[0] YXA[7] YXA[6] YXA[5] YXA[4] YXA[3] YXA[2]
+YXA[1] YXA[0] YXB[7] YXB[6] YXB[5] YXB[4] YXB[3] YXB[2] YXB[1] YXB[0] S55NLLGDPH_X512Y8D16_BW_Y512X8CELL_BW
XI23 BWENA[7] BWENB[7] CLKA CLKB CLKXA CLKXB DATAA[7] DATAB[7] DOUTA[7] DOUTB[7]
+STWLA VSS VSS VSS VSS VSS VSS VSS RWLA[0] RWLA[1]
+RWLB[0] RWLB[1] SACK1A SACK1B SACK4A SACK4B VDD VSS WEA WEB
+WLA[511] WLA[510] WLA[509] WLA[508] WLA[507] WLA[506] WLA[505] WLA[504] WLA[503] WLA[502]
+WLA[501] WLA[500] WLA[499] WLA[498] WLA[497] WLA[496] WLA[495] WLA[494] WLA[493] WLA[492]
+WLA[491] WLA[490] WLA[489] WLA[488] WLA[487] WLA[486] WLA[485] WLA[484] WLA[483] WLA[482]
+WLA[481] WLA[480] WLA[479] WLA[478] WLA[477] WLA[476] WLA[475] WLA[474] WLA[473] WLA[472]
+WLA[471] WLA[470] WLA[469] WLA[468] WLA[467] WLA[466] WLA[465] WLA[464] WLA[463] WLA[462]
+WLA[461] WLA[460] WLA[459] WLA[458] WLA[457] WLA[456] WLA[455] WLA[454] WLA[453] WLA[452]
+WLA[451] WLA[450] WLA[449] WLA[448] WLA[447] WLA[446] WLA[445] WLA[444] WLA[443] WLA[442]
+WLA[441] WLA[440] WLA[439] WLA[438] WLA[437] WLA[436] WLA[435] WLA[434] WLA[433] WLA[432]
+WLA[431] WLA[430] WLA[429] WLA[428] WLA[427] WLA[426] WLA[425] WLA[424] WLA[423] WLA[422]
+WLA[421] WLA[420] WLA[419] WLA[418] WLA[417] WLA[416] WLA[415] WLA[414] WLA[413] WLA[412]
+WLA[411] WLA[410] WLA[409] WLA[408] WLA[407] WLA[406] WLA[405] WLA[404] WLA[403] WLA[402]
+WLA[401] WLA[400] WLA[399] WLA[398] WLA[397] WLA[396] WLA[395] WLA[394] WLA[393] WLA[392]
+WLA[391] WLA[390] WLA[389] WLA[388] WLA[387] WLA[386] WLA[385] WLA[384] WLA[383] WLA[382]
+WLA[381] WLA[380] WLA[379] WLA[378] WLA[377] WLA[376] WLA[375] WLA[374] WLA[373] WLA[372]
+WLA[371] WLA[370] WLA[369] WLA[368] WLA[367] WLA[366] WLA[365] WLA[364] WLA[363] WLA[362]
+WLA[361] WLA[360] WLA[359] WLA[358] WLA[357] WLA[356] WLA[355] WLA[354] WLA[353] WLA[352]
+WLA[351] WLA[350] WLA[349] WLA[348] WLA[347] WLA[346] WLA[345] WLA[344] WLA[343] WLA[342]
+WLA[341] WLA[340] WLA[339] WLA[338] WLA[337] WLA[336] WLA[335] WLA[334] WLA[333] WLA[332]
+WLA[331] WLA[330] WLA[329] WLA[328] WLA[327] WLA[326] WLA[325] WLA[324] WLA[323] WLA[322]
+WLA[321] WLA[320] WLA[319] WLA[318] WLA[317] WLA[316] WLA[315] WLA[314] WLA[313] WLA[312]
+WLA[311] WLA[310] WLA[309] WLA[308] WLA[307] WLA[306] WLA[305] WLA[304] WLA[303] WLA[302]
+WLA[301] WLA[300] WLA[299] WLA[298] WLA[297] WLA[296] WLA[295] WLA[294] WLA[293] WLA[292]
+WLA[291] WLA[290] WLA[289] WLA[288] WLA[287] WLA[286] WLA[285] WLA[284] WLA[283] WLA[282]
+WLA[281] WLA[280] WLA[279] WLA[278] WLA[277] WLA[276] WLA[275] WLA[274] WLA[273] WLA[272]
+WLA[271] WLA[270] WLA[269] WLA[268] WLA[267] WLA[266] WLA[265] WLA[264] WLA[263] WLA[262]
+WLA[261] WLA[260] WLA[259] WLA[258] WLA[257] WLA[256] WLA[255] WLA[254] WLA[253] WLA[252]
+WLA[251] WLA[250] WLA[249] WLA[248] WLA[247] WLA[246] WLA[245] WLA[244] WLA[243] WLA[242]
+WLA[241] WLA[240] WLA[239] WLA[238] WLA[237] WLA[236] WLA[235] WLA[234] WLA[233] WLA[232]
+WLA[231] WLA[230] WLA[229] WLA[228] WLA[227] WLA[226] WLA[225] WLA[224] WLA[223] WLA[222]
+WLA[221] WLA[220] WLA[219] WLA[218] WLA[217] WLA[216] WLA[215] WLA[214] WLA[213] WLA[212]
+WLA[211] WLA[210] WLA[209] WLA[208] WLA[207] WLA[206] WLA[205] WLA[204] WLA[203] WLA[202]
+WLA[201] WLA[200] WLA[199] WLA[198] WLA[197] WLA[196] WLA[195] WLA[194] WLA[193] WLA[192]
+WLA[191] WLA[190] WLA[189] WLA[188] WLA[187] WLA[186] WLA[185] WLA[184] WLA[183] WLA[182]
+WLA[181] WLA[180] WLA[179] WLA[178] WLA[177] WLA[176] WLA[175] WLA[174] WLA[173] WLA[172]
+WLA[171] WLA[170] WLA[169] WLA[168] WLA[167] WLA[166] WLA[165] WLA[164] WLA[163] WLA[162]
+WLA[161] WLA[160] WLA[159] WLA[158] WLA[157] WLA[156] WLA[155] WLA[154] WLA[153] WLA[152]
+WLA[151] WLA[150] WLA[149] WLA[148] WLA[147] WLA[146] WLA[145] WLA[144] WLA[143] WLA[142]
+WLA[141] WLA[140] WLA[139] WLA[138] WLA[137] WLA[136] WLA[135] WLA[134] WLA[133] WLA[132]
+WLA[131] WLA[130] WLA[129] WLA[128] WLA[127] WLA[126] WLA[125] WLA[124] WLA[123] WLA[122]
+WLA[121] WLA[120] WLA[119] WLA[118] WLA[117] WLA[116] WLA[115] WLA[114] WLA[113] WLA[112]
+WLA[111] WLA[110] WLA[109] WLA[108] WLA[107] WLA[106] WLA[105] WLA[104] WLA[103] WLA[102]
+WLA[101] WLA[100] WLA[99] WLA[98] WLA[97] WLA[96] WLA[95] WLA[94] WLA[93] WLA[92]
+WLA[91] WLA[90] WLA[89] WLA[88] WLA[87] WLA[86] WLA[85] WLA[84] WLA[83] WLA[82]
+WLA[81] WLA[80] WLA[79] WLA[78] WLA[77] WLA[76] WLA[75] WLA[74] WLA[73] WLA[72]
+WLA[71] WLA[70] WLA[69] WLA[68] WLA[67] WLA[66] WLA[65] WLA[64] WLA[63] WLA[62]
+WLA[61] WLA[60] WLA[59] WLA[58] WLA[57] WLA[56] WLA[55] WLA[54] WLA[53] WLA[52]
+WLA[51] WLA[50] WLA[49] WLA[48] WLA[47] WLA[46] WLA[45] WLA[44] WLA[43] WLA[42]
+WLA[41] WLA[40] WLA[39] WLA[38] WLA[37] WLA[36] WLA[35] WLA[34] WLA[33] WLA[32]
+WLA[31] WLA[30] WLA[29] WLA[28] WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22]
+WLA[21] WLA[20] WLA[19] WLA[18] WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12]
+WLA[11] WLA[10] WLA[9] WLA[8] WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2]
+WLA[1] WLA[0] WLB[511] WLB[510] WLB[509] WLB[508] WLB[507] WLB[506] WLB[505] WLB[504]
+WLB[503] WLB[502] WLB[501] WLB[500] WLB[499] WLB[498] WLB[497] WLB[496] WLB[495] WLB[494]
+WLB[493] WLB[492] WLB[491] WLB[490] WLB[489] WLB[488] WLB[487] WLB[486] WLB[485] WLB[484]
+WLB[483] WLB[482] WLB[481] WLB[480] WLB[479] WLB[478] WLB[477] WLB[476] WLB[475] WLB[474]
+WLB[473] WLB[472] WLB[471] WLB[470] WLB[469] WLB[468] WLB[467] WLB[466] WLB[465] WLB[464]
+WLB[463] WLB[462] WLB[461] WLB[460] WLB[459] WLB[458] WLB[457] WLB[456] WLB[455] WLB[454]
+WLB[453] WLB[452] WLB[451] WLB[450] WLB[449] WLB[448] WLB[447] WLB[446] WLB[445] WLB[444]
+WLB[443] WLB[442] WLB[441] WLB[440] WLB[439] WLB[438] WLB[437] WLB[436] WLB[435] WLB[434]
+WLB[433] WLB[432] WLB[431] WLB[430] WLB[429] WLB[428] WLB[427] WLB[426] WLB[425] WLB[424]
+WLB[423] WLB[422] WLB[421] WLB[420] WLB[419] WLB[418] WLB[417] WLB[416] WLB[415] WLB[414]
+WLB[413] WLB[412] WLB[411] WLB[410] WLB[409] WLB[408] WLB[407] WLB[406] WLB[405] WLB[404]
+WLB[403] WLB[402] WLB[401] WLB[400] WLB[399] WLB[398] WLB[397] WLB[396] WLB[395] WLB[394]
+WLB[393] WLB[392] WLB[391] WLB[390] WLB[389] WLB[388] WLB[387] WLB[386] WLB[385] WLB[384]
+WLB[383] WLB[382] WLB[381] WLB[380] WLB[379] WLB[378] WLB[377] WLB[376] WLB[375] WLB[374]
+WLB[373] WLB[372] WLB[371] WLB[370] WLB[369] WLB[368] WLB[367] WLB[366] WLB[365] WLB[364]
+WLB[363] WLB[362] WLB[361] WLB[360] WLB[359] WLB[358] WLB[357] WLB[356] WLB[355] WLB[354]
+WLB[353] WLB[352] WLB[351] WLB[350] WLB[349] WLB[348] WLB[347] WLB[346] WLB[345] WLB[344]
+WLB[343] WLB[342] WLB[341] WLB[340] WLB[339] WLB[338] WLB[337] WLB[336] WLB[335] WLB[334]
+WLB[333] WLB[332] WLB[331] WLB[330] WLB[329] WLB[328] WLB[327] WLB[326] WLB[325] WLB[324]
+WLB[323] WLB[322] WLB[321] WLB[320] WLB[319] WLB[318] WLB[317] WLB[316] WLB[315] WLB[314]
+WLB[313] WLB[312] WLB[311] WLB[310] WLB[309] WLB[308] WLB[307] WLB[306] WLB[305] WLB[304]
+WLB[303] WLB[302] WLB[301] WLB[300] WLB[299] WLB[298] WLB[297] WLB[296] WLB[295] WLB[294]
+WLB[293] WLB[292] WLB[291] WLB[290] WLB[289] WLB[288] WLB[287] WLB[286] WLB[285] WLB[284]
+WLB[283] WLB[282] WLB[281] WLB[280] WLB[279] WLB[278] WLB[277] WLB[276] WLB[275] WLB[274]
+WLB[273] WLB[272] WLB[271] WLB[270] WLB[269] WLB[268] WLB[267] WLB[266] WLB[265] WLB[264]
+WLB[263] WLB[262] WLB[261] WLB[260] WLB[259] WLB[258] WLB[257] WLB[256] WLB[255] WLB[254]
+WLB[253] WLB[252] WLB[251] WLB[250] WLB[249] WLB[248] WLB[247] WLB[246] WLB[245] WLB[244]
+WLB[243] WLB[242] WLB[241] WLB[240] WLB[239] WLB[238] WLB[237] WLB[236] WLB[235] WLB[234]
+WLB[233] WLB[232] WLB[231] WLB[230] WLB[229] WLB[228] WLB[227] WLB[226] WLB[225] WLB[224]
+WLB[223] WLB[222] WLB[221] WLB[220] WLB[219] WLB[218] WLB[217] WLB[216] WLB[215] WLB[214]
+WLB[213] WLB[212] WLB[211] WLB[210] WLB[209] WLB[208] WLB[207] WLB[206] WLB[205] WLB[204]
+WLB[203] WLB[202] WLB[201] WLB[200] WLB[199] WLB[198] WLB[197] WLB[196] WLB[195] WLB[194]
+WLB[193] WLB[192] WLB[191] WLB[190] WLB[189] WLB[188] WLB[187] WLB[186] WLB[185] WLB[184]
+WLB[183] WLB[182] WLB[181] WLB[180] WLB[179] WLB[178] WLB[177] WLB[176] WLB[175] WLB[174]
+WLB[173] WLB[172] WLB[171] WLB[170] WLB[169] WLB[168] WLB[167] WLB[166] WLB[165] WLB[164]
+WLB[163] WLB[162] WLB[161] WLB[160] WLB[159] WLB[158] WLB[157] WLB[156] WLB[155] WLB[154]
+WLB[153] WLB[152] WLB[151] WLB[150] WLB[149] WLB[148] WLB[147] WLB[146] WLB[145] WLB[144]
+WLB[143] WLB[142] WLB[141] WLB[140] WLB[139] WLB[138] WLB[137] WLB[136] WLB[135] WLB[134]
+WLB[133] WLB[132] WLB[131] WLB[130] WLB[129] WLB[128] WLB[127] WLB[126] WLB[125] WLB[124]
+WLB[123] WLB[122] WLB[121] WLB[120] WLB[119] WLB[118] WLB[117] WLB[116] WLB[115] WLB[114]
+WLB[113] WLB[112] WLB[111] WLB[110] WLB[109] WLB[108] WLB[107] WLB[106] WLB[105] WLB[104]
+WLB[103] WLB[102] WLB[101] WLB[100] WLB[99] WLB[98] WLB[97] WLB[96] WLB[95] WLB[94]
+WLB[93] WLB[92] WLB[91] WLB[90] WLB[89] WLB[88] WLB[87] WLB[86] WLB[85] WLB[84]
+WLB[83] WLB[82] WLB[81] WLB[80] WLB[79] WLB[78] WLB[77] WLB[76] WLB[75] WLB[74]
+WLB[73] WLB[72] WLB[71] WLB[70] WLB[69] WLB[68] WLB[67] WLB[66] WLB[65] WLB[64]
+WLB[63] WLB[62] WLB[61] WLB[60] WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54]
+WLB[53] WLB[52] WLB[51] WLB[50] WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44]
+WLB[43] WLB[42] WLB[41] WLB[40] WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34]
+WLB[33] WLB[32] WLB[31] WLB[30] WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24]
+WLB[23] WLB[22] WLB[21] WLB[20] WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14]
+WLB[13] WLB[12] WLB[11] WLB[10] WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4]
+WLB[3] WLB[2] WLB[1] WLB[0] YXA[7] YXA[6] YXA[5] YXA[4] YXA[3] YXA[2]
+YXA[1] YXA[0] YXB[7] YXB[6] YXB[5] YXB[4] YXB[3] YXB[2] YXB[1] YXB[0] S55NLLGDPH_X512Y8D16_BW_Y512X8CELL_BW
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    S55NLLGDPH_X512Y8D16_BW_XDEC
* View Name:    schematic
************************************************************************

.SUBCKT S55NLLGDPH_X512Y8D16_BW_XDEC FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA PXB
+PXC VDD VSS WL[7] WL[6] WL[5] WL[4] WL[3] WL[2] WL[1]
+WL[0]
M0 VSS 52 50 VSS N12LL L=6E-08 W=1E-06
M1 50 52 VSS VSS N12LL L=6E-08 W=1E-06
M2 VSS 52 50 VSS N12LL L=6E-08 W=1E-06
M3 52 49 VSS VSS N12LL L=6E-08 W=1E-06
M4 VSS 49 52 VSS N12LL L=6E-08 W=1E-06
M5 52 49 VSS VSS N12LL L=6E-08 W=1E-06
M6 85 PXA 49 VSS N12LL L=6E-08 W=8E-07
M7 86 PXB 85 VSS N12LL L=6E-08 W=8E-07
M8 VSS PXC 86 VSS N12LL L=6E-08 W=8E-07
M9 54 52 FCKX[1] VSS N12LL L=6E-08 W=8E-07
M10 58 52 FCKX[3] VSS N12LL L=6E-08 W=8E-07
M11 59 52 FCKX[5] VSS N12LL L=6E-08 W=8E-07
M12 FCKX[7] 52 55 VSS N12LL L=6E-08 W=8E-07
M13 53 52 FCKX[0] VSS N12LL L=6E-08 W=8E-07
M14 56 52 FCKX[2] VSS N12LL L=6E-08 W=8E-07
M15 57 52 FCKX[4] VSS N12LL L=6E-08 W=8E-07
M16 60 52 FCKX[6] VSS N12LL L=6E-08 W=8E-07
M17 61 53 VSS VSS N12LL L=6E-08 W=3.5E-07
M18 VSS 53 61 VSS N12LL L=6E-08 W=3.5E-07
M19 62 54 VSS VSS N12LL L=6E-08 W=3.5E-07
M20 VSS 54 62 VSS N12LL L=6E-08 W=3.5E-07
M21 63 56 VSS VSS N12LL L=6E-08 W=3.5E-07
M22 VSS 56 63 VSS N12LL L=6E-08 W=3.5E-07
M23 64 58 VSS VSS N12LL L=6E-08 W=3.5E-07
M24 VSS 58 64 VSS N12LL L=6E-08 W=3.5E-07
M25 65 57 VSS VSS N12LL L=6E-08 W=3.5E-07
M26 VSS 57 65 VSS N12LL L=6E-08 W=3.5E-07
M27 66 59 VSS VSS N12LL L=6E-08 W=3.5E-07
M28 VSS 59 66 VSS N12LL L=6E-08 W=3.5E-07
M29 67 60 VSS VSS N12LL L=6E-08 W=3.5E-07
M30 VSS 60 67 VSS N12LL L=6E-08 W=3.5E-07
M31 68 55 VSS VSS N12LL L=6E-08 W=3.5E-07
M32 VSS 55 68 VSS N12LL L=6E-08 W=3.5E-07
M33 69 61 VSS VSS N12LL L=6E-08 W=1.5E-06
M34 VSS 61 69 VSS N12LL L=6E-08 W=1.5E-06
M35 70 62 VSS VSS N12LL L=6E-08 W=1.5E-06
M36 VSS 62 70 VSS N12LL L=6E-08 W=1.5E-06
M37 71 63 VSS VSS N12LL L=6E-08 W=1.5E-06
M38 VSS 63 71 VSS N12LL L=6E-08 W=1.5E-06
M39 72 64 VSS VSS N12LL L=6E-08 W=1.5E-06
M40 VSS 64 72 VSS N12LL L=6E-08 W=1.5E-06
M41 73 65 VSS VSS N12LL L=6E-08 W=1.5E-06
M42 VSS 65 73 VSS N12LL L=6E-08 W=1.5E-06
M43 74 66 VSS VSS N12LL L=6E-08 W=1.5E-06
M44 VSS 66 74 VSS N12LL L=6E-08 W=1.5E-06
M45 75 67 VSS VSS N12LL L=6E-08 W=1.5E-06
M46 VSS 67 75 VSS N12LL L=6E-08 W=1.5E-06
M47 76 68 VSS VSS N12LL L=6E-08 W=1.5E-06
M48 VSS 68 76 VSS N12LL L=6E-08 W=1.5E-06
M49 WL[0] 69 VSS VSS N12LL L=6E-08 W=2E-06
M50 VSS 69 WL[0] VSS N12LL L=6E-08 W=2E-06
M51 WL[1] 70 VSS VSS N12LL L=6E-08 W=2E-06
M52 VSS 70 WL[1] VSS N12LL L=6E-08 W=2E-06
M53 WL[2] 71 VSS VSS N12LL L=6E-08 W=2E-06
M54 VSS 71 WL[2] VSS N12LL L=6E-08 W=2E-06
M55 WL[3] 72 VSS VSS N12LL L=6E-08 W=2E-06
M56 VSS 72 WL[3] VSS N12LL L=6E-08 W=2E-06
M57 WL[4] 73 VSS VSS N12LL L=6E-08 W=2E-06
M58 VSS 73 WL[4] VSS N12LL L=6E-08 W=2E-06
M59 WL[5] 74 VSS VSS N12LL L=6E-08 W=2E-06
M60 VSS 74 WL[5] VSS N12LL L=6E-08 W=2E-06
M61 WL[6] 75 VSS VSS N12LL L=6E-08 W=2E-06
M62 VSS 75 WL[6] VSS N12LL L=6E-08 W=2E-06
M63 WL[7] 76 VSS VSS N12LL L=6E-08 W=2E-06
M64 VSS 76 WL[7] VSS N12LL L=6E-08 W=2E-06
M65 WL[0] 69 VDD VDD PHVT12LL L=6E-08 W=2.5E-06
M66 VDD 69 WL[0] VDD PHVT12LL L=6E-08 W=2.5E-06
M67 WL[1] 70 VDD VDD PHVT12LL L=6E-08 W=2.5E-06
M68 VDD 70 WL[1] VDD PHVT12LL L=6E-08 W=2.5E-06
M69 WL[2] 71 VDD VDD PHVT12LL L=6E-08 W=2.5E-06
M70 VDD 71 WL[2] VDD PHVT12LL L=6E-08 W=2.5E-06
M71 WL[3] 72 VDD VDD PHVT12LL L=6E-08 W=2.5E-06
M72 VDD 72 WL[3] VDD PHVT12LL L=6E-08 W=2.5E-06
M73 WL[4] 73 VDD VDD PHVT12LL L=6E-08 W=2.5E-06
M74 VDD 73 WL[4] VDD PHVT12LL L=6E-08 W=2.5E-06
M75 WL[5] 74 VDD VDD PHVT12LL L=6E-08 W=2.5E-06
M76 VDD 74 WL[5] VDD PHVT12LL L=6E-08 W=2.5E-06
M77 WL[6] 75 VDD VDD PHVT12LL L=6E-08 W=2.5E-06
M78 VDD 75 WL[6] VDD PHVT12LL L=6E-08 W=2.5E-06
M79 WL[7] 76 VDD VDD PHVT12LL L=6E-08 W=2.5E-06
M80 VDD 76 WL[7] VDD PHVT12LL L=6E-08 W=2.5E-06
M81 WL[0] 69 VDD VDD PHVT12LL L=6E-08 W=2.5E-06
M82 VDD 69 WL[0] VDD PHVT12LL L=6E-08 W=2.5E-06
M83 WL[1] 70 VDD VDD PHVT12LL L=6E-08 W=2.5E-06
M84 VDD 70 WL[1] VDD PHVT12LL L=6E-08 W=2.5E-06
M85 WL[2] 71 VDD VDD PHVT12LL L=6E-08 W=2.5E-06
M86 VDD 71 WL[2] VDD PHVT12LL L=6E-08 W=2.5E-06
M87 WL[3] 72 VDD VDD PHVT12LL L=6E-08 W=2.5E-06
M88 VDD 72 WL[3] VDD PHVT12LL L=6E-08 W=2.5E-06
M89 WL[4] 73 VDD VDD PHVT12LL L=6E-08 W=2.5E-06
M90 VDD 73 WL[4] VDD PHVT12LL L=6E-08 W=2.5E-06
M91 WL[5] 74 VDD VDD PHVT12LL L=6E-08 W=2.5E-06
M92 VDD 74 WL[5] VDD PHVT12LL L=6E-08 W=2.5E-06
M93 WL[6] 75 VDD VDD PHVT12LL L=6E-08 W=2.5E-06
M94 VDD 75 WL[6] VDD PHVT12LL L=6E-08 W=2.5E-06
M95 WL[7] 76 VDD VDD PHVT12LL L=6E-08 W=2.5E-06
M96 VDD 76 WL[7] VDD PHVT12LL L=6E-08 W=2.5E-06
M97 VDD 52 50 VDD P12LL L=6E-08 W=1E-06
M98 50 52 VDD VDD P12LL L=6E-08 W=1E-06
M99 VDD 52 50 VDD P12LL L=6E-08 W=1E-06
M100 52 49 VDD VDD P12LL L=6E-08 W=1E-06
M101 VDD 49 52 VDD P12LL L=6E-08 W=1E-06
M102 52 49 VDD VDD P12LL L=6E-08 W=1E-06
M103 VDD PXA 49 VDD P12LL L=6E-08 W=5E-07
M104 49 PXB VDD VDD P12LL L=6E-08 W=5E-07
M105 VDD PXC 49 VDD P12LL L=6E-08 W=5E-07
M106 53 52 VDD VDD P12LL L=6E-08 W=4E-07
M107 VDD 52 54 VDD P12LL L=6E-08 W=4E-07
M108 56 52 VDD VDD P12LL L=6E-08 W=4E-07
M109 VDD 52 58 VDD P12LL L=6E-08 W=4E-07
M110 57 52 VDD VDD P12LL L=6E-08 W=4E-07
M111 VDD 52 59 VDD P12LL L=6E-08 W=4E-07
M112 60 52 VDD VDD P12LL L=6E-08 W=4E-07
M113 VDD 52 55 VDD P12LL L=6E-08 W=4E-07
M114 58 50 FCKX[3] VDD P12LL L=6E-08 W=4E-07
M115 59 50 FCKX[5] VDD P12LL L=6E-08 W=4E-07
M116 FCKX[7] 50 55 VDD P12LL L=6E-08 W=4E-07
M117 54 50 FCKX[1] VDD P12LL L=6E-08 W=4E-07
M118 53 50 FCKX[0] VDD P12LL L=6E-08 W=4E-07
M119 56 50 FCKX[2] VDD P12LL L=6E-08 W=4E-07
M120 57 50 FCKX[4] VDD P12LL L=6E-08 W=4E-07
M121 60 50 FCKX[6] VDD P12LL L=6E-08 W=4E-07
M122 61 53 VDD VDD P12LL L=6E-08 W=7E-07
M123 VDD 53 61 VDD P12LL L=6E-08 W=7E-07
M124 62 54 VDD VDD P12LL L=6E-08 W=7E-07
M125 VDD 54 62 VDD P12LL L=6E-08 W=7E-07
M126 63 56 VDD VDD P12LL L=6E-08 W=7E-07
M127 VDD 56 63 VDD P12LL L=6E-08 W=7E-07
M128 64 58 VDD VDD P12LL L=6E-08 W=7E-07
M129 VDD 58 64 VDD P12LL L=6E-08 W=7E-07
M130 65 57 VDD VDD P12LL L=6E-08 W=7E-07
M131 VDD 57 65 VDD P12LL L=6E-08 W=7E-07
M132 66 59 VDD VDD P12LL L=6E-08 W=7E-07
M133 VDD 59 66 VDD P12LL L=6E-08 W=7E-07
M134 67 60 VDD VDD P12LL L=6E-08 W=7E-07
M135 VDD 60 67 VDD P12LL L=6E-08 W=7E-07
M136 68 55 VDD VDD P12LL L=6E-08 W=7E-07
M137 VDD 55 68 VDD P12LL L=6E-08 W=7E-07
M138 69 61 VDD VDD P12LL L=6E-08 W=1.5E-06
M139 VDD 61 69 VDD P12LL L=6E-08 W=1.5E-06
M140 70 62 VDD VDD P12LL L=6E-08 W=1.5E-06
M141 VDD 62 70 VDD P12LL L=6E-08 W=1.5E-06
M142 71 63 VDD VDD P12LL L=6E-08 W=1.5E-06
M143 VDD 63 71 VDD P12LL L=6E-08 W=1.5E-06
M144 72 64 VDD VDD P12LL L=6E-08 W=1.5E-06
M145 VDD 64 72 VDD P12LL L=6E-08 W=1.5E-06
M146 73 65 VDD VDD P12LL L=6E-08 W=1.5E-06
M147 VDD 65 73 VDD P12LL L=6E-08 W=1.5E-06
M148 74 66 VDD VDD P12LL L=6E-08 W=1.5E-06
M149 VDD 66 74 VDD P12LL L=6E-08 W=1.5E-06
M150 75 67 VDD VDD P12LL L=6E-08 W=1.5E-06
M151 VDD 67 75 VDD P12LL L=6E-08 W=1.5E-06
M152 76 68 VDD VDD P12LL L=6E-08 W=1.5E-06
M153 VDD 68 76 VDD P12LL L=6E-08 W=1.5E-06
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    S55NLLGDPH_X512Y8D16_BW_XDEC64
* View Name:    schematic
************************************************************************

.SUBCKT S55NLLGDPH_X512Y8D16_BW_XDEC64 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[3] PXA[2]
+PXA[1] PXA[0] PXB[3] PXB[2] PXB[1] PXB[0] PXC[3] PXC[2] PXC[1] PXC[0]
+VDD VSS WL[511] WL[510] WL[509] WL[508] WL[507] WL[506] WL[505] WL[504]
+WL[503] WL[502] WL[501] WL[500] WL[499] WL[498] WL[497] WL[496] WL[495] WL[494]
+WL[493] WL[492] WL[491] WL[490] WL[489] WL[488] WL[487] WL[486] WL[485] WL[484]
+WL[483] WL[482] WL[481] WL[480] WL[479] WL[478] WL[477] WL[476] WL[475] WL[474]
+WL[473] WL[472] WL[471] WL[470] WL[469] WL[468] WL[467] WL[466] WL[465] WL[464]
+WL[463] WL[462] WL[461] WL[460] WL[459] WL[458] WL[457] WL[456] WL[455] WL[454]
+WL[453] WL[452] WL[451] WL[450] WL[449] WL[448] WL[447] WL[446] WL[445] WL[444]
+WL[443] WL[442] WL[441] WL[440] WL[439] WL[438] WL[437] WL[436] WL[435] WL[434]
+WL[433] WL[432] WL[431] WL[430] WL[429] WL[428] WL[427] WL[426] WL[425] WL[424]
+WL[423] WL[422] WL[421] WL[420] WL[419] WL[418] WL[417] WL[416] WL[415] WL[414]
+WL[413] WL[412] WL[411] WL[410] WL[409] WL[408] WL[407] WL[406] WL[405] WL[404]
+WL[403] WL[402] WL[401] WL[400] WL[399] WL[398] WL[397] WL[396] WL[395] WL[394]
+WL[393] WL[392] WL[391] WL[390] WL[389] WL[388] WL[387] WL[386] WL[385] WL[384]
+WL[383] WL[382] WL[381] WL[380] WL[379] WL[378] WL[377] WL[376] WL[375] WL[374]
+WL[373] WL[372] WL[371] WL[370] WL[369] WL[368] WL[367] WL[366] WL[365] WL[364]
+WL[363] WL[362] WL[361] WL[360] WL[359] WL[358] WL[357] WL[356] WL[355] WL[354]
+WL[353] WL[352] WL[351] WL[350] WL[349] WL[348] WL[347] WL[346] WL[345] WL[344]
+WL[343] WL[342] WL[341] WL[340] WL[339] WL[338] WL[337] WL[336] WL[335] WL[334]
+WL[333] WL[332] WL[331] WL[330] WL[329] WL[328] WL[327] WL[326] WL[325] WL[324]
+WL[323] WL[322] WL[321] WL[320] WL[319] WL[318] WL[317] WL[316] WL[315] WL[314]
+WL[313] WL[312] WL[311] WL[310] WL[309] WL[308] WL[307] WL[306] WL[305] WL[304]
+WL[303] WL[302] WL[301] WL[300] WL[299] WL[298] WL[297] WL[296] WL[295] WL[294]
+WL[293] WL[292] WL[291] WL[290] WL[289] WL[288] WL[287] WL[286] WL[285] WL[284]
+WL[283] WL[282] WL[281] WL[280] WL[279] WL[278] WL[277] WL[276] WL[275] WL[274]
+WL[273] WL[272] WL[271] WL[270] WL[269] WL[268] WL[267] WL[266] WL[265] WL[264]
+WL[263] WL[262] WL[261] WL[260] WL[259] WL[258] WL[257] WL[256] WL[255] WL[254]
+WL[253] WL[252] WL[251] WL[250] WL[249] WL[248] WL[247] WL[246] WL[245] WL[244]
+WL[243] WL[242] WL[241] WL[240] WL[239] WL[238] WL[237] WL[236] WL[235] WL[234]
+WL[233] WL[232] WL[231] WL[230] WL[229] WL[228] WL[227] WL[226] WL[225] WL[224]
+WL[223] WL[222] WL[221] WL[220] WL[219] WL[218] WL[217] WL[216] WL[215] WL[214]
+WL[213] WL[212] WL[211] WL[210] WL[209] WL[208] WL[207] WL[206] WL[205] WL[204]
+WL[203] WL[202] WL[201] WL[200] WL[199] WL[198] WL[197] WL[196] WL[195] WL[194]
+WL[193] WL[192] WL[191] WL[190] WL[189] WL[188] WL[187] WL[186] WL[185] WL[184]
+WL[183] WL[182] WL[181] WL[180] WL[179] WL[178] WL[177] WL[176] WL[175] WL[174]
+WL[173] WL[172] WL[171] WL[170] WL[169] WL[168] WL[167] WL[166] WL[165] WL[164]
+WL[163] WL[162] WL[161] WL[160] WL[159] WL[158] WL[157] WL[156] WL[155] WL[154]
+WL[153] WL[152] WL[151] WL[150] WL[149] WL[148] WL[147] WL[146] WL[145] WL[144]
+WL[143] WL[142] WL[141] WL[140] WL[139] WL[138] WL[137] WL[136] WL[135] WL[134]
+WL[133] WL[132] WL[131] WL[130] WL[129] WL[128] WL[127] WL[126] WL[125] WL[124]
+WL[123] WL[122] WL[121] WL[120] WL[119] WL[118] WL[117] WL[116] WL[115] WL[114]
+WL[113] WL[112] WL[111] WL[110] WL[109] WL[108] WL[107] WL[106] WL[105] WL[104]
+WL[103] WL[102] WL[101] WL[100] WL[99] WL[98] WL[97] WL[96] WL[95] WL[94]
+WL[93] WL[92] WL[91] WL[90] WL[89] WL[88] WL[87] WL[86] WL[85] WL[84]
+WL[83] WL[82] WL[81] WL[80] WL[79] WL[78] WL[77] WL[76] WL[75] WL[74]
+WL[73] WL[72] WL[71] WL[70] WL[69] WL[68] WL[67] WL[66] WL[65] WL[64]
+WL[63] WL[62] WL[61] WL[60] WL[59] WL[58] WL[57] WL[56] WL[55] WL[54]
+WL[53] WL[52] WL[51] WL[50] WL[49] WL[48] WL[47] WL[46] WL[45] WL[44]
+WL[43] WL[42] WL[41] WL[40] WL[39] WL[38] WL[37] WL[36] WL[35] WL[34]
+WL[33] WL[32] WL[31] WL[30] WL[29] WL[28] WL[27] WL[26] WL[25] WL[24]
+WL[23] WL[22] WL[21] WL[20] WL[19] WL[18] WL[17] WL[16] WL[15] WL[14]
+WL[13] WL[12] WL[11] WL[10] WL[9] WL[8] WL[7] WL[6] WL[5] WL[4]
+WL[3] WL[2] WL[1] WL[0]
XI0 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[3] PXB[3]
+PXC[3] VDD VSS WL[511] WL[510] WL[509] WL[508] WL[507] WL[506] WL[505]
+WL[504] S55NLLGDPH_X512Y8D16_BW_XDEC
XI1 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[2] PXB[3]
+PXC[3] VDD VSS WL[503] WL[502] WL[501] WL[500] WL[499] WL[498] WL[497]
+WL[496] S55NLLGDPH_X512Y8D16_BW_XDEC
XI2 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[1] PXB[3]
+PXC[3] VDD VSS WL[495] WL[494] WL[493] WL[492] WL[491] WL[490] WL[489]
+WL[488] S55NLLGDPH_X512Y8D16_BW_XDEC
XI3 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[0] PXB[3]
+PXC[3] VDD VSS WL[487] WL[486] WL[485] WL[484] WL[483] WL[482] WL[481]
+WL[480] S55NLLGDPH_X512Y8D16_BW_XDEC
XI4 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[3] PXB[2]
+PXC[3] VDD VSS WL[479] WL[478] WL[477] WL[476] WL[475] WL[474] WL[473]
+WL[472] S55NLLGDPH_X512Y8D16_BW_XDEC
XI5 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[2] PXB[2]
+PXC[3] VDD VSS WL[471] WL[470] WL[469] WL[468] WL[467] WL[466] WL[465]
+WL[464] S55NLLGDPH_X512Y8D16_BW_XDEC
XI6 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[1] PXB[2]
+PXC[3] VDD VSS WL[463] WL[462] WL[461] WL[460] WL[459] WL[458] WL[457]
+WL[456] S55NLLGDPH_X512Y8D16_BW_XDEC
XI7 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[0] PXB[2]
+PXC[3] VDD VSS WL[455] WL[454] WL[453] WL[452] WL[451] WL[450] WL[449]
+WL[448] S55NLLGDPH_X512Y8D16_BW_XDEC
XI8 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[3] PXB[1]
+PXC[3] VDD VSS WL[447] WL[446] WL[445] WL[444] WL[443] WL[442] WL[441]
+WL[440] S55NLLGDPH_X512Y8D16_BW_XDEC
XI9 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[2] PXB[1]
+PXC[3] VDD VSS WL[439] WL[438] WL[437] WL[436] WL[435] WL[434] WL[433]
+WL[432] S55NLLGDPH_X512Y8D16_BW_XDEC
XI10 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[1] PXB[1]
+PXC[3] VDD VSS WL[431] WL[430] WL[429] WL[428] WL[427] WL[426] WL[425]
+WL[424] S55NLLGDPH_X512Y8D16_BW_XDEC
XI11 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[0] PXB[1]
+PXC[3] VDD VSS WL[423] WL[422] WL[421] WL[420] WL[419] WL[418] WL[417]
+WL[416] S55NLLGDPH_X512Y8D16_BW_XDEC
XI12 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[3] PXB[0]
+PXC[3] VDD VSS WL[415] WL[414] WL[413] WL[412] WL[411] WL[410] WL[409]
+WL[408] S55NLLGDPH_X512Y8D16_BW_XDEC
XI13 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[2] PXB[0]
+PXC[3] VDD VSS WL[407] WL[406] WL[405] WL[404] WL[403] WL[402] WL[401]
+WL[400] S55NLLGDPH_X512Y8D16_BW_XDEC
XI14 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[1] PXB[0]
+PXC[3] VDD VSS WL[399] WL[398] WL[397] WL[396] WL[395] WL[394] WL[393]
+WL[392] S55NLLGDPH_X512Y8D16_BW_XDEC
XI15 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[0] PXB[0]
+PXC[3] VDD VSS WL[391] WL[390] WL[389] WL[388] WL[387] WL[386] WL[385]
+WL[384] S55NLLGDPH_X512Y8D16_BW_XDEC
XI16 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[3] PXB[3]
+PXC[2] VDD VSS WL[383] WL[382] WL[381] WL[380] WL[379] WL[378] WL[377]
+WL[376] S55NLLGDPH_X512Y8D16_BW_XDEC
XI17 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[2] PXB[3]
+PXC[2] VDD VSS WL[375] WL[374] WL[373] WL[372] WL[371] WL[370] WL[369]
+WL[368] S55NLLGDPH_X512Y8D16_BW_XDEC
XI18 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[1] PXB[3]
+PXC[2] VDD VSS WL[367] WL[366] WL[365] WL[364] WL[363] WL[362] WL[361]
+WL[360] S55NLLGDPH_X512Y8D16_BW_XDEC
XI19 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[0] PXB[3]
+PXC[2] VDD VSS WL[359] WL[358] WL[357] WL[356] WL[355] WL[354] WL[353]
+WL[352] S55NLLGDPH_X512Y8D16_BW_XDEC
XI20 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[3] PXB[2]
+PXC[2] VDD VSS WL[351] WL[350] WL[349] WL[348] WL[347] WL[346] WL[345]
+WL[344] S55NLLGDPH_X512Y8D16_BW_XDEC
XI21 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[2] PXB[2]
+PXC[2] VDD VSS WL[343] WL[342] WL[341] WL[340] WL[339] WL[338] WL[337]
+WL[336] S55NLLGDPH_X512Y8D16_BW_XDEC
XI22 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[1] PXB[2]
+PXC[2] VDD VSS WL[335] WL[334] WL[333] WL[332] WL[331] WL[330] WL[329]
+WL[328] S55NLLGDPH_X512Y8D16_BW_XDEC
XI23 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[0] PXB[2]
+PXC[2] VDD VSS WL[327] WL[326] WL[325] WL[324] WL[323] WL[322] WL[321]
+WL[320] S55NLLGDPH_X512Y8D16_BW_XDEC
XI24 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[3] PXB[1]
+PXC[2] VDD VSS WL[319] WL[318] WL[317] WL[316] WL[315] WL[314] WL[313]
+WL[312] S55NLLGDPH_X512Y8D16_BW_XDEC
XI25 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[2] PXB[1]
+PXC[2] VDD VSS WL[311] WL[310] WL[309] WL[308] WL[307] WL[306] WL[305]
+WL[304] S55NLLGDPH_X512Y8D16_BW_XDEC
XI26 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[1] PXB[1]
+PXC[2] VDD VSS WL[303] WL[302] WL[301] WL[300] WL[299] WL[298] WL[297]
+WL[296] S55NLLGDPH_X512Y8D16_BW_XDEC
XI27 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[0] PXB[1]
+PXC[2] VDD VSS WL[295] WL[294] WL[293] WL[292] WL[291] WL[290] WL[289]
+WL[288] S55NLLGDPH_X512Y8D16_BW_XDEC
XI28 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[3] PXB[0]
+PXC[2] VDD VSS WL[287] WL[286] WL[285] WL[284] WL[283] WL[282] WL[281]
+WL[280] S55NLLGDPH_X512Y8D16_BW_XDEC
XI29 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[2] PXB[0]
+PXC[2] VDD VSS WL[279] WL[278] WL[277] WL[276] WL[275] WL[274] WL[273]
+WL[272] S55NLLGDPH_X512Y8D16_BW_XDEC
XI30 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[1] PXB[0]
+PXC[2] VDD VSS WL[271] WL[270] WL[269] WL[268] WL[267] WL[266] WL[265]
+WL[264] S55NLLGDPH_X512Y8D16_BW_XDEC
XI31 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[0] PXB[0]
+PXC[2] VDD VSS WL[263] WL[262] WL[261] WL[260] WL[259] WL[258] WL[257]
+WL[256] S55NLLGDPH_X512Y8D16_BW_XDEC
XI32 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[3] PXB[3]
+PXC[1] VDD VSS WL[255] WL[254] WL[253] WL[252] WL[251] WL[250] WL[249]
+WL[248] S55NLLGDPH_X512Y8D16_BW_XDEC
XI33 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[2] PXB[3]
+PXC[1] VDD VSS WL[247] WL[246] WL[245] WL[244] WL[243] WL[242] WL[241]
+WL[240] S55NLLGDPH_X512Y8D16_BW_XDEC
XI34 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[1] PXB[3]
+PXC[1] VDD VSS WL[239] WL[238] WL[237] WL[236] WL[235] WL[234] WL[233]
+WL[232] S55NLLGDPH_X512Y8D16_BW_XDEC
XI35 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[0] PXB[3]
+PXC[1] VDD VSS WL[231] WL[230] WL[229] WL[228] WL[227] WL[226] WL[225]
+WL[224] S55NLLGDPH_X512Y8D16_BW_XDEC
XI36 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[3] PXB[2]
+PXC[1] VDD VSS WL[223] WL[222] WL[221] WL[220] WL[219] WL[218] WL[217]
+WL[216] S55NLLGDPH_X512Y8D16_BW_XDEC
XI37 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[2] PXB[2]
+PXC[1] VDD VSS WL[215] WL[214] WL[213] WL[212] WL[211] WL[210] WL[209]
+WL[208] S55NLLGDPH_X512Y8D16_BW_XDEC
XI38 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[1] PXB[2]
+PXC[1] VDD VSS WL[207] WL[206] WL[205] WL[204] WL[203] WL[202] WL[201]
+WL[200] S55NLLGDPH_X512Y8D16_BW_XDEC
XI39 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[0] PXB[2]
+PXC[1] VDD VSS WL[199] WL[198] WL[197] WL[196] WL[195] WL[194] WL[193]
+WL[192] S55NLLGDPH_X512Y8D16_BW_XDEC
XI40 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[3] PXB[1]
+PXC[1] VDD VSS WL[191] WL[190] WL[189] WL[188] WL[187] WL[186] WL[185]
+WL[184] S55NLLGDPH_X512Y8D16_BW_XDEC
XI41 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[2] PXB[1]
+PXC[1] VDD VSS WL[183] WL[182] WL[181] WL[180] WL[179] WL[178] WL[177]
+WL[176] S55NLLGDPH_X512Y8D16_BW_XDEC
XI42 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[1] PXB[1]
+PXC[1] VDD VSS WL[175] WL[174] WL[173] WL[172] WL[171] WL[170] WL[169]
+WL[168] S55NLLGDPH_X512Y8D16_BW_XDEC
XI43 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[0] PXB[1]
+PXC[1] VDD VSS WL[167] WL[166] WL[165] WL[164] WL[163] WL[162] WL[161]
+WL[160] S55NLLGDPH_X512Y8D16_BW_XDEC
XI44 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[3] PXB[0]
+PXC[1] VDD VSS WL[159] WL[158] WL[157] WL[156] WL[155] WL[154] WL[153]
+WL[152] S55NLLGDPH_X512Y8D16_BW_XDEC
XI45 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[2] PXB[0]
+PXC[1] VDD VSS WL[151] WL[150] WL[149] WL[148] WL[147] WL[146] WL[145]
+WL[144] S55NLLGDPH_X512Y8D16_BW_XDEC
XI46 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[1] PXB[0]
+PXC[1] VDD VSS WL[143] WL[142] WL[141] WL[140] WL[139] WL[138] WL[137]
+WL[136] S55NLLGDPH_X512Y8D16_BW_XDEC
XI47 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[0] PXB[0]
+PXC[1] VDD VSS WL[135] WL[134] WL[133] WL[132] WL[131] WL[130] WL[129]
+WL[128] S55NLLGDPH_X512Y8D16_BW_XDEC
XI48 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[3] PXB[3]
+PXC[0] VDD VSS WL[127] WL[126] WL[125] WL[124] WL[123] WL[122] WL[121]
+WL[120] S55NLLGDPH_X512Y8D16_BW_XDEC
XI49 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[2] PXB[3]
+PXC[0] VDD VSS WL[119] WL[118] WL[117] WL[116] WL[115] WL[114] WL[113]
+WL[112] S55NLLGDPH_X512Y8D16_BW_XDEC
XI50 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[1] PXB[3]
+PXC[0] VDD VSS WL[111] WL[110] WL[109] WL[108] WL[107] WL[106] WL[105]
+WL[104] S55NLLGDPH_X512Y8D16_BW_XDEC
XI51 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[0] PXB[3]
+PXC[0] VDD VSS WL[103] WL[102] WL[101] WL[100] WL[99] WL[98] WL[97]
+WL[96] S55NLLGDPH_X512Y8D16_BW_XDEC
XI52 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[3] PXB[2]
+PXC[0] VDD VSS WL[95] WL[94] WL[93] WL[92] WL[91] WL[90] WL[89]
+WL[88] S55NLLGDPH_X512Y8D16_BW_XDEC
XI53 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[2] PXB[2]
+PXC[0] VDD VSS WL[87] WL[86] WL[85] WL[84] WL[83] WL[82] WL[81]
+WL[80] S55NLLGDPH_X512Y8D16_BW_XDEC
XI54 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[1] PXB[2]
+PXC[0] VDD VSS WL[79] WL[78] WL[77] WL[76] WL[75] WL[74] WL[73]
+WL[72] S55NLLGDPH_X512Y8D16_BW_XDEC
XI55 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[0] PXB[2]
+PXC[0] VDD VSS WL[71] WL[70] WL[69] WL[68] WL[67] WL[66] WL[65]
+WL[64] S55NLLGDPH_X512Y8D16_BW_XDEC
XI56 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[3] PXB[1]
+PXC[0] VDD VSS WL[63] WL[62] WL[61] WL[60] WL[59] WL[58] WL[57]
+WL[56] S55NLLGDPH_X512Y8D16_BW_XDEC
XI57 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[2] PXB[1]
+PXC[0] VDD VSS WL[55] WL[54] WL[53] WL[52] WL[51] WL[50] WL[49]
+WL[48] S55NLLGDPH_X512Y8D16_BW_XDEC
XI58 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[1] PXB[1]
+PXC[0] VDD VSS WL[47] WL[46] WL[45] WL[44] WL[43] WL[42] WL[41]
+WL[40] S55NLLGDPH_X512Y8D16_BW_XDEC
XI59 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[0] PXB[1]
+PXC[0] VDD VSS WL[39] WL[38] WL[37] WL[36] WL[35] WL[34] WL[33]
+WL[32] S55NLLGDPH_X512Y8D16_BW_XDEC
XI60 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[3] PXB[0]
+PXC[0] VDD VSS WL[31] WL[30] WL[29] WL[28] WL[27] WL[26] WL[25]
+WL[24] S55NLLGDPH_X512Y8D16_BW_XDEC
XI61 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[2] PXB[0]
+PXC[0] VDD VSS WL[23] WL[22] WL[21] WL[20] WL[19] WL[18] WL[17]
+WL[16] S55NLLGDPH_X512Y8D16_BW_XDEC
XI62 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[1] PXB[0]
+PXC[0] VDD VSS WL[15] WL[14] WL[13] WL[12] WL[11] WL[10] WL[9]
+WL[8] S55NLLGDPH_X512Y8D16_BW_XDEC
XI63 FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[0] PXB[0]
+PXC[0] VDD VSS WL[7] WL[6] WL[5] WL[4] WL[3] WL[2] WL[1]
+WL[0] S55NLLGDPH_X512Y8D16_BW_XDEC
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    S55NLLGDPH_X512Y8D16_BW_PX4
* View Name:    schematic
************************************************************************

.SUBCKT S55NLLGDPH_X512Y8D16_BW_PX4 A[0] A[1] CLK CLKX PX[3] PX[2] PX[1] PX[0] VDD VSS
M0 PX[3] 38 VSS VSS N12LL L=6E-08 W=1.5E-06
M1 40 PX[2] VSS VSS N12LL L=6E-07 W=1.2E-07
M2 50 47 37 VSS N12LL L=6E-08 W=1.495E-06
M3 51 A[0] 36 VSS N12LL L=6E-08 W=4E-07
M4 38 CLKX 37 VSS N12LL L=6E-08 W=2.5E-06
M5 VSS PX[3] 38 VSS N12LL L=6E-07 W=1.2E-07
M6 VSS 38 PX[3] VSS N12LL L=6E-08 W=1.5E-06
M7 VSS 43 50 VSS N12LL L=6E-08 W=1.495E-06
M8 VSS 36 47 VSS N12LL L=6E-08 W=7E-07
M9 VSS VDD 51 VSS N12LL L=3E-07 W=4E-07
M10 52 43 VSS VSS N12LL L=6E-08 W=1.495E-06
M11 PX[2] 40 VSS VSS N12LL L=6E-08 W=1.5E-06
M12 32 47 VSS VSS N12LL L=6E-08 W=7E-07
M13 39 CLKX 40 VSS N12LL L=6E-08 W=2.5E-06
M14 39 32 52 VSS N12LL L=6E-08 W=1.495E-06
M15 VSS 40 PX[2] VSS N12LL L=6E-08 W=1.5E-06
M16 PX[0] 41 VSS VSS N12LL L=6E-08 W=1.5E-06
M17 46 PX[1] VSS VSS N12LL L=6E-07 W=1.2E-07
M18 53 32 42 VSS N12LL L=6E-08 W=1.495E-06
M19 41 CLKX 42 VSS N12LL L=6E-08 W=2.5E-06
M20 54 VDD VSS VSS N12LL L=3E-07 W=4E-07
M21 VSS 49 43 VSS N12LL L=6E-08 W=7E-07
M22 VSS PX[0] 41 VSS N12LL L=6E-07 W=1.2E-07
M23 VSS 41 PX[0] VSS N12LL L=6E-08 W=1.5E-06
M24 VSS 45 53 VSS N12LL L=6E-08 W=1.495E-06
M25 45 43 VSS VSS N12LL L=6E-08 W=7E-07
M26 55 45 VSS VSS N12LL L=6E-08 W=1.495E-06
M27 PX[1] 46 VSS VSS N12LL L=6E-08 W=1.5E-06
M28 48 CLKX 46 VSS N12LL L=6E-08 W=2.5E-06
M29 49 A[1] 54 VSS N12LL L=6E-08 W=4E-07
M30 48 47 55 VSS N12LL L=6E-08 W=1.495E-06
M31 VSS 46 PX[1] VSS N12LL L=6E-08 W=1.5E-06
M32 PX[3] 38 VDD VDD P12LL L=6E-08 W=3.5E-06
M33 37 47 VDD VDD P12LL L=6E-08 W=1.5E-06
M34 56 A[0] 36 VDD P12LL L=6E-08 W=4E-07
M35 38 CLK 37 VDD P12LL L=6E-08 W=2.5E-06
M36 40 PX[2] VDD VDD P12LL L=3E-07 W=1.2E-07
M37 VDD 38 PX[3] VDD P12LL L=6E-08 W=3.5E-06
M38 VDD 43 37 VDD P12LL L=6E-08 W=1.5E-06
M39 VDD 36 47 VDD P12LL L=6E-08 W=1.4E-06
M40 VDD VSS 56 VDD P12LL L=1E-07 W=4E-07
M41 VDD PX[3] 38 VDD P12LL L=3E-07 W=1.2E-07
M42 39 43 VDD VDD P12LL L=6E-08 W=1.5E-06
M43 PX[2] 40 VDD VDD P12LL L=6E-08 W=3.5E-06
M44 32 47 VDD VDD P12LL L=6E-08 W=1.4E-06
M45 39 CLK 40 VDD P12LL L=6E-08 W=2.5E-06
M46 VDD 32 39 VDD P12LL L=6E-08 W=1.5E-06
M47 VDD 40 PX[2] VDD P12LL L=6E-08 W=3.5E-06
M48 PX[0] 41 VDD VDD P12LL L=6E-08 W=3.5E-06
M49 42 32 VDD VDD P12LL L=6E-08 W=1.5E-06
M50 46 PX[1] VDD VDD P12LL L=3E-07 W=1.2E-07
M51 41 CLK 42 VDD P12LL L=6E-08 W=2.5E-06
M52 57 VSS VDD VDD P12LL L=1E-07 W=4E-07
M53 VDD 49 43 VDD P12LL L=6E-08 W=1.4E-06
M54 VDD 41 PX[0] VDD P12LL L=6E-08 W=3.5E-06
M55 VDD 45 42 VDD P12LL L=6E-08 W=1.5E-06
M56 VDD PX[0] 41 VDD P12LL L=3E-07 W=1.2E-07
M57 45 43 VDD VDD P12LL L=6E-08 W=1.4E-06
M58 48 45 VDD VDD P12LL L=6E-08 W=1.5E-06
M59 PX[1] 46 VDD VDD P12LL L=6E-08 W=3.5E-06
M60 48 CLK 46 VDD P12LL L=6E-08 W=2.5E-06
M61 49 A[1] 57 VDD P12LL L=6E-08 W=4E-07
M62 VDD 47 48 VDD P12LL L=6E-08 W=1.5E-06
M63 VDD 46 PX[1] VDD P12LL L=6E-08 W=3.5E-06
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    S55NLLGDPH_X512Y8D16_BW_YPREDEC_Y8
* View Name:    schematic
************************************************************************

.SUBCKT S55NLLGDPH_X512Y8D16_BW_YPREDEC_Y8 A[0] A[1] A[2] CLK CLKX VDD VSS YCKX YX[7] YX[6]
+YX[5] YX[4] YX[3] YX[2] YX[1] YX[0]
M0 51 64 VSS VSS N12LL L=6E-08 W=4E-07
M1 YX[3] 51 YCKX VSS N12LL L=6E-08 W=1.25E-06
M2 65 CLKX 64 VSS N12LL L=6E-08 W=5E-07
M3 VSS 51 64 VSS N12LL L=6E-07 W=1.2E-07
M4 VSS 64 51 VSS N12LL L=6E-08 W=4E-07
M5 YCKX 51 YX[3] VSS N12LL L=6E-08 W=1.25E-06
M6 94 6 65 VSS N12LL L=6E-08 W=1E-06
M7 64 CLKX 65 VSS N12LL L=6E-08 W=5E-07
M8 51 64 VSS VSS N12LL L=6E-08 W=4E-07
M9 YX[3] 51 YCKX VSS N12LL L=6E-08 W=1.25E-06
M10 95 5 94 VSS N12LL L=6E-08 W=1E-06
M11 65 CLKX 64 VSS N12LL L=6E-08 W=5E-07
M12 73 87 VSS VSS N12LL L=6E-08 W=5E-07
M13 VSS 73 95 VSS N12LL L=6E-08 W=1E-06
M14 VSS 64 51 VSS N12LL L=6E-08 W=4E-07
M15 YCKX 51 YX[3] VSS N12LL L=6E-08 W=1.25E-06
M16 VSS 87 73 VSS N12LL L=6E-08 W=5E-07
M17 96 73 VSS VSS N12LL L=6E-08 W=1E-06
M18 52 67 VSS VSS N12LL L=6E-08 W=4E-07
M19 YX[1] 52 YCKX VSS N12LL L=6E-08 W=1.25E-06
M20 67 52 VSS VSS N12LL L=6E-07 W=1.2E-07
M21 67 CLKX 53 VSS N12LL L=6E-08 W=5E-07
M22 87 69 VSS VSS N12LL L=6E-08 W=5E-07
M23 97 5 96 VSS N12LL L=6E-08 W=1E-06
M24 VSS 67 52 VSS N12LL L=6E-08 W=4E-07
M25 YCKX 52 YX[1] VSS N12LL L=6E-08 W=1.25E-06
M26 53 CLKX 67 VSS N12LL L=6E-08 W=5E-07
M27 53 4 97 VSS N12LL L=6E-08 W=1E-06
M28 VSS 69 87 VSS N12LL L=6E-08 W=5E-07
M29 52 67 VSS VSS N12LL L=6E-08 W=4E-07
M30 YX[1] 52 YCKX VSS N12LL L=6E-08 W=1.25E-06
M31 67 CLKX 53 VSS N12LL L=6E-08 W=5E-07
M32 VSS 67 52 VSS N12LL L=6E-08 W=4E-07
M33 YCKX 52 YX[1] VSS N12LL L=6E-08 W=1.25E-06
M34 98 A[2] 69 VSS N12LL L=6E-08 W=4E-07
M35 55 71 VSS VSS N12LL L=6E-08 W=4E-07
M36 YX[0] 55 YCKX VSS N12LL L=6E-08 W=1.25E-06
M37 54 CLKX 71 VSS N12LL L=6E-08 W=5E-07
M38 VSS VDD 98 VSS N12LL L=3E-07 W=4E-07
M39 VSS 55 71 VSS N12LL L=6E-07 W=1.2E-07
M40 VSS 71 55 VSS N12LL L=6E-08 W=4E-07
M41 YCKX 55 YX[0] VSS N12LL L=6E-08 W=1.25E-06
M42 99 4 54 VSS N12LL L=6E-08 W=1E-06
M43 71 CLKX 54 VSS N12LL L=6E-08 W=5E-07
M44 55 71 VSS VSS N12LL L=6E-08 W=4E-07
M45 YX[0] 55 YCKX VSS N12LL L=6E-08 W=1.25E-06
M46 100 88 99 VSS N12LL L=6E-08 W=1E-06
M47 54 CLKX 71 VSS N12LL L=6E-08 W=5E-07
M48 VSS 73 100 VSS N12LL L=6E-08 W=1E-06
M49 VSS 71 55 VSS N12LL L=6E-08 W=4E-07
M50 YCKX 55 YX[0] VSS N12LL L=6E-08 W=1.25E-06
M51 101 73 VSS VSS N12LL L=6E-08 W=1E-06
M52 56 74 VSS VSS N12LL L=6E-08 W=4E-07
M53 YX[2] 56 YCKX VSS N12LL L=6E-08 W=1.25E-06
M54 74 56 VSS VSS N12LL L=6E-07 W=1.2E-07
M55 74 CLKX 75 VSS N12LL L=6E-08 W=5E-07
M56 102 88 101 VSS N12LL L=6E-08 W=1E-06
M57 103 VDD VSS VSS N12LL L=3E-07 W=4E-07
M58 VSS 74 56 VSS N12LL L=6E-08 W=4E-07
M59 YCKX 56 YX[2] VSS N12LL L=6E-08 W=1.25E-06
M60 75 CLKX 74 VSS N12LL L=6E-08 W=5E-07
M61 75 6 102 VSS N12LL L=6E-08 W=1E-06
M62 56 74 VSS VSS N12LL L=6E-08 W=4E-07
M63 YX[2] 56 YCKX VSS N12LL L=6E-08 W=1.25E-06
M64 74 CLKX 75 VSS N12LL L=6E-08 W=5E-07
M65 78 A[1] 103 VSS N12LL L=6E-08 W=4E-07
M66 VSS 74 56 VSS N12LL L=6E-08 W=4E-07
M67 YCKX 56 YX[2] VSS N12LL L=6E-08 W=1.25E-06
M68 58 79 VSS VSS N12LL L=6E-08 W=4E-07
M69 YX[7] 58 YCKX VSS N12LL L=6E-08 W=1.25E-06
M70 57 CLKX 79 VSS N12LL L=6E-08 W=5E-07
M71 6 78 VSS VSS N12LL L=6E-08 W=5E-07
M72 VSS 58 79 VSS N12LL L=6E-07 W=1.2E-07
M73 VSS 79 58 VSS N12LL L=6E-08 W=4E-07
M74 YCKX 58 YX[7] VSS N12LL L=6E-08 W=1.25E-06
M75 104 6 57 VSS N12LL L=6E-08 W=1E-06
M76 79 CLKX 57 VSS N12LL L=6E-08 W=5E-07
M77 VSS 78 6 VSS N12LL L=6E-08 W=5E-07
M78 58 79 VSS VSS N12LL L=6E-08 W=4E-07
M79 YX[7] 58 YCKX VSS N12LL L=6E-08 W=1.25E-06
M80 105 5 104 VSS N12LL L=6E-08 W=1E-06
M81 57 CLKX 79 VSS N12LL L=6E-08 W=5E-07
M82 4 6 VSS VSS N12LL L=6E-08 W=5E-07
M83 VSS 87 105 VSS N12LL L=6E-08 W=1E-06
M84 VSS 79 58 VSS N12LL L=6E-08 W=4E-07
M85 YCKX 58 YX[7] VSS N12LL L=6E-08 W=1.25E-06
M86 VSS 6 4 VSS N12LL L=6E-08 W=5E-07
M87 106 87 VSS VSS N12LL L=6E-08 W=1E-06
M88 59 81 VSS VSS N12LL L=6E-08 W=4E-07
M89 YX[5] 59 YCKX VSS N12LL L=6E-08 W=1.25E-06
M90 81 59 VSS VSS N12LL L=6E-07 W=1.2E-07
M91 81 CLKX 60 VSS N12LL L=6E-08 W=5E-07
M92 107 5 106 VSS N12LL L=6E-08 W=1E-06
M93 VSS 81 59 VSS N12LL L=6E-08 W=4E-07
M94 YCKX 59 YX[5] VSS N12LL L=6E-08 W=1.25E-06
M95 60 CLKX 81 VSS N12LL L=6E-08 W=5E-07
M96 60 4 107 VSS N12LL L=6E-08 W=1E-06
M97 59 81 VSS VSS N12LL L=6E-08 W=4E-07
M98 YX[5] 59 YCKX VSS N12LL L=6E-08 W=1.25E-06
M99 81 CLKX 60 VSS N12LL L=6E-08 W=5E-07
M100 108 VDD VSS VSS N12LL L=3E-07 W=4E-07
M101 VSS 81 59 VSS N12LL L=6E-08 W=4E-07
M102 YCKX 59 YX[5] VSS N12LL L=6E-08 W=1.25E-06
M103 62 83 VSS VSS N12LL L=6E-08 W=4E-07
M104 YX[4] 62 YCKX VSS N12LL L=6E-08 W=1.25E-06
M105 85 A[0] 108 VSS N12LL L=6E-08 W=4E-07
M106 61 CLKX 83 VSS N12LL L=6E-08 W=5E-07
M107 VSS 62 83 VSS N12LL L=6E-07 W=1.2E-07
M108 VSS 83 62 VSS N12LL L=6E-08 W=4E-07
M109 YCKX 62 YX[4] VSS N12LL L=6E-08 W=1.25E-06
M110 109 4 61 VSS N12LL L=6E-08 W=1E-06
M111 83 CLKX 61 VSS N12LL L=6E-08 W=5E-07
M112 62 83 VSS VSS N12LL L=6E-08 W=4E-07
M113 YX[4] 62 YCKX VSS N12LL L=6E-08 W=1.25E-06
M114 110 88 109 VSS N12LL L=6E-08 W=1E-06
M115 61 CLKX 83 VSS N12LL L=6E-08 W=5E-07
M116 5 85 VSS VSS N12LL L=6E-08 W=5E-07
M117 VSS 87 110 VSS N12LL L=6E-08 W=1E-06
M118 VSS 83 62 VSS N12LL L=6E-08 W=4E-07
M119 YCKX 62 YX[4] VSS N12LL L=6E-08 W=1.25E-06
M120 VSS 85 5 VSS N12LL L=6E-08 W=5E-07
M121 111 87 VSS VSS N12LL L=6E-08 W=1E-06
M122 63 89 VSS VSS N12LL L=6E-08 W=4E-07
M123 YX[6] 63 YCKX VSS N12LL L=6E-08 W=1.25E-06
M124 89 63 VSS VSS N12LL L=6E-07 W=1.2E-07
M125 89 CLKX 90 VSS N12LL L=6E-08 W=5E-07
M126 88 5 VSS VSS N12LL L=6E-08 W=5E-07
M127 112 88 111 VSS N12LL L=6E-08 W=1E-06
M128 VSS 89 63 VSS N12LL L=6E-08 W=4E-07
M129 YCKX 63 YX[6] VSS N12LL L=6E-08 W=1.25E-06
M130 90 CLKX 89 VSS N12LL L=6E-08 W=5E-07
M131 90 6 112 VSS N12LL L=6E-08 W=1E-06
M132 VSS 5 88 VSS N12LL L=6E-08 W=5E-07
M133 63 89 VSS VSS N12LL L=6E-08 W=4E-07
M134 YX[6] 63 YCKX VSS N12LL L=6E-08 W=1.25E-06
M135 89 CLKX 90 VSS N12LL L=6E-08 W=5E-07
M136 VSS 89 63 VSS N12LL L=6E-08 W=4E-07
M137 YCKX 63 YX[6] VSS N12LL L=6E-08 W=1.25E-06
M138 51 64 VDD VDD P12LL L=6E-08 W=4E-07
M139 YX[3] 64 YCKX VDD P12LL L=6E-08 W=1.25E-06
M140 YX[3] 51 VDD VDD P12LL L=6E-08 W=1.25E-06
M141 65 CLK 64 VDD P12LL L=6E-08 W=5E-07
M142 VDD 6 65 VDD P12LL L=6E-08 W=1E-06
M143 VDD 64 51 VDD P12LL L=6E-08 W=4E-07
M144 YCKX 64 YX[3] VDD P12LL L=6E-08 W=1.25E-06
M145 VDD 51 YX[3] VDD P12LL L=6E-08 W=1.25E-06
M146 64 CLK 65 VDD P12LL L=6E-08 W=5E-07
M147 VDD 51 64 VDD P12LL L=3E-07 W=1.2E-07
M148 65 5 VDD VDD P12LL L=6E-08 W=1E-06
M149 51 64 VDD VDD P12LL L=6E-08 W=4E-07
M150 YX[3] 64 YCKX VDD P12LL L=6E-08 W=1.25E-06
M151 YX[3] 51 VDD VDD P12LL L=6E-08 W=1.25E-06
M152 65 CLK 64 VDD P12LL L=6E-08 W=5E-07
M153 73 87 VDD VDD P12LL L=6E-08 W=1E-06
M154 VDD 73 65 VDD P12LL L=6E-08 W=1E-06
M155 VDD 64 51 VDD P12LL L=6E-08 W=4E-07
M156 YCKX 64 YX[3] VDD P12LL L=6E-08 W=1.25E-06
M157 VDD 51 YX[3] VDD P12LL L=6E-08 W=1.25E-06
M158 VDD 87 73 VDD P12LL L=6E-08 W=1E-06
M159 53 73 VDD VDD P12LL L=6E-08 W=1E-06
M160 52 67 VDD VDD P12LL L=6E-08 W=4E-07
M161 YX[1] 67 YCKX VDD P12LL L=6E-08 W=1.25E-06
M162 YX[1] 52 VDD VDD P12LL L=6E-08 W=1.25E-06
M163 67 52 VDD VDD P12LL L=3E-07 W=1.2E-07
M164 67 CLK 53 VDD P12LL L=6E-08 W=5E-07
M165 87 69 VDD VDD P12LL L=6E-08 W=1E-06
M166 VDD 5 53 VDD P12LL L=6E-08 W=1E-06
M167 VDD 67 52 VDD P12LL L=6E-08 W=4E-07
M168 YCKX 67 YX[1] VDD P12LL L=6E-08 W=1.25E-06
M169 VDD 52 YX[1] VDD P12LL L=6E-08 W=1.25E-06
M170 53 CLK 67 VDD P12LL L=6E-08 W=5E-07
M171 VDD 69 87 VDD P12LL L=6E-08 W=1E-06
M172 53 4 VDD VDD P12LL L=6E-08 W=1E-06
M173 52 67 VDD VDD P12LL L=6E-08 W=4E-07
M174 YX[1] 67 YCKX VDD P12LL L=6E-08 W=1.25E-06
M175 YX[1] 52 VDD VDD P12LL L=6E-08 W=1.25E-06
M176 67 CLK 53 VDD P12LL L=6E-08 W=5E-07
M177 VDD 67 52 VDD P12LL L=6E-08 W=4E-07
M178 YCKX 67 YX[1] VDD P12LL L=6E-08 W=1.25E-06
M179 VDD 52 YX[1] VDD P12LL L=6E-08 W=1.25E-06
M180 113 A[2] 69 VDD P12LL L=6E-08 W=4E-07
M181 55 71 VDD VDD P12LL L=6E-08 W=4E-07
M182 YX[0] 71 YCKX VDD P12LL L=6E-08 W=1.25E-06
M183 YX[0] 55 VDD VDD P12LL L=6E-08 W=1.25E-06
M184 54 CLK 71 VDD P12LL L=6E-08 W=5E-07
M185 VDD VSS 113 VDD P12LL L=1E-07 W=4E-07
M186 VDD 4 54 VDD P12LL L=6E-08 W=1E-06
M187 VDD 71 55 VDD P12LL L=6E-08 W=4E-07
M188 YCKX 71 YX[0] VDD P12LL L=6E-08 W=1.25E-06
M189 VDD 55 YX[0] VDD P12LL L=6E-08 W=1.25E-06
M190 71 CLK 54 VDD P12LL L=6E-08 W=5E-07
M191 VDD 55 71 VDD P12LL L=3E-07 W=1.2E-07
M192 54 88 VDD VDD P12LL L=6E-08 W=1E-06
M193 55 71 VDD VDD P12LL L=6E-08 W=4E-07
M194 YX[0] 71 YCKX VDD P12LL L=6E-08 W=1.25E-06
M195 YX[0] 55 VDD VDD P12LL L=6E-08 W=1.25E-06
M196 54 CLK 71 VDD P12LL L=6E-08 W=5E-07
M197 VDD 73 54 VDD P12LL L=6E-08 W=1E-06
M198 VDD 71 55 VDD P12LL L=6E-08 W=4E-07
M199 YCKX 71 YX[0] VDD P12LL L=6E-08 W=1.25E-06
M200 VDD 55 YX[0] VDD P12LL L=6E-08 W=1.25E-06
M201 75 73 VDD VDD P12LL L=6E-08 W=1E-06
M202 56 74 VDD VDD P12LL L=6E-08 W=4E-07
M203 YX[2] 74 YCKX VDD P12LL L=6E-08 W=1.25E-06
M204 YX[2] 56 VDD VDD P12LL L=6E-08 W=1.25E-06
M205 74 56 VDD VDD P12LL L=3E-07 W=1.2E-07
M206 74 CLK 75 VDD P12LL L=6E-08 W=5E-07
M207 114 VSS VDD VDD P12LL L=1E-07 W=4E-07
M208 VDD 88 75 VDD P12LL L=6E-08 W=1E-06
M209 VDD 74 56 VDD P12LL L=6E-08 W=4E-07
M210 YCKX 74 YX[2] VDD P12LL L=6E-08 W=1.25E-06
M211 VDD 56 YX[2] VDD P12LL L=6E-08 W=1.25E-06
M212 75 CLK 74 VDD P12LL L=6E-08 W=5E-07
M213 75 6 VDD VDD P12LL L=6E-08 W=1E-06
M214 56 74 VDD VDD P12LL L=6E-08 W=4E-07
M215 YX[2] 74 YCKX VDD P12LL L=6E-08 W=1.25E-06
M216 YX[2] 56 VDD VDD P12LL L=6E-08 W=1.25E-06
M217 74 CLK 75 VDD P12LL L=6E-08 W=5E-07
M218 78 A[1] 114 VDD P12LL L=6E-08 W=4E-07
M219 VDD 74 56 VDD P12LL L=6E-08 W=4E-07
M220 YCKX 74 YX[2] VDD P12LL L=6E-08 W=1.25E-06
M221 VDD 56 YX[2] VDD P12LL L=6E-08 W=1.25E-06
M222 58 79 VDD VDD P12LL L=6E-08 W=4E-07
M223 YX[7] 79 YCKX VDD P12LL L=6E-08 W=1.25E-06
M224 YX[7] 58 VDD VDD P12LL L=6E-08 W=1.25E-06
M225 57 CLK 79 VDD P12LL L=6E-08 W=5E-07
M226 6 78 VDD VDD P12LL L=6E-08 W=1E-06
M227 VDD 6 57 VDD P12LL L=6E-08 W=1E-06
M228 VDD 79 58 VDD P12LL L=6E-08 W=4E-07
M229 YCKX 79 YX[7] VDD P12LL L=6E-08 W=1.25E-06
M230 VDD 58 YX[7] VDD P12LL L=6E-08 W=1.25E-06
M231 79 CLK 57 VDD P12LL L=6E-08 W=5E-07
M232 VDD 78 6 VDD P12LL L=6E-08 W=1E-06
M233 VDD 58 79 VDD P12LL L=3E-07 W=1.2E-07
M234 57 5 VDD VDD P12LL L=6E-08 W=1E-06
M235 58 79 VDD VDD P12LL L=6E-08 W=4E-07
M236 YX[7] 79 YCKX VDD P12LL L=6E-08 W=1.25E-06
M237 YX[7] 58 VDD VDD P12LL L=6E-08 W=1.25E-06
M238 57 CLK 79 VDD P12LL L=6E-08 W=5E-07
M239 4 6 VDD VDD P12LL L=6E-08 W=1E-06
M240 VDD 87 57 VDD P12LL L=6E-08 W=1E-06
M241 VDD 79 58 VDD P12LL L=6E-08 W=4E-07
M242 YCKX 79 YX[7] VDD P12LL L=6E-08 W=1.25E-06
M243 VDD 58 YX[7] VDD P12LL L=6E-08 W=1.25E-06
M244 VDD 6 4 VDD P12LL L=6E-08 W=1E-06
M245 60 87 VDD VDD P12LL L=6E-08 W=1E-06
M246 59 81 VDD VDD P12LL L=6E-08 W=4E-07
M247 YX[5] 81 YCKX VDD P12LL L=6E-08 W=1.25E-06
M248 YX[5] 59 VDD VDD P12LL L=6E-08 W=1.25E-06
M249 81 59 VDD VDD P12LL L=3E-07 W=1.2E-07
M250 81 CLK 60 VDD P12LL L=6E-08 W=5E-07
M251 VDD 5 60 VDD P12LL L=6E-08 W=1E-06
M252 VDD 81 59 VDD P12LL L=6E-08 W=4E-07
M253 YCKX 81 YX[5] VDD P12LL L=6E-08 W=1.25E-06
M254 VDD 59 YX[5] VDD P12LL L=6E-08 W=1.25E-06
M255 60 CLK 81 VDD P12LL L=6E-08 W=5E-07
M256 60 4 VDD VDD P12LL L=6E-08 W=1E-06
M257 59 81 VDD VDD P12LL L=6E-08 W=4E-07
M258 YX[5] 81 YCKX VDD P12LL L=6E-08 W=1.25E-06
M259 YX[5] 59 VDD VDD P12LL L=6E-08 W=1.25E-06
M260 81 CLK 60 VDD P12LL L=6E-08 W=5E-07
M261 115 VSS VDD VDD P12LL L=1E-07 W=4E-07
M262 VDD 81 59 VDD P12LL L=6E-08 W=4E-07
M263 YCKX 81 YX[5] VDD P12LL L=6E-08 W=1.25E-06
M264 VDD 59 YX[5] VDD P12LL L=6E-08 W=1.25E-06
M265 62 83 VDD VDD P12LL L=6E-08 W=4E-07
M266 YX[4] 83 YCKX VDD P12LL L=6E-08 W=1.25E-06
M267 YX[4] 62 VDD VDD P12LL L=6E-08 W=1.25E-06
M268 85 A[0] 115 VDD P12LL L=6E-08 W=4E-07
M269 61 CLK 83 VDD P12LL L=6E-08 W=5E-07
M270 VDD 4 61 VDD P12LL L=6E-08 W=1E-06
M271 VDD 83 62 VDD P12LL L=6E-08 W=4E-07
M272 YCKX 83 YX[4] VDD P12LL L=6E-08 W=1.25E-06
M273 VDD 62 YX[4] VDD P12LL L=6E-08 W=1.25E-06
M274 83 CLK 61 VDD P12LL L=6E-08 W=5E-07
M275 VDD 62 83 VDD P12LL L=3E-07 W=1.2E-07
M276 61 88 VDD VDD P12LL L=6E-08 W=1E-06
M277 62 83 VDD VDD P12LL L=6E-08 W=4E-07
M278 YX[4] 83 YCKX VDD P12LL L=6E-08 W=1.25E-06
M279 YX[4] 62 VDD VDD P12LL L=6E-08 W=1.25E-06
M280 61 CLK 83 VDD P12LL L=6E-08 W=5E-07
M281 5 85 VDD VDD P12LL L=6E-08 W=1E-06
M282 VDD 87 61 VDD P12LL L=6E-08 W=1E-06
M283 VDD 83 62 VDD P12LL L=6E-08 W=4E-07
M284 YCKX 83 YX[4] VDD P12LL L=6E-08 W=1.25E-06
M285 VDD 62 YX[4] VDD P12LL L=6E-08 W=1.25E-06
M286 VDD 85 5 VDD P12LL L=6E-08 W=1E-06
M287 90 87 VDD VDD P12LL L=6E-08 W=1E-06
M288 63 89 VDD VDD P12LL L=6E-08 W=4E-07
M289 YX[6] 89 YCKX VDD P12LL L=6E-08 W=1.25E-06
M290 YX[6] 63 VDD VDD P12LL L=6E-08 W=1.25E-06
M291 89 63 VDD VDD P12LL L=3E-07 W=1.2E-07
M292 89 CLK 90 VDD P12LL L=6E-08 W=5E-07
M293 88 5 VDD VDD P12LL L=6E-08 W=1E-06
M294 VDD 88 90 VDD P12LL L=6E-08 W=1E-06
M295 VDD 89 63 VDD P12LL L=6E-08 W=4E-07
M296 YCKX 89 YX[6] VDD P12LL L=6E-08 W=1.25E-06
M297 VDD 63 YX[6] VDD P12LL L=6E-08 W=1.25E-06
M298 90 CLK 89 VDD P12LL L=6E-08 W=5E-07
M299 VDD 5 88 VDD P12LL L=6E-08 W=1E-06
M300 90 6 VDD VDD P12LL L=6E-08 W=1E-06
M301 63 89 VDD VDD P12LL L=6E-08 W=4E-07
M302 YX[6] 89 YCKX VDD P12LL L=6E-08 W=1.25E-06
M303 YX[6] 63 VDD VDD P12LL L=6E-08 W=1.25E-06
M304 89 CLK 90 VDD P12LL L=6E-08 W=5E-07
M305 VDD 89 63 VDD P12LL L=6E-08 W=4E-07
M306 YCKX 89 YX[6] VDD P12LL L=6E-08 W=1.25E-06
M307 VDD 63 YX[6] VDD P12LL L=6E-08 W=1.25E-06
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    S55NLLGDPH_X512Y8D16_BW_LOGIC_BASE
* View Name:    schematic
************************************************************************

.SUBCKT S55NLLGDPH_X512Y8D16_BW_LOGIC_BASE ACTRCLK ACTRCLKX DCTRCLK DCTRCLKX EMCLK FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3]
+FCKX[2] FCKX[1] FCKX[0] PXA[3] PXA[2] PXA[1] PXA[0] RWL SACK1 SACK4
+WE A[4] A[3] A[2] A[1] A[0] CEN CLK FB RDE
+WEN INTCLKX S[1] S[0] VDD VSS
M0 4 7 INTCLKX VSS N12LL L=6E-08 W=5E-07 $X=5365 $Y=27535 $D=0
M1 RWL 4 VSS VSS N12LL L=6E-08 W=1E-06 $X=5365 $Y=28740 $D=0
M2 VSS 11 6 VSS N12LL L=6E-08 W=4E-07 $X=5565 $Y=15355 $D=0
M3 6 ACTRCLKX 13 VSS N12LL L=6E-08 W=5E-07 $X=5565 $Y=16300 $D=0
M4 VSS 13 12 VSS N12LL L=6E-08 W=4E-07 $X=5565 $Y=20640 $D=0
M5 INTCLKX 7 4 VSS N12LL L=6E-08 W=5E-07 $X=5655 $Y=27535 $D=0
M6 VSS 4 RWL VSS N12LL L=6E-08 W=1E-06 $X=5655 $Y=28740 $D=0
M7 525 VDD VSS VSS N12LL L=3E-07 W=4E-07 $X=5665 $Y=11140 $D=0
M8 13 ACTRCLKX 6 VSS N12LL L=6E-08 W=5E-07 $X=5835 $Y=16300 $D=0
M9 VSS S[0] 8 VSS N12LL L=6E-08 W=4E-07 $X=5850 $Y=6115 $D=0
M10 VSS S[1] 9 VSS N12LL L=6E-08 W=4E-07 $X=5850 $Y=7145 $D=0
M11 4 7 INTCLKX VSS N12LL L=6E-08 W=5E-07 $X=5925 $Y=27535 $D=0
M12 RWL 4 VSS VSS N12LL L=6E-08 W=1E-06 $X=5945 $Y=28740 $D=0
M13 13 12 VSS VSS N12LL L=6E-07 W=1.2E-07 $X=6025 $Y=20875 $D=0
M14 7 12 VSS VSS N12LL L=6E-08 W=4E-07 $X=6035 $Y=22125 $D=0
M15 23 8 VSS VSS N12LL L=6E-08 W=4E-07 $X=6120 $Y=6115 $D=0
M16 16 9 VSS VSS N12LL L=6E-08 W=4E-07 $X=6120 $Y=7145 $D=0
M17 VSS 19 11 VSS N12LL L=6E-08 W=4E-07 $X=6155 $Y=15355 $D=0
M18 INTCLKX 7 4 VSS N12LL L=6E-08 W=5E-07 $X=6215 $Y=27535 $D=0
M19 17 RDE 525 VSS N12LL L=6E-08 W=4E-07 $X=6230 $Y=11140 $D=0
M20 VSS 4 RWL VSS N12LL L=6E-08 W=1E-06 $X=6235 $Y=28740 $D=0
M21 19 17 VSS VSS N12LL L=6E-08 W=4E-07 $X=6425 $Y=15355 $D=0
M22 529 9 21 VSS N12LL L=6E-08 W=4E-07 $X=6720 $Y=6115 $D=0
M23 530 9 22 VSS N12LL L=6E-08 W=4E-07 $X=6720 $Y=7145 $D=0
M24 VSS 8 529 VSS N12LL L=6E-08 W=4E-07 $X=6990 $Y=6115 $D=0
M25 VSS 23 530 VSS N12LL L=6E-08 W=4E-07 $X=6990 $Y=7145 $D=0
M26 532 8 VSS VSS N12LL L=6E-08 W=4E-07 $X=7260 $Y=6115 $D=0
M27 533 23 VSS VSS N12LL L=6E-08 W=4E-07 $X=7260 $Y=7145 $D=0
M28 24 16 532 VSS N12LL L=6E-08 W=4E-07 $X=7530 $Y=6115 $D=0
M29 25 16 533 VSS N12LL L=6E-08 W=4E-07 $X=7530 $Y=7145 $D=0
M30 46 30 VSS VSS N12LL L=6E-08 W=5E-07 $X=7565 $Y=15325 $D=0
M31 PXA[3] 29 VSS VSS N12LL L=6E-08 W=1.5E-06 $X=7810 $Y=28665 $D=0
M32 VSS RDE 46 VSS N12LL L=6E-08 W=5E-07 $X=7855 $Y=15325 $D=0
M33 36 PXA[2] VSS VSS N12LL L=6E-07 W=1.2E-07 $X=7890 $Y=27880 $D=0
M34 535 46 27 VSS N12LL L=6E-08 W=1.5E-06 $X=7920 $Y=16875 $D=0
M35 VSS A[3] 30 VSS N12LL L=6E-08 W=4E-07 $X=7950 $Y=11140 $D=0
M36 29 ACTRCLKX 27 VSS N12LL L=6E-08 W=2.5E-06 $X=7955 $Y=21115 $D=0
M37 40 45 VSS VSS N12LL L=6E-08 W=5E-07 $X=8010 $Y=1910 $D=0
M38 VSS PXA[3] 29 VSS N12LL L=6E-07 W=1.2E-07 $X=8060 $Y=27195 $D=0
M39 VSS 29 PXA[3] VSS N12LL L=6E-08 W=1.5E-06 $X=8100 $Y=28665 $D=0
M40 VSS 42 535 VSS N12LL L=6E-08 W=1.5E-06 $X=8110 $Y=16875 $D=0
M41 32 RDE VSS VSS N12LL L=6E-08 W=7E-07 $X=8145 $Y=15325 $D=0
M42 VSS 45 40 VSS N12LL L=6E-08 W=5E-07 $X=8280 $Y=1910 $D=0
M43 VSS 25 37 VSS N12LL L=6E-08 W=4E-07 $X=8280 $Y=8585 $D=0
M44 31 30 VSS VSS N12LL L=6E-08 W=4E-07 $X=8280 $Y=11140 $D=0
M45 537 42 VSS VSS N12LL L=6E-08 W=1.5E-06 $X=8380 $Y=16875 $D=0
M46 PXA[2] 36 VSS VSS N12LL L=6E-08 W=1.5E-06 $X=8390 $Y=28665 $D=0
M47 VSS 31 32 VSS N12LL L=6E-08 W=7E-07 $X=8435 $Y=15325 $D=0
M48 34 ACTRCLKX 36 VSS N12LL L=6E-08 W=2.5E-06 $X=8535 $Y=21115 $D=0
M49 34 32 537 VSS N12LL L=6E-08 W=1.5E-06 $X=8570 $Y=16875 $D=0
M50 EMCLK 37 40 VSS N12LL L=6E-08 W=1E-06 $X=8630 $Y=7220 $D=0
M51 VSS 36 PXA[2] VSS N12LL L=6E-08 W=1.5E-06 $X=8680 $Y=28665 $D=0
M52 40 37 EMCLK VSS N12LL L=6E-08 W=1.5E-06 $X=8900 $Y=7220 $D=0
M53 PXA[0] 38 VSS VSS N12LL L=6E-08 W=1.5E-06 $X=9020 $Y=28665 $D=0
M54 48 PXA[1] VSS VSS N12LL L=6E-07 W=1.2E-07 $X=9100 $Y=27195 $D=0
M55 539 32 41 VSS N12LL L=6E-08 W=1.5E-06 $X=9130 $Y=16875 $D=0
M56 38 ACTRCLKX 41 VSS N12LL L=6E-08 W=2.5E-06 $X=9165 $Y=21115 $D=0
M57 540 VDD VSS VSS N12LL L=3E-07 W=4E-07 $X=9205 $Y=11140 $D=0
M58 VSS 45 40 VSS N12LL L=6E-08 W=1.5E-06 $X=9215 $Y=7220 $D=0
M59 VSS 49 42 VSS N12LL L=6E-08 W=7E-07 $X=9265 $Y=15325 $D=0
M60 VSS PXA[0] 38 VSS N12LL L=6E-07 W=1.2E-07 $X=9270 $Y=27880 $D=0
M61 VSS 38 PXA[0] VSS N12LL L=6E-08 W=1.5E-06 $X=9310 $Y=28665 $D=0
M62 VSS 47 539 VSS N12LL L=6E-08 W=1.5E-06 $X=9320 $Y=16875 $D=0
M63 45 102 VSS VSS N12LL L=6E-08 W=7.5E-07 $X=9515 $Y=7220 $D=0
M64 47 42 VSS VSS N12LL L=6E-08 W=7E-07 $X=9555 $Y=15325 $D=0
M65 542 47 VSS VSS N12LL L=6E-08 W=1.5E-06 $X=9590 $Y=16875 $D=0
M66 PXA[1] 48 VSS VSS N12LL L=6E-08 W=1.5E-06 $X=9600 $Y=28665 $D=0
M67 50 ACTRCLKX 48 VSS N12LL L=6E-08 W=2.5E-06 $X=9745 $Y=21115 $D=0
M68 49 A[4] 540 VSS N12LL L=6E-08 W=4E-07 $X=9770 $Y=11140 $D=0
M69 50 46 542 VSS N12LL L=6E-08 W=1.5E-06 $X=9780 $Y=16875 $D=0
M70 VSS 48 PXA[1] VSS N12LL L=6E-08 W=1.5E-06 $X=9890 $Y=28665 $D=0
M71 VSS FB 52 VSS N12LL L=6E-08 W=8E-07 $X=10135 $Y=7215 $D=0
M72 80 52 VSS VSS N12LL L=6E-08 W=1.25E-06 $X=10495 $Y=7215 $D=0
M73 VSS 52 80 VSS N12LL L=6E-08 W=1.25E-06 $X=10765 $Y=7215 $D=0
M74 VSS 40 55 VSS N12LL L=3E-07 W=7E-07 $X=10815 $Y=9090 $D=0
M75 VSS 24 53 VSS N12LL L=6E-08 W=4E-07 $X=10890 $Y=15230 $D=0
M76 54 55 VSS VSS N12LL L=6E-08 W=6.25E-07 $X=11115 $Y=7470 $D=0
M77 62 22 VSS VSS N12LL L=6E-08 W=4E-07 $X=11160 $Y=15230 $D=0
M78 54 55 VSS VSS N12LL L=6E-08 W=1.25E-06 $X=11385 $Y=8540 $D=0
M79 VSS 55 54 VSS N12LL L=6E-08 W=6.25E-07 $X=11410 $Y=7470 $D=0
M80 59 57 VSS VSS N12LL L=6E-08 W=4E-07 $X=11485 $Y=29110 $D=0
M81 FCKX[3] 59 INTCLKX VSS N12LL L=6E-08 W=1.25E-06 $X=11485 $Y=33030 $D=0
M82 60 ACTRCLKX 57 VSS N12LL L=6E-08 W=5E-07 $X=11645 $Y=25070 $D=0
M83 EMCLK 53 54 VSS N12LL L=6E-08 W=1.25E-06 $X=11715 $Y=8540 $D=0
M84 VSS 59 57 VSS N12LL L=6E-07 W=1.2E-07 $X=11735 $Y=30405 $D=0
M85 67 21 VSS VSS N12LL L=6E-08 W=4E-07 $X=11760 $Y=14620 $D=0
M86 VSS 57 59 VSS N12LL L=6E-08 W=4E-07 $X=11775 $Y=29110 $D=0
M87 INTCLKX 59 FCKX[3] VSS N12LL L=6E-08 W=1.25E-06 $X=11775 $Y=33030 $D=0
M88 548 58 60 VSS N12LL L=6E-08 W=1E-06 $X=11875 $Y=23525 $D=0
M89 57 ACTRCLKX 60 VSS N12LL L=6E-08 W=5E-07 $X=11915 $Y=25070 $D=0
M90 54 53 EMCLK VSS N12LL L=6E-08 W=1.25E-06 $X=11985 $Y=8540 $D=0
M91 VSS 66 65 VSS N12LL L=3E-07 W=7E-07 $X=12010 $Y=15390 $D=0
M92 59 57 VSS VSS N12LL L=6E-08 W=4E-07 $X=12065 $Y=29110 $D=0
M93 FCKX[3] 59 INTCLKX VSS N12LL L=6E-08 W=1.25E-06 $X=12065 $Y=33030 $D=0
M94 551 63 548 VSS N12LL L=6E-08 W=1E-06 $X=12115 $Y=23525 $D=0
M95 60 ACTRCLKX 57 VSS N12LL L=6E-08 W=5E-07 $X=12195 $Y=25070 $D=0
M96 VSS 65 77 VSS N12LL L=6E-08 W=6.25E-07 $X=12230 $Y=16900 $D=0
M97 84 118 VSS VSS N12LL L=6E-08 W=5E-07 $X=12265 $Y=19040 $D=0
M98 VSS CLK 64 VSS N12LL L=6E-08 W=4E-07 $X=12330 $Y=6620 $D=0
M99 VSS 84 551 VSS N12LL L=6E-08 W=1E-06 $X=12355 $Y=23525 $D=0
M100 VSS 57 59 VSS N12LL L=6E-08 W=4E-07 $X=12355 $Y=29110 $D=0
M101 INTCLKX 59 FCKX[3] VSS N12LL L=6E-08 W=1.25E-06 $X=12355 $Y=33030 $D=0
M102 77 65 VSS VSS N12LL L=6E-08 W=1.25E-06 $X=12530 $Y=15390 $D=0
M103 77 65 VSS VSS N12LL L=6E-08 W=6.25E-07 $X=12530 $Y=16900 $D=0
M104 VSS 118 84 VSS N12LL L=6E-08 W=5E-07 $X=12555 $Y=19040 $D=0
M105 EMCLK 62 66 VSS N12LL L=6E-08 W=1.25E-06 $X=12595 $Y=8540 $D=0
M106 554 84 VSS VSS N12LL L=6E-08 W=1E-06 $X=12645 $Y=23525 $D=0
M107 68 70 VSS VSS N12LL L=6E-08 W=4E-07 $X=12645 $Y=29110 $D=0
M108 FCKX[1] 68 INTCLKX VSS N12LL L=6E-08 W=1.25E-06 $X=12645 $Y=33030 $D=0
M109 555 64 VSS VSS N12LL L=6E-08 W=1E-06 $X=12670 $Y=6620 $D=0
M110 70 68 VSS VSS N12LL L=6E-07 W=1.2E-07 $X=12725 $Y=30405 $D=0
M111 70 ACTRCLKX 69 VSS N12LL L=6E-08 W=5E-07 $X=12805 $Y=25070 $D=0
M112 118 75 VSS VSS N12LL L=6E-08 W=5E-07 $X=12845 $Y=19040 $D=0
M113 EMCLK 67 77 VSS N12LL L=6E-08 W=1.25E-06 $X=12860 $Y=15390 $D=0
M114 66 62 EMCLK VSS N12LL L=6E-08 W=1.25E-06 $X=12865 $Y=8540 $D=0
M115 557 63 554 VSS N12LL L=6E-08 W=1E-06 $X=12885 $Y=23525 $D=0
M116 78 CEN 555 VSS N12LL L=6E-08 W=1E-06 $X=12910 $Y=6620 $D=0
M117 VSS 70 68 VSS N12LL L=6E-08 W=4E-07 $X=12935 $Y=29110 $D=0
M118 INTCLKX 68 FCKX[1] VSS N12LL L=6E-08 W=1.25E-06 $X=12935 $Y=33030 $D=0
M119 69 ACTRCLKX 70 VSS N12LL L=6E-08 W=5E-07 $X=13085 $Y=25070 $D=0
M120 69 74 557 VSS N12LL L=6E-08 W=1E-06 $X=13125 $Y=23525 $D=0
M121 77 67 EMCLK VSS N12LL L=6E-08 W=1.25E-06 $X=13130 $Y=15390 $D=0
M122 VSS 75 118 VSS N12LL L=6E-08 W=5E-07 $X=13135 $Y=19040 $D=0
M123 VSS 79 66 VSS N12LL L=6E-08 W=1.25E-06 $X=13155 $Y=8540 $D=0
M124 68 70 VSS VSS N12LL L=6E-08 W=4E-07 $X=13225 $Y=29110 $D=0
M125 FCKX[1] 68 INTCLKX VSS N12LL L=6E-08 W=1.25E-06 $X=13225 $Y=33030 $D=0
M126 VSS 85 78 VSS N12LL L=6E-07 W=1.2E-07 $X=13270 $Y=6620 $D=0
M127 70 ACTRCLKX 69 VSS N12LL L=6E-08 W=5E-07 $X=13355 $Y=25070 $D=0
M128 79 54 VSS VSS N12LL L=3E-07 W=7E-07 $X=13485 $Y=9090 $D=0
M129 VSS 70 68 VSS N12LL L=6E-08 W=4E-07 $X=13515 $Y=29110 $D=0
M130 INTCLKX 68 FCKX[1] VSS N12LL L=6E-08 W=1.25E-06 $X=13515 $Y=33030 $D=0
M131 VSS 79 66 VSS N12LL L=6E-08 W=6.25E-07 $X=13735 $Y=8005 $D=0
M132 560 A[2] 75 VSS N12LL L=6E-08 W=4E-07 $X=13765 $Y=19085 $D=0
M133 VSS 86 106 VSS N12LL L=6E-08 W=2.5E-06 $X=13770 $Y=14750 $D=0
M134 81 76 VSS VSS N12LL L=6E-08 W=4E-07 $X=13805 $Y=29110 $D=0
M135 FCKX[0] 81 INTCLKX VSS N12LL L=6E-08 W=1.25E-06 $X=13805 $Y=33030 $D=0
M136 82 ACTRCLKX 76 VSS N12LL L=6E-08 W=5E-07 $X=13965 $Y=25070 $D=0
M137 66 79 VSS VSS N12LL L=6E-08 W=6.25E-07 $X=14035 $Y=8005 $D=0
M138 106 86 VSS VSS N12LL L=6E-08 W=2.5E-06 $X=14040 $Y=14750 $D=0
M139 VSS VDD 560 VSS N12LL L=3E-07 W=4E-07 $X=14045 $Y=19085 $D=0
M140 VSS 81 76 VSS N12LL L=6E-07 W=1.2E-07 $X=14055 $Y=30405 $D=0
M141 VSS 76 81 VSS N12LL L=6E-08 W=4E-07 $X=14095 $Y=29110 $D=0
M142 INTCLKX 81 FCKX[0] VSS N12LL L=6E-08 W=1.25E-06 $X=14095 $Y=33030 $D=0
M143 562 74 82 VSS N12LL L=6E-08 W=1E-06 $X=14195 $Y=23525 $D=0
M144 85 78 VSS VSS N12LL L=6E-08 W=4E-07 $X=14200 $Y=6620 $D=0
M145 76 ACTRCLKX 82 VSS N12LL L=6E-08 W=5E-07 $X=14235 $Y=25070 $D=0
M146 VSS 86 106 VSS N12LL L=6E-08 W=2.5E-06 $X=14310 $Y=14750 $D=0
M147 81 76 VSS VSS N12LL L=6E-08 W=4E-07 $X=14385 $Y=29110 $D=0
M148 FCKX[0] 81 INTCLKX VSS N12LL L=6E-08 W=1.25E-06 $X=14385 $Y=33030 $D=0
M149 563 121 562 VSS N12LL L=6E-08 W=1E-06 $X=14435 $Y=23525 $D=0
M150 82 ACTRCLKX 76 VSS N12LL L=6E-08 W=5E-07 $X=14515 $Y=25070 $D=0
M151 106 86 VSS VSS N12LL L=6E-08 W=2.5E-06 $X=14580 $Y=14750 $D=0
M152 VSS 84 563 VSS N12LL L=6E-08 W=1E-06 $X=14675 $Y=23525 $D=0
M153 VSS 76 81 VSS N12LL L=6E-08 W=4E-07 $X=14675 $Y=29110 $D=0
M154 INTCLKX 81 FCKX[0] VSS N12LL L=6E-08 W=1.25E-06 $X=14675 $Y=33030 $D=0
M155 VSS 116 102 VSS N12LL L=1E-06 W=1.2E-07 $X=14795 $Y=8155 $D=0
M156 VSS 86 106 VSS N12LL L=6E-08 W=2.5E-06 $X=14850 $Y=14750 $D=0
M157 87 85 VSS VSS N12LL L=6E-08 W=5E-07 $X=14895 $Y=6520 $D=0
M158 VSS 116 89 VSS N12LL L=3E-07 W=3E-07 $X=14910 $Y=8855 $D=0
M159 566 84 VSS VSS N12LL L=6E-08 W=1E-06 $X=14965 $Y=23525 $D=0
M160 90 91 VSS VSS N12LL L=6E-08 W=4E-07 $X=14965 $Y=29110 $D=0
M161 FCKX[2] 90 INTCLKX VSS N12LL L=6E-08 W=1.25E-06 $X=14965 $Y=33030 $D=0
M162 91 90 VSS VSS N12LL L=6E-07 W=1.2E-07 $X=15045 $Y=30405 $D=0
M163 106 86 VSS VSS N12LL L=6E-08 W=2.5E-06 $X=15120 $Y=14750 $D=0
M164 91 ACTRCLKX 93 VSS N12LL L=6E-08 W=5E-07 $X=15125 $Y=25070 $D=0
M165 VSS CLK 87 VSS N12LL L=6E-08 W=5E-07 $X=15165 $Y=6520 $D=0
M166 569 121 566 VSS N12LL L=6E-08 W=1E-06 $X=15205 $Y=23525 $D=0
M167 570 VDD VSS VSS N12LL L=3E-07 W=4E-07 $X=15225 $Y=19085 $D=0
M168 VSS 91 90 VSS N12LL L=6E-08 W=4E-07 $X=15255 $Y=29110 $D=0
M169 INTCLKX 90 FCKX[2] VSS N12LL L=6E-08 W=1.25E-06 $X=15255 $Y=33030 $D=0
M170 VSS 86 106 VSS N12LL L=6E-08 W=2.5E-06 $X=15390 $Y=14750 $D=0
M171 95 89 VSS VSS N12LL L=2E-07 W=4E-07 $X=15400 $Y=8855 $D=0
M172 93 ACTRCLKX 91 VSS N12LL L=6E-08 W=5E-07 $X=15405 $Y=25070 $D=0
M173 92 87 VSS VSS N12LL L=6E-08 W=5E-07 $X=15435 $Y=6520 $D=0
M174 93 58 569 VSS N12LL L=6E-08 W=1E-06 $X=15445 $Y=23525 $D=0
M175 90 91 VSS VSS N12LL L=6E-08 W=4E-07 $X=15545 $Y=29110 $D=0
M176 FCKX[2] 90 INTCLKX VSS N12LL L=6E-08 W=1.25E-06 $X=15545 $Y=33030 $D=0
M177 106 86 VSS VSS N12LL L=6E-08 W=2.5E-06 $X=15660 $Y=14750 $D=0
M178 91 ACTRCLKX 93 VSS N12LL L=6E-08 W=5E-07 $X=15675 $Y=25070 $D=0
M179 96 A[1] 570 VSS N12LL L=6E-08 W=4E-07 $X=15745 $Y=19085 $D=0
M180 VSS 91 90 VSS N12LL L=6E-08 W=4E-07 $X=15835 $Y=29110 $D=0
M181 INTCLKX 90 FCKX[2] VSS N12LL L=6E-08 W=1.25E-06 $X=15835 $Y=33030 $D=0
M182 102 CLK 106 VSS N12LL L=6E-08 W=2.5E-06 $X=15930 $Y=14750 $D=0
M183 86 92 VSS VSS N12LL L=6E-08 W=5E-07 $X=16045 $Y=6520 $D=0
M184 98 97 VSS VSS N12LL L=6E-08 W=4E-07 $X=16125 $Y=29110 $D=0
M185 FCKX[7] 98 INTCLKX VSS N12LL L=6E-08 W=1.25E-06 $X=16125 $Y=33030 $D=0
M186 106 CLK 102 VSS N12LL L=6E-08 W=2.5E-06 $X=16200 $Y=14750 $D=0
M187 99 ACTRCLKX 97 VSS N12LL L=6E-08 W=5E-07 $X=16285 $Y=25070 $D=0
M188 VSS 92 86 VSS N12LL L=6E-08 W=5E-07 $X=16315 $Y=6520 $D=0
M189 58 96 VSS VSS N12LL L=6E-08 W=5E-07 $X=16375 $Y=19040 $D=0
M190 VSS 98 97 VSS N12LL L=6E-07 W=1.2E-07 $X=16375 $Y=30405 $D=0
M191 VSS 97 98 VSS N12LL L=6E-08 W=4E-07 $X=16415 $Y=29110 $D=0
M192 INTCLKX 98 FCKX[7] VSS N12LL L=6E-08 W=1.25E-06 $X=16415 $Y=33030 $D=0
M193 102 CLK 106 VSS N12LL L=6E-08 W=2.5E-06 $X=16470 $Y=14750 $D=0
M194 141 116 VSS VSS N12LL L=6E-08 W=7.5E-07 $X=16500 $Y=8005 $D=0
M195 574 58 99 VSS N12LL L=6E-08 W=1E-06 $X=16515 $Y=23525 $D=0
M196 97 ACTRCLKX 99 VSS N12LL L=6E-08 W=5E-07 $X=16555 $Y=25070 $D=0
M197 86 92 VSS VSS N12LL L=6E-08 W=5E-07 $X=16585 $Y=6520 $D=0
M198 VSS 96 58 VSS N12LL L=6E-08 W=5E-07 $X=16665 $Y=19040 $D=0
M199 98 97 VSS VSS N12LL L=6E-08 W=4E-07 $X=16705 $Y=29110 $D=0
M200 FCKX[7] 98 INTCLKX VSS N12LL L=6E-08 W=1.25E-06 $X=16705 $Y=33030 $D=0
M201 106 CLK 102 VSS N12LL L=6E-08 W=2.5E-06 $X=16740 $Y=14750 $D=0
M202 576 63 574 VSS N12LL L=6E-08 W=1E-06 $X=16755 $Y=23525 $D=0
M203 VSS 95 141 VSS N12LL L=6E-08 W=7.5E-07 $X=16770 $Y=8005 $D=0
M204 99 ACTRCLKX 97 VSS N12LL L=6E-08 W=5E-07 $X=16835 $Y=25070 $D=0
M205 74 58 VSS VSS N12LL L=6E-08 W=5E-07 $X=16955 $Y=19040 $D=0
M206 VSS 118 576 VSS N12LL L=6E-08 W=1E-06 $X=16995 $Y=23525 $D=0
M207 VSS 97 98 VSS N12LL L=6E-08 W=4E-07 $X=16995 $Y=29110 $D=0
M208 INTCLKX 98 FCKX[7] VSS N12LL L=6E-08 W=1.25E-06 $X=16995 $Y=33030 $D=0
M209 102 CLK 106 VSS N12LL L=6E-08 W=2.5E-06 $X=17010 $Y=14750 $D=0
M210 141 95 VSS VSS N12LL L=6E-08 W=7.5E-07 $X=17040 $Y=8005 $D=0
M211 VSS 58 74 VSS N12LL L=6E-08 W=5E-07 $X=17245 $Y=19040 $D=0
M212 WE 144 VSS VSS N12LL L=6E-08 W=5E-07 $X=17255 $Y=6540 $D=0
M213 106 CLK 102 VSS N12LL L=6E-08 W=2.5E-06 $X=17280 $Y=14750 $D=0
M214 579 118 VSS VSS N12LL L=6E-08 W=1E-06 $X=17285 $Y=23525 $D=0
M215 103 105 VSS VSS N12LL L=6E-08 W=4E-07 $X=17285 $Y=29110 $D=0
M216 FCKX[5] 103 INTCLKX VSS N12LL L=6E-08 W=1.25E-06 $X=17285 $Y=33030 $D=0
M217 VSS 116 141 VSS N12LL L=6E-08 W=7.5E-07 $X=17310 $Y=8005 $D=0
M218 105 103 VSS VSS N12LL L=6E-07 W=1.2E-07 $X=17365 $Y=30405 $D=0
M219 105 ACTRCLKX 104 VSS N12LL L=6E-08 W=5E-07 $X=17445 $Y=25070 $D=0
M220 VSS 144 WE VSS N12LL L=6E-08 W=5E-07 $X=17525 $Y=6540 $D=0
M221 581 63 579 VSS N12LL L=6E-08 W=1E-06 $X=17525 $Y=23525 $D=0
M222 102 CLK 106 VSS N12LL L=6E-08 W=2.5E-06 $X=17550 $Y=14750 $D=0
M223 VSS 105 103 VSS N12LL L=6E-08 W=4E-07 $X=17575 $Y=29110 $D=0
M224 INTCLKX 103 FCKX[5] VSS N12LL L=6E-08 W=1.25E-06 $X=17575 $Y=33030 $D=0
M225 104 ACTRCLKX 105 VSS N12LL L=6E-08 W=5E-07 $X=17725 $Y=25070 $D=0
M226 104 74 581 VSS N12LL L=6E-08 W=1E-06 $X=17765 $Y=23525 $D=0
M227 WE 144 VSS VSS N12LL L=6E-08 W=5E-07 $X=17795 $Y=6540 $D=0
M228 106 CLK 102 VSS N12LL L=6E-08 W=2.5E-06 $X=17820 $Y=14750 $D=0
M229 103 105 VSS VSS N12LL L=6E-08 W=4E-07 $X=17865 $Y=29110 $D=0
M230 FCKX[5] 103 INTCLKX VSS N12LL L=6E-08 W=1.25E-06 $X=17865 $Y=33030 $D=0
M231 107 116 VSS VSS N12LL L=2E-07 W=4E-07 $X=17960 $Y=8390 $D=0
M232 105 ACTRCLKX 104 VSS N12LL L=6E-08 W=5E-07 $X=17995 $Y=25070 $D=0
M233 VSS 144 WE VSS N12LL L=6E-08 W=5E-07 $X=18055 $Y=6540 $D=0
M234 584 VDD VSS VSS N12LL L=3E-07 W=4E-07 $X=18080 $Y=19085 $D=0
M235 VSS 105 103 VSS N12LL L=6E-08 W=4E-07 $X=18155 $Y=29110 $D=0
M236 INTCLKX 103 FCKX[5] VSS N12LL L=6E-08 W=1.25E-06 $X=18155 $Y=33030 $D=0
M237 112 107 VSS VSS N12LL L=2E-07 W=4E-07 $X=18250 $Y=7475 $D=0
M238 WE 144 VSS VSS N12LL L=6E-08 W=5E-07 $X=18325 $Y=6540 $D=0
M239 113 111 VSS VSS N12LL L=6E-08 W=4E-07 $X=18445 $Y=29110 $D=0
M240 FCKX[4] 113 INTCLKX VSS N12LL L=6E-08 W=1.25E-06 $X=18445 $Y=33030 $D=0
M241 VSS VSS 107 VSS N12LL L=2E-07 W=4E-07 $X=18450 $Y=8390 $D=0
M242 116 102 VSS VSS N12LL L=6E-08 W=2.5E-06 $X=18480 $Y=14750 $D=0
M243 VSS 144 WE VSS N12LL L=6E-08 W=5E-07 $X=18595 $Y=6540 $D=0
M244 114 A[0] 584 VSS N12LL L=6E-08 W=4E-07 $X=18600 $Y=19085 $D=0
M245 115 ACTRCLKX 111 VSS N12LL L=6E-08 W=5E-07 $X=18605 $Y=25070 $D=0
M246 VSS 113 111 VSS N12LL L=6E-07 W=1.2E-07 $X=18695 $Y=30405 $D=0
M247 VSS 111 113 VSS N12LL L=6E-08 W=4E-07 $X=18735 $Y=29110 $D=0
M248 INTCLKX 113 FCKX[4] VSS N12LL L=6E-08 W=1.25E-06 $X=18735 $Y=33030 $D=0
M249 VSS 102 116 VSS N12LL L=6E-08 W=2.5E-06 $X=18750 $Y=14750 $D=0
M250 586 74 115 VSS N12LL L=6E-08 W=1E-06 $X=18835 $Y=23525 $D=0
M251 WE 144 VSS VSS N12LL L=6E-08 W=5E-07 $X=18865 $Y=6540 $D=0
M252 111 ACTRCLKX 115 VSS N12LL L=6E-08 W=5E-07 $X=18875 $Y=25070 $D=0
M253 116 102 VSS VSS N12LL L=6E-08 W=2.5E-06 $X=19020 $Y=14750 $D=0
M254 113 111 VSS VSS N12LL L=6E-08 W=4E-07 $X=19025 $Y=29110 $D=0
M255 FCKX[4] 113 INTCLKX VSS N12LL L=6E-08 W=1.25E-06 $X=19025 $Y=33030 $D=0
M256 587 121 586 VSS N12LL L=6E-08 W=1E-06 $X=19075 $Y=23525 $D=0
M257 VSS 144 WE VSS N12LL L=6E-08 W=5E-07 $X=19135 $Y=6540 $D=0
M258 115 ACTRCLKX 111 VSS N12LL L=6E-08 W=5E-07 $X=19155 $Y=25070 $D=0
M259 136 116 VSS VSS N12LL L=6E-08 W=1.25E-06 $X=19200 $Y=7510 $D=0
M260 63 114 VSS VSS N12LL L=6E-08 W=5E-07 $X=19230 $Y=19040 $D=0
M261 VSS 102 116 VSS N12LL L=6E-08 W=2.5E-06 $X=19290 $Y=14750 $D=0
M262 VSS 118 587 VSS N12LL L=6E-08 W=1E-06 $X=19315 $Y=23525 $D=0
M263 VSS 111 113 VSS N12LL L=6E-08 W=4E-07 $X=19315 $Y=29110 $D=0
M264 INTCLKX 113 FCKX[4] VSS N12LL L=6E-08 W=1.25E-06 $X=19315 $Y=33030 $D=0
M265 WE 144 VSS VSS N12LL L=6E-08 W=5E-07 $X=19395 $Y=6540 $D=0
M266 VSS 112 136 VSS N12LL L=6E-08 W=1.25E-06 $X=19470 $Y=7510 $D=0
M267 VSS 114 63 VSS N12LL L=6E-08 W=5E-07 $X=19520 $Y=19040 $D=0
M268 INTCLKX 116 VSS VSS N12LL L=6E-08 W=2.5E-06 $X=19560 $Y=14750 $D=0
M269 590 118 VSS VSS N12LL L=6E-08 W=1E-06 $X=19605 $Y=23525 $D=0
M270 122 123 VSS VSS N12LL L=6E-08 W=4E-07 $X=19605 $Y=29110 $D=0
M271 FCKX[6] 122 INTCLKX VSS N12LL L=6E-08 W=1.25E-06 $X=19605 $Y=33030 $D=0
M272 VSS 144 WE VSS N12LL L=6E-08 W=5E-07 $X=19665 $Y=6540 $D=0
M273 123 122 VSS VSS N12LL L=6E-07 W=1.2E-07 $X=19685 $Y=30405 $D=0
M274 136 112 VSS VSS N12LL L=6E-08 W=1.25E-06 $X=19740 $Y=7510 $D=0
M275 123 ACTRCLKX 124 VSS N12LL L=6E-08 W=5E-07 $X=19765 $Y=25070 $D=0
M276 121 63 VSS VSS N12LL L=6E-08 W=5E-07 $X=19810 $Y=19040 $D=0
M277 VSS 116 INTCLKX VSS N12LL L=6E-08 W=2.5E-06 $X=19830 $Y=14750 $D=0
M278 591 121 590 VSS N12LL L=6E-08 W=1E-06 $X=19845 $Y=23525 $D=0
M279 VSS 123 122 VSS N12LL L=6E-08 W=4E-07 $X=19895 $Y=29110 $D=0
M280 INTCLKX 122 FCKX[6] VSS N12LL L=6E-08 W=1.25E-06 $X=19895 $Y=33030 $D=0
M281 VSS 116 136 VSS N12LL L=6E-08 W=1.25E-06 $X=20010 $Y=7510 $D=0
M282 124 ACTRCLKX 123 VSS N12LL L=6E-08 W=5E-07 $X=20045 $Y=25070 $D=0
M283 124 58 591 VSS N12LL L=6E-08 W=1E-06 $X=20085 $Y=23525 $D=0
M284 INTCLKX 116 VSS VSS N12LL L=6E-08 W=2.5E-06 $X=20100 $Y=14750 $D=0
M285 VSS 63 121 VSS N12LL L=6E-08 W=5E-07 $X=20100 $Y=19040 $D=0
M286 122 123 VSS VSS N12LL L=6E-08 W=4E-07 $X=20185 $Y=29110 $D=0
M287 FCKX[6] 122 INTCLKX VSS N12LL L=6E-08 W=1.25E-06 $X=20185 $Y=33030 $D=0
M288 126 WEN VSS VSS N12LL L=6E-08 W=4E-07 $X=20315 $Y=6565 $D=0
M289 123 ACTRCLKX 124 VSS N12LL L=6E-08 W=5E-07 $X=20315 $Y=25070 $D=0
M290 VSS 116 INTCLKX VSS N12LL L=6E-08 W=2.5E-06 $X=20370 $Y=14750 $D=0
M291 VSS 123 122 VSS N12LL L=6E-08 W=4E-07 $X=20475 $Y=29110 $D=0
M292 INTCLKX 122 FCKX[6] VSS N12LL L=6E-08 W=1.25E-06 $X=20475 $Y=33030 $D=0
M293 129 136 VSS VSS N12LL L=6E-08 W=1E-06 $X=20610 $Y=7760 $D=0
M294 INTCLKX 116 VSS VSS N12LL L=6E-08 W=2.5E-06 $X=20640 $Y=14750 $D=0
M295 VSS 136 129 VSS N12LL L=6E-08 W=1E-06 $X=20880 $Y=7760 $D=0
M296 VSS 116 INTCLKX VSS N12LL L=6E-08 W=2.5E-06 $X=20910 $Y=14750 $D=0
M297 VSS 126 130 VSS N12LL L=3E-07 W=4E-07 $X=20990 $Y=6565 $D=0
M298 129 136 VSS VSS N12LL L=6E-08 W=1E-06 $X=21150 $Y=7760 $D=0
M299 INTCLKX 116 VSS VSS N12LL L=6E-08 W=2.5E-06 $X=21180 $Y=14750 $D=0
M300 VSS 116 INTCLKX VSS N12LL L=6E-08 W=2.5E-06 $X=21450 $Y=14750 $D=0
M301 133 130 VSS VSS N12LL L=2E-07 W=4E-07 $X=21580 $Y=6565 $D=0
M302 DCTRCLKX 129 VSS VSS N12LL L=6E-08 W=2.5E-06 $X=22110 $Y=14750 $D=0
M303 VSS 129 DCTRCLKX VSS N12LL L=6E-08 W=2.5E-06 $X=22380 $Y=14750 $D=0
M304 134 133 VSS VSS N12LL L=6E-08 W=1E-06 $X=22390 $Y=6585 $D=0
M305 DCTRCLK 136 VSS VSS N12LL L=6E-08 W=2.5E-06 $X=22650 $Y=14750 $D=0
M306 138 ACTRCLKX 134 VSS N12LL L=6E-08 W=1E-06 $X=22660 $Y=6585 $D=0
M307 VSS 136 DCTRCLK VSS N12LL L=6E-08 W=2.5E-06 $X=22920 $Y=14750 $D=0
M308 ACTRCLK 136 VSS VSS N12LL L=6E-08 W=2.5E-06 $X=23190 $Y=14750 $D=0
M309 VSS 140 138 VSS N12LL L=6E-07 W=1.2E-07 $X=23355 $Y=6840 $D=0
M310 VSS 136 ACTRCLK VSS N12LL L=6E-08 W=2.5E-06 $X=23460 $Y=14750 $D=0
M311 ACTRCLKX ACTRCLK VSS VSS N12LL L=6E-08 W=2.5E-06 $X=23730 $Y=14750 $D=0
M312 VSS ACTRCLK ACTRCLKX VSS N12LL L=6E-08 W=2.5E-06 $X=24000 $Y=14750 $D=0
M313 VSS 138 140 VSS N12LL L=6E-08 W=1E-06 $X=24020 $Y=6560 $D=0
M314 SACK1 116 VSS VSS N12LL L=6E-08 W=2.5E-06 $X=24270 $Y=14750 $D=0
M315 143 116 VSS VSS N12LL L=6E-08 W=1.5E-06 $X=24290 $Y=6560 $D=0
M316 VSS 116 SACK1 VSS N12LL L=6E-08 W=2.5E-06 $X=24540 $Y=14750 $D=0
M317 144 140 143 VSS N12LL L=6E-08 W=1.5E-06 $X=24560 $Y=6560 $D=0
M318 SACK4 141 VSS VSS N12LL L=6E-08 W=2.5E-06 $X=24810 $Y=14750 $D=0
M319 143 140 144 VSS N12LL L=6E-08 W=1.5E-06 $X=24830 $Y=6560 $D=0
M320 VSS 141 SACK4 VSS N12LL L=6E-08 W=2.5E-06 $X=25080 $Y=14750 $D=0
M321 VSS 116 143 VSS N12LL L=6E-08 W=1.5E-06 $X=25110 $Y=6560 $D=0
M322 4 12 INTCLKX VDD P12LL L=6E-08 W=5E-07 $X=5365 $Y=24635 $D=1
M323 RWL 4 VDD VDD P12LL L=6E-08 W=2.5E-06 $X=5365 $Y=30345 $D=1
M324 VDD 11 6 VDD P12LL L=6E-08 W=8E-07 $X=5565 $Y=13735 $D=1
M325 6 ACTRCLK 13 VDD P12LL L=6E-08 W=5E-07 $X=5565 $Y=17440 $D=1
M326 VDD 13 12 VDD P12LL L=6E-08 W=8E-07 $X=5565 $Y=19260 $D=1
M327 INTCLKX 12 4 VDD P12LL L=6E-08 W=5E-07 $X=5655 $Y=24635 $D=1
M328 VDD 7 4 VDD P12LL L=6E-08 W=1E-06 $X=5655 $Y=25875 $D=1
M329 VDD 4 RWL VDD P12LL L=6E-08 W=2.5E-06 $X=5655 $Y=30345 $D=1
M330 13 ACTRCLK 6 VDD P12LL L=6E-08 W=5E-07 $X=5835 $Y=17440 $D=1
M331 VDD S[0] 8 VDD P12LL L=6E-08 W=4E-07 $X=5850 $Y=5075 $D=1
M332 VDD S[1] 9 VDD P12LL L=6E-08 W=4E-07 $X=5850 $Y=8185 $D=1
M333 13 12 VDD VDD P12LL L=3E-07 W=1.2E-07 $X=5895 $Y=19940 $D=1
M334 4 12 INTCLKX VDD P12LL L=6E-08 W=5E-07 $X=5925 $Y=24635 $D=1
M335 4 7 VDD VDD P12LL L=6E-08 W=1E-06 $X=5925 $Y=25875 $D=1
M336 RWL 4 VDD VDD P12LL L=6E-08 W=2.5E-06 $X=5945 $Y=30345 $D=1
M337 617 VSS VDD VDD P12LL L=1E-07 W=4E-07 $X=5960 $Y=12400 $D=1
M338 7 12 VDD VDD P12LL L=6E-08 W=8E-07 $X=6035 $Y=23075 $D=1
M339 23 8 VDD VDD P12LL L=6E-08 W=4E-07 $X=6120 $Y=5075 $D=1
M340 16 9 VDD VDD P12LL L=6E-08 W=4E-07 $X=6120 $Y=8185 $D=1
M341 VDD 19 11 VDD P12LL L=6E-08 W=8E-07 $X=6155 $Y=13735 $D=1
M342 INTCLKX 12 4 VDD P12LL L=6E-08 W=5E-07 $X=6215 $Y=24635 $D=1
M343 17 RDE 617 VDD P12LL L=6E-08 W=4E-07 $X=6230 $Y=12400 $D=1
M344 VDD 4 RWL VDD P12LL L=6E-08 W=2.5E-06 $X=6235 $Y=30345 $D=1
M345 19 17 VDD VDD P12LL L=6E-08 W=8E-07 $X=6425 $Y=13735 $D=1
M346 21 9 VDD VDD P12LL L=6E-08 W=4E-07 $X=6720 $Y=5075 $D=1
M347 22 9 VDD VDD P12LL L=6E-08 W=4E-07 $X=6720 $Y=8185 $D=1
M348 VDD 8 21 VDD P12LL L=6E-08 W=4E-07 $X=6990 $Y=5075 $D=1
M349 VDD 23 22 VDD P12LL L=6E-08 W=4E-07 $X=6990 $Y=8185 $D=1
M350 24 8 VDD VDD P12LL L=6E-08 W=4E-07 $X=7260 $Y=5075 $D=1
M351 25 23 VDD VDD P12LL L=6E-08 W=4E-07 $X=7260 $Y=8185 $D=1
M352 VDD 16 24 VDD P12LL L=6E-08 W=4E-07 $X=7530 $Y=5075 $D=1
M353 VDD 16 25 VDD P12LL L=6E-08 W=4E-07 $X=7530 $Y=8185 $D=1
M354 621 30 46 VDD P12LL L=6E-08 W=7E-07 $X=7565 $Y=14015 $D=1
M355 VDD RDE 621 VDD P12LL L=6E-08 W=7E-07 $X=7795 $Y=14015 $D=1
M356 PXA[3] 29 VDD VDD P12LL L=6E-08 W=3.5E-06 $X=7810 $Y=30770 $D=1
M357 27 46 VDD VDD P12LL L=6E-08 W=1.5E-06 $X=7830 $Y=19095 $D=1
M358 VDD A[3] 30 VDD P12LL L=6E-08 W=4E-07 $X=7950 $Y=12400 $D=1
M359 29 ACTRCLK 27 VDD P12LL L=6E-08 W=2.5E-06 $X=7955 $Y=24130 $D=1
M360 40 45 VDD VDD P12LL L=6E-08 W=1E-06 $X=8010 $Y=2955 $D=1
M361 36 PXA[2] VDD VDD P12LL L=3E-07 W=1.2E-07 $X=8090 $Y=34920 $D=1
M362 VDD 29 PXA[3] VDD P12LL L=6E-08 W=3.5E-06 $X=8100 $Y=30770 $D=1
M363 VDD 42 27 VDD P12LL L=6E-08 W=1.5E-06 $X=8110 $Y=19095 $D=1
M364 622 RDE VDD VDD P12LL L=6E-08 W=1.4E-06 $X=8145 $Y=13315 $D=1
M365 VDD 25 37 VDD P12LL L=6E-08 W=4E-07 $X=8220 $Y=4860 $D=1
M366 31 30 VDD VDD P12LL L=6E-08 W=4E-07 $X=8280 $Y=12400 $D=1
M367 VDD PXA[3] 29 VDD P12LL L=3E-07 W=1.2E-07 $X=8345 $Y=35525 $D=1
M368 34 42 VDD VDD P12LL L=6E-08 W=1.5E-06 $X=8380 $Y=19095 $D=1
M369 PXA[2] 36 VDD VDD P12LL L=6E-08 W=3.5E-06 $X=8390 $Y=30770 $D=1
M370 32 31 622 VDD P12LL L=6E-08 W=1.4E-06 $X=8435 $Y=13315 $D=1
M371 34 ACTRCLK 36 VDD P12LL L=6E-08 W=2.5E-06 $X=8535 $Y=24130 $D=1
M372 EMCLK 25 40 VDD P12LL L=6E-08 W=1E-06 $X=8630 $Y=5420 $D=1
M373 VDD 32 34 VDD P12LL L=6E-08 W=1.5E-06 $X=8660 $Y=19095 $D=1
M374 VDD 36 PXA[2] VDD P12LL L=6E-08 W=3.5E-06 $X=8680 $Y=30770 $D=1
M375 40 25 EMCLK VDD P12LL L=6E-08 W=1.5E-06 $X=8900 $Y=4920 $D=1
M376 PXA[0] 38 VDD VDD P12LL L=6E-08 W=3.5E-06 $X=9020 $Y=30770 $D=1
M377 41 32 VDD VDD P12LL L=6E-08 W=1.5E-06 $X=9040 $Y=19095 $D=1
M378 48 PXA[1] VDD VDD P12LL L=3E-07 W=1.2E-07 $X=9115 $Y=35525 $D=1
M379 38 ACTRCLK 41 VDD P12LL L=6E-08 W=2.5E-06 $X=9165 $Y=24130 $D=1
M380 VDD 45 40 VDD P12LL L=6E-08 W=1.5E-06 $X=9215 $Y=4920 $D=1
M381 VDD 49 42 VDD P12LL L=6E-08 W=1.4E-06 $X=9265 $Y=13315 $D=1
M382 VDD 38 PXA[0] VDD P12LL L=6E-08 W=3.5E-06 $X=9310 $Y=30770 $D=1
M383 VDD 47 41 VDD P12LL L=6E-08 W=1.5E-06 $X=9320 $Y=19095 $D=1
M384 VDD PXA[0] 38 VDD P12LL L=3E-07 W=1.2E-07 $X=9370 $Y=34920 $D=1
M385 623 VSS VDD VDD P12LL L=1E-07 W=4E-07 $X=9405 $Y=12400 $D=1
M386 45 102 VDD VDD P12LL L=6E-08 W=1.5E-06 $X=9515 $Y=4920 $D=1
M387 47 42 VDD VDD P12LL L=6E-08 W=1.4E-06 $X=9555 $Y=13315 $D=1
M388 50 47 VDD VDD P12LL L=6E-08 W=1.5E-06 $X=9590 $Y=19095 $D=1
M389 PXA[1] 48 VDD VDD P12LL L=6E-08 W=3.5E-06 $X=9600 $Y=30770 $D=1
M390 50 ACTRCLK 48 VDD P12LL L=6E-08 W=2.5E-06 $X=9745 $Y=24130 $D=1
M391 49 A[4] 623 VDD P12LL L=6E-08 W=4E-07 $X=9770 $Y=12400 $D=1
M392 VDD 46 50 VDD P12LL L=6E-08 W=1.5E-06 $X=9870 $Y=19095 $D=1
M393 VDD 48 PXA[1] VDD P12LL L=6E-08 W=3.5E-06 $X=9890 $Y=30770 $D=1
M394 VDD FB 52 VDD P12LL L=6E-08 W=8E-07 $X=10135 $Y=5645 $D=1
M395 80 52 VDD VDD P12LL L=6E-08 W=1.25E-06 $X=10495 $Y=5195 $D=1
M396 VDD 52 80 VDD P12LL L=6E-08 W=1.25E-06 $X=10765 $Y=5195 $D=1
M397 VDD 24 53 VDD P12LL L=6E-08 W=4E-07 $X=10890 $Y=13475 $D=1
M398 VDD 40 55 VDD P12LL L=1.5E-07 W=7E-07 $X=10945 $Y=10650 $D=1
M399 VDD 55 54 VDD P12LL L=6E-08 W=6.25E-07 $X=11085 $Y=12110 $D=1
M400 62 22 VDD VDD P12LL L=6E-08 W=4E-07 $X=11160 $Y=13475 $D=1
M401 54 55 VDD VDD P12LL L=6E-08 W=1.25E-06 $X=11385 $Y=10650 $D=1
M402 54 55 VDD VDD P12LL L=6E-08 W=6.25E-07 $X=11385 $Y=12110 $D=1
M403 FB 45 VDD VDD P12LL L=6E-08 W=1.2E-06 $X=11410 $Y=4770 $D=1
M404 59 57 VDD VDD P12LL L=6E-08 W=4E-07 $X=11485 $Y=28025 $D=1
M405 FCKX[3] 57 INTCLKX VDD P12LL L=6E-08 W=1.25E-06 $X=11485 $Y=31220 $D=1
M406 FCKX[3] 59 VDD VDD P12LL L=6E-08 W=1.25E-06 $X=11485 $Y=34780 $D=1
M407 60 ACTRCLK 57 VDD P12LL L=6E-08 W=5E-07 $X=11645 $Y=26070 $D=1
M408 VDD 45 FB VDD P12LL L=6E-08 W=1.2E-06 $X=11680 $Y=4770 $D=1
M409 EMCLK 24 54 VDD P12LL L=6E-08 W=1.25E-06 $X=11715 $Y=10650 $D=1
M410 67 21 VDD VDD P12LL L=6E-08 W=4E-07 $X=11760 $Y=13475 $D=1
M411 VDD 58 60 VDD P12LL L=6E-08 W=1E-06 $X=11775 $Y=21925 $D=1
M412 VDD 57 59 VDD P12LL L=6E-08 W=4E-07 $X=11775 $Y=28025 $D=1
M413 INTCLKX 57 FCKX[3] VDD P12LL L=6E-08 W=1.25E-06 $X=11775 $Y=31220 $D=1
M414 VDD 59 FCKX[3] VDD P12LL L=6E-08 W=1.25E-06 $X=11775 $Y=34780 $D=1
M415 57 ACTRCLK 60 VDD P12LL L=6E-08 W=5E-07 $X=11915 $Y=26070 $D=1
M416 54 24 EMCLK VDD P12LL L=6E-08 W=1.25E-06 $X=11985 $Y=10650 $D=1
M417 VDD 59 57 VDD P12LL L=3E-07 W=1.2E-07 $X=12025 $Y=27185 $D=1
M418 60 63 VDD VDD P12LL L=6E-08 W=1E-06 $X=12065 $Y=21925 $D=1
M419 59 57 VDD VDD P12LL L=6E-08 W=4E-07 $X=12065 $Y=28025 $D=1
M420 FCKX[3] 57 INTCLKX VDD P12LL L=6E-08 W=1.25E-06 $X=12065 $Y=31220 $D=1
M421 FCKX[3] 59 VDD VDD P12LL L=6E-08 W=1.25E-06 $X=12065 $Y=34780 $D=1
M422 60 ACTRCLK 57 VDD P12LL L=6E-08 W=5E-07 $X=12195 $Y=26070 $D=1
M423 84 118 VDD VDD P12LL L=6E-08 W=1E-06 $X=12265 $Y=20095 $D=1
M424 VDD CLK 64 VDD P12LL L=6E-08 W=4E-07 $X=12330 $Y=5455 $D=1
M425 VDD 84 60 VDD P12LL L=6E-08 W=1E-06 $X=12355 $Y=21925 $D=1
M426 VDD 57 59 VDD P12LL L=6E-08 W=4E-07 $X=12355 $Y=28025 $D=1
M427 INTCLKX 57 FCKX[3] VDD P12LL L=6E-08 W=1.25E-06 $X=12355 $Y=31220 $D=1
M428 VDD 59 FCKX[3] VDD P12LL L=6E-08 W=1.25E-06 $X=12355 $Y=34780 $D=1
M429 VDD 118 84 VDD P12LL L=6E-08 W=1E-06 $X=12555 $Y=20095 $D=1
M430 EMCLK 22 66 VDD P12LL L=6E-08 W=1.25E-06 $X=12595 $Y=10650 $D=1
M431 69 84 VDD VDD P12LL L=6E-08 W=1E-06 $X=12645 $Y=21925 $D=1
M432 68 70 VDD VDD P12LL L=6E-08 W=4E-07 $X=12645 $Y=28025 $D=1
M433 FCKX[1] 70 INTCLKX VDD P12LL L=6E-08 W=1.25E-06 $X=12645 $Y=31220 $D=1
M434 FCKX[1] 68 VDD VDD P12LL L=6E-08 W=1.25E-06 $X=12645 $Y=34780 $D=1
M435 626 CLK VDD VDD P12LL L=6E-08 W=1E-06 $X=12670 $Y=4855 $D=1
M436 70 68 VDD VDD P12LL L=3E-07 W=1.2E-07 $X=12735 $Y=27185 $D=1
M437 VDD 66 65 VDD P12LL L=1.5E-07 W=7E-07 $X=12740 $Y=13120 $D=1
M438 70 ACTRCLK 69 VDD P12LL L=6E-08 W=5E-07 $X=12805 $Y=26070 $D=1
M439 118 75 VDD VDD P12LL L=6E-08 W=1E-06 $X=12845 $Y=20095 $D=1
M440 66 22 EMCLK VDD P12LL L=6E-08 W=1.25E-06 $X=12865 $Y=10650 $D=1
M441 78 CEN 626 VDD P12LL L=6E-08 W=1E-06 $X=12910 $Y=4855 $D=1
M442 VDD 63 69 VDD P12LL L=6E-08 W=1E-06 $X=12935 $Y=21925 $D=1
M443 VDD 70 68 VDD P12LL L=6E-08 W=4E-07 $X=12935 $Y=28025 $D=1
M444 INTCLKX 70 FCKX[1] VDD P12LL L=6E-08 W=1.25E-06 $X=12935 $Y=31220 $D=1
M445 VDD 68 FCKX[1] VDD P12LL L=6E-08 W=1.25E-06 $X=12935 $Y=34780 $D=1
M446 69 ACTRCLK 70 VDD P12LL L=6E-08 W=5E-07 $X=13085 $Y=26070 $D=1
M447 VDD 75 118 VDD P12LL L=6E-08 W=1E-06 $X=13135 $Y=20095 $D=1
M448 VDD 79 66 VDD P12LL L=6E-08 W=1.25E-06 $X=13155 $Y=10650 $D=1
M449 69 74 VDD VDD P12LL L=6E-08 W=1E-06 $X=13225 $Y=21925 $D=1
M450 68 70 VDD VDD P12LL L=6E-08 W=4E-07 $X=13225 $Y=28025 $D=1
M451 FCKX[1] 70 INTCLKX VDD P12LL L=6E-08 W=1.25E-06 $X=13225 $Y=31220 $D=1
M452 FCKX[1] 68 VDD VDD P12LL L=6E-08 W=1.25E-06 $X=13225 $Y=34780 $D=1
M453 VDD 85 78 VDD P12LL L=3E-07 W=1.2E-07 $X=13270 $Y=5735 $D=1
M454 70 ACTRCLK 69 VDD P12LL L=6E-08 W=5E-07 $X=13355 $Y=26070 $D=1
M455 VDD 65 77 VDD P12LL L=6E-08 W=1.25E-06 $X=13420 $Y=12570 $D=1
M456 66 79 VDD VDD P12LL L=6E-08 W=1.25E-06 $X=13425 $Y=10650 $D=1
M457 VDD 70 68 VDD P12LL L=6E-08 W=4E-07 $X=13515 $Y=28025 $D=1
M458 INTCLKX 70 FCKX[1] VDD P12LL L=6E-08 W=1.25E-06 $X=13515 $Y=31220 $D=1
M459 VDD 68 FCKX[1] VDD P12LL L=6E-08 W=1.25E-06 $X=13515 $Y=34780 $D=1
M460 77 65 VDD VDD P12LL L=6E-08 W=1.25E-06 $X=13750 $Y=12570 $D=1
M461 629 A[2] 75 VDD P12LL L=6E-08 W=4E-07 $X=13765 $Y=20425 $D=1
M462 81 76 VDD VDD P12LL L=6E-08 W=4E-07 $X=13805 $Y=28025 $D=1
M463 FCKX[0] 76 INTCLKX VDD P12LL L=6E-08 W=1.25E-06 $X=13805 $Y=31220 $D=1
M464 FCKX[0] 81 VDD VDD P12LL L=6E-08 W=1.25E-06 $X=13805 $Y=34780 $D=1
M465 82 ACTRCLK 76 VDD P12LL L=6E-08 W=5E-07 $X=13965 $Y=26070 $D=1
M466 EMCLK 21 77 VDD P12LL L=6E-08 W=1.25E-06 $X=14020 $Y=12570 $D=1
M467 79 54 VDD VDD P12LL L=1.5E-07 W=7E-07 $X=14035 $Y=10650 $D=1
M468 VDD 74 82 VDD P12LL L=6E-08 W=1E-06 $X=14095 $Y=21925 $D=1
M469 VDD 76 81 VDD P12LL L=6E-08 W=4E-07 $X=14095 $Y=28025 $D=1
M470 INTCLKX 76 FCKX[0] VDD P12LL L=6E-08 W=1.25E-06 $X=14095 $Y=31220 $D=1
M471 VDD 81 FCKX[0] VDD P12LL L=6E-08 W=1.25E-06 $X=14095 $Y=34780 $D=1
M472 85 78 VDD VDD P12LL L=6E-08 W=8E-07 $X=14200 $Y=5055 $D=1
M473 76 ACTRCLK 82 VDD P12LL L=6E-08 W=5E-07 $X=14235 $Y=26070 $D=1
M474 VDD VSS 629 VDD P12LL L=1E-07 W=4E-07 $X=14245 $Y=20425 $D=1
M475 77 21 EMCLK VDD P12LL L=6E-08 W=1.25E-06 $X=14310 $Y=12570 $D=1
M476 VDD 81 76 VDD P12LL L=3E-07 W=1.2E-07 $X=14345 $Y=27185 $D=1
M477 82 121 VDD VDD P12LL L=6E-08 W=1E-06 $X=14385 $Y=21925 $D=1
M478 81 76 VDD VDD P12LL L=6E-08 W=4E-07 $X=14385 $Y=28025 $D=1
M479 FCKX[0] 76 INTCLKX VDD P12LL L=6E-08 W=1.25E-06 $X=14385 $Y=31220 $D=1
M480 FCKX[0] 81 VDD VDD P12LL L=6E-08 W=1.25E-06 $X=14385 $Y=34780 $D=1
M481 82 ACTRCLK 76 VDD P12LL L=6E-08 W=5E-07 $X=14515 $Y=26070 $D=1
M482 VDD 84 82 VDD P12LL L=6E-08 W=1E-06 $X=14675 $Y=21925 $D=1
M483 VDD 76 81 VDD P12LL L=6E-08 W=4E-07 $X=14675 $Y=28025 $D=1
M484 INTCLKX 76 FCKX[0] VDD P12LL L=6E-08 W=1.25E-06 $X=14675 $Y=31220 $D=1
M485 VDD 81 FCKX[0] VDD P12LL L=6E-08 W=1.25E-06 $X=14675 $Y=34780 $D=1
M486 631 85 87 VDD P12LL L=6E-08 W=1E-06 $X=14895 $Y=4920 $D=1
M487 102 80 VDD VDD P12LL L=6E-08 W=1.25E-06 $X=14900 $Y=12600 $D=1
M488 VDD 116 89 VDD P12LL L=3E-07 W=3E-07 $X=14910 $Y=10010 $D=1
M489 93 84 VDD VDD P12LL L=6E-08 W=1E-06 $X=14965 $Y=21925 $D=1
M490 90 91 VDD VDD P12LL L=6E-08 W=4E-07 $X=14965 $Y=28025 $D=1
M491 FCKX[2] 91 INTCLKX VDD P12LL L=6E-08 W=1.25E-06 $X=14965 $Y=31220 $D=1
M492 FCKX[2] 90 VDD VDD P12LL L=6E-08 W=1.25E-06 $X=14965 $Y=34780 $D=1
M493 VDD 116 102 VDD P12LL L=2E-07 W=1.2E-07 $X=15000 $Y=11125 $D=1
M494 91 90 VDD VDD P12LL L=3E-07 W=1.2E-07 $X=15055 $Y=27185 $D=1
M495 91 ACTRCLK 93 VDD P12LL L=6E-08 W=5E-07 $X=15125 $Y=26070 $D=1
M496 VDD CLK 631 VDD P12LL L=6E-08 W=1E-06 $X=15165 $Y=4920 $D=1
M497 VDD 80 102 VDD P12LL L=6E-08 W=1.25E-06 $X=15170 $Y=12600 $D=1
M498 633 VSS VDD VDD P12LL L=1E-07 W=4E-07 $X=15225 $Y=20425 $D=1
M499 VDD 121 93 VDD P12LL L=6E-08 W=1E-06 $X=15255 $Y=21925 $D=1
M500 VDD 91 90 VDD P12LL L=6E-08 W=4E-07 $X=15255 $Y=28025 $D=1
M501 INTCLKX 91 FCKX[2] VDD P12LL L=6E-08 W=1.25E-06 $X=15255 $Y=31220 $D=1
M502 VDD 90 FCKX[2] VDD P12LL L=6E-08 W=1.25E-06 $X=15255 $Y=34780 $D=1
M503 95 89 VDD VDD P12LL L=2E-07 W=4E-07 $X=15400 $Y=10010 $D=1
M504 93 ACTRCLK 91 VDD P12LL L=6E-08 W=5E-07 $X=15405 $Y=26070 $D=1
M505 92 87 VDD VDD P12LL L=6E-08 W=1E-06 $X=15435 $Y=4920 $D=1
M506 102 80 VDD VDD P12LL L=6E-08 W=1.25E-06 $X=15440 $Y=12600 $D=1
M507 93 58 VDD VDD P12LL L=6E-08 W=1E-06 $X=15545 $Y=21925 $D=1
M508 90 91 VDD VDD P12LL L=6E-08 W=4E-07 $X=15545 $Y=28025 $D=1
M509 FCKX[2] 91 INTCLKX VDD P12LL L=6E-08 W=1.25E-06 $X=15545 $Y=31220 $D=1
M510 FCKX[2] 90 VDD VDD P12LL L=6E-08 W=1.25E-06 $X=15545 $Y=34780 $D=1
M511 91 ACTRCLK 93 VDD P12LL L=6E-08 W=5E-07 $X=15675 $Y=26070 $D=1
M512 VDD 80 102 VDD P12LL L=6E-08 W=1.25E-06 $X=15710 $Y=12600 $D=1
M513 96 A[1] 633 VDD P12LL L=6E-08 W=4E-07 $X=15745 $Y=20425 $D=1
M514 VDD 91 90 VDD P12LL L=6E-08 W=4E-07 $X=15835 $Y=28025 $D=1
M515 INTCLKX 91 FCKX[2] VDD P12LL L=6E-08 W=1.25E-06 $X=15835 $Y=31220 $D=1
M516 VDD 90 FCKX[2] VDD P12LL L=6E-08 W=1.25E-06 $X=15835 $Y=34780 $D=1
M517 102 80 VDD VDD P12LL L=6E-08 W=1.25E-06 $X=15980 $Y=12600 $D=1
M518 86 92 VDD VDD P12LL L=6E-08 W=1E-06 $X=16045 $Y=4920 $D=1
M519 98 97 VDD VDD P12LL L=6E-08 W=4E-07 $X=16125 $Y=28025 $D=1
M520 FCKX[7] 97 INTCLKX VDD P12LL L=6E-08 W=1.25E-06 $X=16125 $Y=31220 $D=1
M521 FCKX[7] 98 VDD VDD P12LL L=6E-08 W=1.25E-06 $X=16125 $Y=34780 $D=1
M522 VDD 80 102 VDD P12LL L=6E-08 W=1.25E-06 $X=16250 $Y=12600 $D=1
M523 99 ACTRCLK 97 VDD P12LL L=6E-08 W=5E-07 $X=16285 $Y=26070 $D=1
M524 VDD 92 86 VDD P12LL L=6E-08 W=1E-06 $X=16315 $Y=4920 $D=1
M525 58 96 VDD VDD P12LL L=6E-08 W=1E-06 $X=16375 $Y=20095 $D=1
M526 VDD 58 99 VDD P12LL L=6E-08 W=1E-06 $X=16415 $Y=21925 $D=1
M527 VDD 97 98 VDD P12LL L=6E-08 W=4E-07 $X=16415 $Y=28025 $D=1
M528 INTCLKX 97 FCKX[7] VDD P12LL L=6E-08 W=1.25E-06 $X=16415 $Y=31220 $D=1
M529 VDD 98 FCKX[7] VDD P12LL L=6E-08 W=1.25E-06 $X=16415 $Y=34780 $D=1
M530 101 116 141 VDD P12LL L=6E-08 W=1E-06 $X=16500 $Y=9395 $D=1
M531 102 80 VDD VDD P12LL L=6E-08 W=1.25E-06 $X=16520 $Y=12600 $D=1
M532 97 ACTRCLK 99 VDD P12LL L=6E-08 W=5E-07 $X=16555 $Y=26070 $D=1
M533 86 92 VDD VDD P12LL L=6E-08 W=1E-06 $X=16585 $Y=4920 $D=1
M534 VDD 96 58 VDD P12LL L=6E-08 W=1E-06 $X=16665 $Y=20095 $D=1
M535 VDD 98 97 VDD P12LL L=3E-07 W=1.2E-07 $X=16665 $Y=27185 $D=1
M536 99 63 VDD VDD P12LL L=6E-08 W=1E-06 $X=16705 $Y=21925 $D=1
M537 98 97 VDD VDD P12LL L=6E-08 W=4E-07 $X=16705 $Y=28025 $D=1
M538 FCKX[7] 97 INTCLKX VDD P12LL L=6E-08 W=1.25E-06 $X=16705 $Y=31220 $D=1
M539 FCKX[7] 98 VDD VDD P12LL L=6E-08 W=1.25E-06 $X=16705 $Y=34780 $D=1
M540 VDD 95 101 VDD P12LL L=6E-08 W=1E-06 $X=16770 $Y=9395 $D=1
M541 VDD 80 102 VDD P12LL L=6E-08 W=1.25E-06 $X=16790 $Y=12600 $D=1
M542 99 ACTRCLK 97 VDD P12LL L=6E-08 W=5E-07 $X=16835 $Y=26070 $D=1
M543 74 58 VDD VDD P12LL L=6E-08 W=1E-06 $X=16955 $Y=20095 $D=1
M544 VDD 118 99 VDD P12LL L=6E-08 W=1E-06 $X=16995 $Y=21925 $D=1
M545 VDD 97 98 VDD P12LL L=6E-08 W=4E-07 $X=16995 $Y=28025 $D=1
M546 INTCLKX 97 FCKX[7] VDD P12LL L=6E-08 W=1.25E-06 $X=16995 $Y=31220 $D=1
M547 VDD 98 FCKX[7] VDD P12LL L=6E-08 W=1.25E-06 $X=16995 $Y=34780 $D=1
M548 101 95 VDD VDD P12LL L=6E-08 W=1E-06 $X=17040 $Y=9395 $D=1
M549 VDD 58 74 VDD P12LL L=6E-08 W=1E-06 $X=17245 $Y=20095 $D=1
M550 WE 144 VDD VDD P12LL L=6E-08 W=1E-06 $X=17255 $Y=4905 $D=1
M551 104 118 VDD VDD P12LL L=6E-08 W=1E-06 $X=17285 $Y=21925 $D=1
M552 103 105 VDD VDD P12LL L=6E-08 W=4E-07 $X=17285 $Y=28025 $D=1
M553 FCKX[5] 105 INTCLKX VDD P12LL L=6E-08 W=1.25E-06 $X=17285 $Y=31220 $D=1
M554 FCKX[5] 103 VDD VDD P12LL L=6E-08 W=1.25E-06 $X=17285 $Y=34780 $D=1
M555 141 116 101 VDD P12LL L=6E-08 W=1E-06 $X=17310 $Y=9395 $D=1
M556 105 103 VDD VDD P12LL L=3E-07 W=1.2E-07 $X=17375 $Y=27185 $D=1
M557 116 102 VDD VDD P12LL L=6E-08 W=2.5E-06 $X=17400 $Y=11350 $D=1
M558 105 ACTRCLK 104 VDD P12LL L=6E-08 W=5E-07 $X=17445 $Y=26070 $D=1
M559 VDD 144 WE VDD P12LL L=6E-08 W=1E-06 $X=17525 $Y=4905 $D=1
M560 VDD 63 104 VDD P12LL L=6E-08 W=1E-06 $X=17575 $Y=21925 $D=1
M561 VDD 105 103 VDD P12LL L=6E-08 W=4E-07 $X=17575 $Y=28025 $D=1
M562 INTCLKX 105 FCKX[5] VDD P12LL L=6E-08 W=1.25E-06 $X=17575 $Y=31220 $D=1
M563 VDD 103 FCKX[5] VDD P12LL L=6E-08 W=1.25E-06 $X=17575 $Y=34780 $D=1
M564 VDD 102 116 VDD P12LL L=6E-08 W=2.5E-06 $X=17670 $Y=11350 $D=1
M565 104 ACTRCLK 105 VDD P12LL L=6E-08 W=5E-07 $X=17725 $Y=26070 $D=1
M566 WE 144 VDD VDD P12LL L=6E-08 W=1E-06 $X=17795 $Y=4905 $D=1
M567 104 74 VDD VDD P12LL L=6E-08 W=1E-06 $X=17865 $Y=21925 $D=1
M568 103 105 VDD VDD P12LL L=6E-08 W=4E-07 $X=17865 $Y=28025 $D=1
M569 FCKX[5] 105 INTCLKX VDD P12LL L=6E-08 W=1.25E-06 $X=17865 $Y=31220 $D=1
M570 FCKX[5] 103 VDD VDD P12LL L=6E-08 W=1.25E-06 $X=17865 $Y=34780 $D=1
M571 116 102 VDD VDD P12LL L=6E-08 W=2.5E-06 $X=17940 $Y=11350 $D=1
M572 638 116 107 VDD P12LL L=2E-07 W=8E-07 $X=17960 $Y=9190 $D=1
M573 105 ACTRCLK 104 VDD P12LL L=6E-08 W=5E-07 $X=17995 $Y=26070 $D=1
M574 VDD 144 WE VDD P12LL L=6E-08 W=1E-06 $X=18055 $Y=4905 $D=1
M575 639 VSS VDD VDD P12LL L=1E-07 W=4E-07 $X=18080 $Y=20425 $D=1
M576 VDD 105 103 VDD P12LL L=6E-08 W=4E-07 $X=18155 $Y=28025 $D=1
M577 INTCLKX 105 FCKX[5] VDD P12LL L=6E-08 W=1.25E-06 $X=18155 $Y=31220 $D=1
M578 VDD 103 FCKX[5] VDD P12LL L=6E-08 W=1.25E-06 $X=18155 $Y=34780 $D=1
M579 VDD 102 116 VDD P12LL L=6E-08 W=2.5E-06 $X=18210 $Y=11350 $D=1
M580 WE 144 VDD VDD P12LL L=6E-08 W=1E-06 $X=18325 $Y=4905 $D=1
M581 VDD VSS 638 VDD P12LL L=2E-07 W=8E-07 $X=18350 $Y=9190 $D=1
M582 VDD 107 112 VDD P12LL L=2E-07 W=4E-07 $X=18410 $Y=10505 $D=1
M583 113 111 VDD VDD P12LL L=6E-08 W=4E-07 $X=18445 $Y=28025 $D=1
M584 FCKX[4] 111 INTCLKX VDD P12LL L=6E-08 W=1.25E-06 $X=18445 $Y=31220 $D=1
M585 FCKX[4] 113 VDD VDD P12LL L=6E-08 W=1.25E-06 $X=18445 $Y=34780 $D=1
M586 116 102 VDD VDD P12LL L=6E-08 W=2.5E-06 $X=18480 $Y=11350 $D=1
M587 VDD 144 WE VDD P12LL L=6E-08 W=1E-06 $X=18595 $Y=4905 $D=1
M588 114 A[0] 639 VDD P12LL L=6E-08 W=4E-07 $X=18600 $Y=20425 $D=1
M589 115 ACTRCLK 111 VDD P12LL L=6E-08 W=5E-07 $X=18605 $Y=26070 $D=1
M590 VDD 74 115 VDD P12LL L=6E-08 W=1E-06 $X=18735 $Y=21925 $D=1
M591 VDD 111 113 VDD P12LL L=6E-08 W=4E-07 $X=18735 $Y=28025 $D=1
M592 INTCLKX 111 FCKX[4] VDD P12LL L=6E-08 W=1.25E-06 $X=18735 $Y=31220 $D=1
M593 VDD 113 FCKX[4] VDD P12LL L=6E-08 W=1.25E-06 $X=18735 $Y=34780 $D=1
M594 VDD 102 116 VDD P12LL L=6E-08 W=2.5E-06 $X=18750 $Y=11350 $D=1
M595 WE 144 VDD VDD P12LL L=6E-08 W=1E-06 $X=18865 $Y=4905 $D=1
M596 111 ACTRCLK 115 VDD P12LL L=6E-08 W=5E-07 $X=18875 $Y=26070 $D=1
M597 VDD 113 111 VDD P12LL L=3E-07 W=1.2E-07 $X=18985 $Y=27185 $D=1
M598 116 102 VDD VDD P12LL L=6E-08 W=2.5E-06 $X=19020 $Y=11350 $D=1
M599 115 121 VDD VDD P12LL L=6E-08 W=1E-06 $X=19025 $Y=21925 $D=1
M600 113 111 VDD VDD P12LL L=6E-08 W=4E-07 $X=19025 $Y=28025 $D=1
M601 FCKX[4] 111 INTCLKX VDD P12LL L=6E-08 W=1.25E-06 $X=19025 $Y=31220 $D=1
M602 FCKX[4] 113 VDD VDD P12LL L=6E-08 W=1.25E-06 $X=19025 $Y=34780 $D=1
M603 VDD 144 WE VDD P12LL L=6E-08 W=1E-06 $X=19135 $Y=4905 $D=1
M604 115 ACTRCLK 111 VDD P12LL L=6E-08 W=5E-07 $X=19155 $Y=26070 $D=1
M605 120 116 136 VDD P12LL L=6E-08 W=1.25E-06 $X=19200 $Y=9420 $D=1
M606 63 114 VDD VDD P12LL L=6E-08 W=1E-06 $X=19230 $Y=20095 $D=1
M607 VDD 102 116 VDD P12LL L=6E-08 W=2.5E-06 $X=19290 $Y=11350 $D=1
M608 VDD 118 115 VDD P12LL L=6E-08 W=1E-06 $X=19315 $Y=21925 $D=1
M609 VDD 111 113 VDD P12LL L=6E-08 W=4E-07 $X=19315 $Y=28025 $D=1
M610 INTCLKX 111 FCKX[4] VDD P12LL L=6E-08 W=1.25E-06 $X=19315 $Y=31220 $D=1
M611 VDD 113 FCKX[4] VDD P12LL L=6E-08 W=1.25E-06 $X=19315 $Y=34780 $D=1
M612 WE 144 VDD VDD P12LL L=6E-08 W=1E-06 $X=19395 $Y=4905 $D=1
M613 VDD 112 120 VDD P12LL L=6E-08 W=1.25E-06 $X=19470 $Y=9420 $D=1
M614 VDD 114 63 VDD P12LL L=6E-08 W=1E-06 $X=19520 $Y=20095 $D=1
M615 INTCLKX 116 VDD VDD P12LL L=6E-08 W=2.5E-06 $X=19560 $Y=11350 $D=1
M616 124 118 VDD VDD P12LL L=6E-08 W=1E-06 $X=19605 $Y=21925 $D=1
M617 122 123 VDD VDD P12LL L=6E-08 W=4E-07 $X=19605 $Y=28025 $D=1
M618 FCKX[6] 123 INTCLKX VDD P12LL L=6E-08 W=1.25E-06 $X=19605 $Y=31220 $D=1
M619 FCKX[6] 122 VDD VDD P12LL L=6E-08 W=1.25E-06 $X=19605 $Y=34780 $D=1
M620 VDD 144 WE VDD P12LL L=6E-08 W=1E-06 $X=19665 $Y=4905 $D=1
M621 123 122 VDD VDD P12LL L=3E-07 W=1.2E-07 $X=19695 $Y=27185 $D=1
M622 120 112 VDD VDD P12LL L=6E-08 W=1.25E-06 $X=19740 $Y=9420 $D=1
M623 123 ACTRCLK 124 VDD P12LL L=6E-08 W=5E-07 $X=19765 $Y=26070 $D=1
M624 121 63 VDD VDD P12LL L=6E-08 W=1E-06 $X=19810 $Y=20095 $D=1
M625 VDD 116 INTCLKX VDD P12LL L=6E-08 W=2.5E-06 $X=19830 $Y=11350 $D=1
M626 VDD 121 124 VDD P12LL L=6E-08 W=1E-06 $X=19895 $Y=21925 $D=1
M627 VDD 123 122 VDD P12LL L=6E-08 W=4E-07 $X=19895 $Y=28025 $D=1
M628 INTCLKX 123 FCKX[6] VDD P12LL L=6E-08 W=1.25E-06 $X=19895 $Y=31220 $D=1
M629 VDD 122 FCKX[6] VDD P12LL L=6E-08 W=1.25E-06 $X=19895 $Y=34780 $D=1
M630 136 116 120 VDD P12LL L=6E-08 W=1.25E-06 $X=20010 $Y=9420 $D=1
M631 124 ACTRCLK 123 VDD P12LL L=6E-08 W=5E-07 $X=20045 $Y=26070 $D=1
M632 INTCLKX 116 VDD VDD P12LL L=6E-08 W=2.5E-06 $X=20100 $Y=11350 $D=1
M633 VDD 63 121 VDD P12LL L=6E-08 W=1E-06 $X=20100 $Y=20095 $D=1
M634 124 58 VDD VDD P12LL L=6E-08 W=1E-06 $X=20185 $Y=21925 $D=1
M635 122 123 VDD VDD P12LL L=6E-08 W=4E-07 $X=20185 $Y=28025 $D=1
M636 FCKX[6] 123 INTCLKX VDD P12LL L=6E-08 W=1.25E-06 $X=20185 $Y=31220 $D=1
M637 FCKX[6] 122 VDD VDD P12LL L=6E-08 W=1.25E-06 $X=20185 $Y=34780 $D=1
M638 126 WEN VDD VDD P12LL L=6E-08 W=4E-07 $X=20315 $Y=5390 $D=1
M639 123 ACTRCLK 124 VDD P12LL L=6E-08 W=5E-07 $X=20315 $Y=26070 $D=1
M640 VDD 116 INTCLKX VDD P12LL L=6E-08 W=2.5E-06 $X=20370 $Y=11350 $D=1
M641 VDD 123 122 VDD P12LL L=6E-08 W=4E-07 $X=20475 $Y=28025 $D=1
M642 INTCLKX 123 FCKX[6] VDD P12LL L=6E-08 W=1.25E-06 $X=20475 $Y=31220 $D=1
M643 VDD 122 FCKX[6] VDD P12LL L=6E-08 W=1.25E-06 $X=20475 $Y=34780 $D=1
M644 129 136 VDD VDD P12LL L=6E-08 W=1E-06 $X=20610 $Y=9485 $D=1
M645 VDD 136 129 VDD P12LL L=6E-08 W=1E-06 $X=20880 $Y=9485 $D=1
M646 VDD 126 130 VDD P12LL L=3E-07 W=4E-07 $X=20990 $Y=5390 $D=1
M647 129 136 VDD VDD P12LL L=6E-08 W=1E-06 $X=21150 $Y=9485 $D=1
M648 133 130 VDD VDD P12LL L=2E-07 W=4E-07 $X=21580 $Y=5390 $D=1
M649 DCTRCLKX 129 VDD VDD P12LL L=6E-08 W=5E-06 $X=22110 $Y=8750 $D=1
M650 VDD 129 DCTRCLKX VDD P12LL L=6E-08 W=5E-06 $X=22380 $Y=8750 $D=1
M651 134 133 VDD VDD P12LL L=6E-08 W=1E-06 $X=22390 $Y=4985 $D=1
M652 DCTRCLK 136 VDD VDD P12LL L=6E-08 W=5E-06 $X=22650 $Y=8750 $D=1
M653 138 ACTRCLK 134 VDD P12LL L=6E-08 W=1E-06 $X=22660 $Y=4985 $D=1
M654 VDD 136 DCTRCLK VDD P12LL L=6E-08 W=5E-06 $X=22920 $Y=8750 $D=1
M655 ACTRCLK 136 VDD VDD P12LL L=6E-08 W=5E-06 $X=23190 $Y=8750 $D=1
M656 138 140 VDD VDD P12LL L=3E-07 W=1.2E-07 $X=23355 $Y=5460 $D=1
M657 VDD 136 ACTRCLK VDD P12LL L=6E-08 W=5E-06 $X=23460 $Y=8750 $D=1
M658 ACTRCLKX ACTRCLK VDD VDD P12LL L=6E-08 W=5E-06 $X=23730 $Y=8750 $D=1
M659 VDD ACTRCLK ACTRCLKX VDD P12LL L=6E-08 W=5E-06 $X=24000 $Y=8750 $D=1
M660 VDD 138 140 VDD P12LL L=6E-08 W=1E-06 $X=24020 $Y=4985 $D=1
M661 SACK1 116 VDD VDD P12LL L=6E-08 W=5E-06 $X=24270 $Y=8750 $D=1
M662 144 116 VDD VDD P12LL L=6E-08 W=1E-06 $X=24290 $Y=4985 $D=1
M663 VDD 116 SACK1 VDD P12LL L=6E-08 W=5E-06 $X=24540 $Y=8750 $D=1
M664 VDD 140 144 VDD P12LL L=6E-08 W=1E-06 $X=24560 $Y=4985 $D=1
M665 SACK4 141 VDD VDD P12LL L=6E-08 W=5E-06 $X=24810 $Y=8750 $D=1
M666 144 140 VDD VDD P12LL L=6E-08 W=1E-06 $X=24830 $Y=4985 $D=1
M667 VDD 141 SACK4 VDD P12LL L=6E-08 W=5E-06 $X=25080 $Y=8750 $D=1
M668 VDD 116 144 VDD P12LL L=6E-08 W=1E-06 $X=25110 $Y=4985 $D=1
M669 144 116 VDD VDD P12LL L=6E-08 W=1E-06 $X=25390 $Y=4985 $D=1
M670 VDD 140 144 VDD P12LL L=6E-08 W=1E-06 $X=25670 $Y=4985 $D=1
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    S55NLLGDPH_X512Y8D16_BW_LOGIC_BASE_Y8
* View Name:    schematic
************************************************************************

.SUBCKT S55NLLGDPH_X512Y8D16_BW_LOGIC_BASE_Y8 A[7] A[6] A[5] A[4] A[3] A[2] A[1] A[0] ACTRCLK ACTRCLKX
+CEN CLK DCTRCLK DCTRCLKX EMCLK FB FCKX[7] FCKX[6] FCKX[5] FCKX[4]
+FCKX[3] FCKX[2] FCKX[1] FCKX[0] PXA[3] PXA[2] PXA[1] PXA[0] RDE RWL
+S[1] S[0] SACK1 SACK4 VDD VSS WE WEN YX[7] YX[6]
+YX[5] YX[4] YX[3] YX[2] YX[1] YX[0]
XI0 A[0] A[1] A[2] ACTRCLK ACTRCLKX VDD VSS INTCLKX YX[7] YX[6]
+YX[5] YX[4] YX[3] YX[2] YX[1] YX[0] S55NLLGDPH_X512Y8D16_BW_YPREDEC_Y8
XI1 ACTRCLK ACTRCLKX DCTRCLK DCTRCLKX EMCLK FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3]
+FCKX[2] FCKX[1] FCKX[0] PXA[3] PXA[2] PXA[1] PXA[0] RWL SACK1 SACK4
+WE A[7] A[6] A[5] A[4] A[3] CEN CLK FB RDE
+WEN INTCLKX S[1] S[0] VDD VSS S55NLLGDPH_X512Y8D16_BW_LOGIC_BASE
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    S55NLLGDPH_X512Y8D16_BW_ESDA11
* View Name:    schematic
************************************************************************

.SUBCKT S55NLLGDPH_X512Y8D16_BW_ESDA11 A[11] A[10] A[9] A[8] A[7] A[6] A[5] A[4] A[3] A[2]
+A[1] A[0] CEN CLK WEN VDD VSS
MN11 A[11] VSS VSS VSS N12LL W=0.2U L=0.06U M=1
MP11 VDD VDD A[11] VDD P12LL W=0.2U L=0.06U M=1
MN10 A[10] VSS VSS VSS N12LL W=0.2U L=0.06U M=1
MP10 VDD VDD A[10] VDD P12LL W=0.2U L=0.06U M=1
MN9 A[9] VSS VSS VSS N12LL W=0.2U L=0.06U M=1
MP9 VDD VDD A[9] VDD P12LL W=0.2U L=0.06U M=1
MN8 A[8] VSS VSS VSS N12LL W=0.2U L=0.06U M=1
MP8 VDD VDD A[8] VDD P12LL W=0.2U L=0.06U M=1
MN7 A[7] VSS VSS VSS N12LL W=0.2U L=0.06U M=1
MP7 VDD VDD A[7] VDD P12LL W=0.2U L=0.06U M=1
MN6 A[6] VSS VSS VSS N12LL W=0.2U L=0.06U M=1
MP6 VDD VDD A[6] VDD P12LL W=0.2U L=0.06U M=1
MN5 A[5] VSS VSS VSS N12LL W=0.2U L=0.06U M=1
MP5 VDD VDD A[5] VDD P12LL W=0.2U L=0.06U M=1
MN4 A[4] VSS VSS VSS N12LL W=0.2U L=0.06U M=1
MP4 VDD VDD A[4] VDD P12LL W=0.2U L=0.06U M=1
MN3 A[3] VSS VSS VSS N12LL W=0.2U L=0.06U M=1
MP3 VDD VDD A[3] VDD P12LL W=0.2U L=0.06U M=1
MN2 A[2] VSS VSS VSS N12LL W=0.2U L=0.06U M=1
MP2 VDD VDD A[2] VDD P12LL W=0.2U L=0.06U M=1
MN1 A[1] VSS VSS VSS N12LL W=0.2U L=0.06U M=1
MP1 VDD VDD A[1] VDD P12LL W=0.2U L=0.06U M=1
MN0 A[0] VSS VSS VSS N12LL W=0.2U L=0.06U M=1
MP0 VDD VDD A[0] VDD P12LL W=0.2U L=0.06U M=1
MN93 CEN VSS VSS VSS N12LL W=0.2U L=0.06U M=1
MN91 WEN VSS VSS VSS N12LL W=0.2U L=0.06U M=1
MN90 CLK VSS VSS VSS N12LL W=0.2U L=0.06U M=1
MP93 VDD VDD CEN VDD P12LL W=0.2U L=0.06U M=1
MP91 VDD VDD WEN VDD P12LL W=0.2U L=0.06U M=1
MP90 VDD VDD CLK VDD P12LL W=0.2U L=0.06U M=1
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    S55NLLGDPH_X512Y8D16_BW_TIE_LOW_S
* View Name:    schematic
************************************************************************

.SUBCKT S55NLLGDPH_X512Y8D16_BW_TIE_LOW_S PULL0 VSS VDD
MP18 VDD NET2 NET2 VDD P12LL W=2U L=0.06U M=1
MN18 PULL0 NET2 VSS VSS N12LL W=3U L=0.06U M=1
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    S55NLLGDPH_X512Y8D16_BW_TIE_HIGH_S
* View Name:    schematic
************************************************************************

.SUBCKT S55NLLGDPH_X512Y8D16_BW_TIE_HIGH_S PULL1 VSS VDD
MP18 VDD NET2 PULL1 VDD P12LL W=4U L=0.06U M=1
MN18 NET2 NET2 VSS VSS N12LL W=2U L=0.06U M=1
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    S55NLLGDPH_X512Y8D16_BW_OPDEC
* View Name:    schematic
************************************************************************

.SUBCKT S55NLLGDPH_X512Y8D16_BW_OPDEC OP[1] OP[0] S[2] S[1] S[0] VDD VSS
M0 VSS OP[0] 6 VSS N12LL L=6E-08 W=4E-07
M1 8 OP[1] VSS VSS N12LL L=6E-08 W=4E-07
M2 14 6 S[0] VSS N12LL L=6E-08 W=4E-07
M3 VSS 8 14 VSS N12LL L=6E-08 W=4E-07
M4 VSS 8 S[1] VSS N12LL L=6E-08 W=4E-07
M5 VSS 8 S[2] VSS N12LL L=6E-08 W=4E-07
M6 S[2] 6 VSS VSS N12LL L=6E-08 W=4E-07
M9 VDD OP[0] 6 VDD P12LL L=6E-08 W=4E-07
M10 8 OP[1] VDD VDD P12LL L=6E-08 W=4E-07
M11 VDD 6 S[0] VDD P12LL L=6E-08 W=4E-07
M12 S[0] 8 VDD VDD P12LL L=6E-08 W=4E-07
M13 VDD 8 S[1] VDD P12LL L=6E-08 W=4E-07
M14 15 8 S[2] VDD P12LL L=6E-08 W=4E-07
M15 VDD 6 15 VDD P12LL L=6E-08 W=4E-07
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    S55NLLGDPH_X512Y8D16_BW_TIE_LOW_X2
* View Name:    schematic
************************************************************************

.SUBCKT S55NLLGDPH_X512Y8D16_BW_TIE_LOW_X2 PULL0 VSS VDD
MP18 VDD NET2 NET2 VDD P12LL W=0.4U L=0.06U M=1
MN18 PULL0 NET2 VSS VSS N12LL W=1U L=0.06U M=1
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    S55NLLGDPH_X512Y8D16_BW_DISCHARGECELLS
* View Name:    schematic
************************************************************************

.SUBCKT S55NLLGDPH_X512Y8D16_BW_DISCHARGECELLS DUM_BL EMCLK S[2] S[1] S[0] VDD VSS
M0 4 EMCLK DUM_BL VSS DPNPGBHVT L=8.5E-08 W=1E-07
M1 4 EMCLK DUM_BL VSS DPNPGBHVT L=8.5E-08 W=1E-07
M2 4 EMCLK DUM_BL VSS DPNPGBHVT L=8.5E-08 W=1E-07
M3 4 EMCLK DUM_BL VSS DPNPGBHVT L=8.5E-08 W=1E-07
M4 DUM_BL EMCLK 6 VSS DPNPGBHVT L=8.5E-08 W=1E-07
M5 DUM_BL EMCLK 6 VSS DPNPGBHVT L=8.5E-08 W=1E-07
M6 DUM_BL EMCLK 6 VSS DPNPGBHVT L=8.5E-08 W=1E-07
M7 DUM_BL EMCLK 6 VSS DPNPGBHVT L=8.5E-08 W=1E-07
M8 8 EMCLK DUM_BL VSS DPNPGBHVT L=8.5E-08 W=1E-07
M9 8 EMCLK DUM_BL VSS DPNPGBHVT L=8.5E-08 W=1E-07
M10 8 EMCLK DUM_BL VSS DPNPGBHVT L=8.5E-08 W=1E-07
M11 8 EMCLK DUM_BL VSS DPNPGBHVT L=8.5E-08 W=1E-07
M12 DUM_BL EMCLK 10 VSS DPNPGBHVT L=8.5E-08 W=1E-07
M13 DUM_BL EMCLK 10 VSS DPNPGBHVT L=8.5E-08 W=1E-07
M14 DUM_BL EMCLK 10 VSS DPNPGBHVT L=8.5E-08 W=1E-07
M15 DUM_BL EMCLK 10 VSS DPNPGBHVT L=8.5E-08 W=1E-07
M16 10 EMCLK DUM_BL VSS DPNPGBHVT L=8.5E-08 W=1E-07
M17 10 EMCLK DUM_BL VSS DPNPGBHVT L=8.5E-08 W=1E-07
M18 10 EMCLK DUM_BL VSS DPNPGBHVT L=8.5E-08 W=1E-07
M19 10 EMCLK DUM_BL VSS DPNPGBHVT L=8.5E-08 W=1E-07
M20 VSS VDD 4 VSS DPNPDHVT L=7.0E-08 W=3.1E-07
M21 VSS VDD 4 VSS DPNPDHVT L=7.0E-08 W=3.1E-07
M22 VSS VDD 4 VSS DPNPDHVT L=7.0E-08 W=3.1E-07
M23 VSS VDD 4 VSS DPNPDHVT L=7.0E-08 W=3.1E-07
M24 6 S[0] VSS VSS DPNPDHVT L=7.0E-08 W=3.1E-07
M25 6 S[0] VSS VSS DPNPDHVT L=7.0E-08 W=3.1E-07
M26 6 S[0] VSS VSS DPNPDHVT L=7.0E-08 W=3.1E-07
M27 6 S[0] VSS VSS DPNPDHVT L=7.0E-08 W=3.1E-07
M28 VSS S[1] 8 VSS DPNPDHVT L=7.0E-08 W=3.1E-07
M29 VSS S[1] 8 VSS DPNPDHVT L=7.0E-08 W=3.1E-07
M30 VSS S[1] 8 VSS DPNPDHVT L=7.0E-08 W=3.1E-07
M31 VSS S[1] 8 VSS DPNPDHVT L=7.0E-08 W=3.1E-07
M32 10 S[2] VSS VSS DPNPDHVT L=7.0E-08 W=3.1E-07
M33 10 S[2] VSS VSS DPNPDHVT L=7.0E-08 W=3.1E-07
M34 10 S[2] VSS VSS DPNPDHVT L=7.0E-08 W=3.1E-07
M35 10 S[2] VSS VSS DPNPDHVT L=7.0E-08 W=3.1E-07
M36 VSS S[2] 10 VSS DPNPDHVT L=7.0E-08 W=3.1E-07
M37 VSS S[2] 10 VSS DPNPDHVT L=7.0E-08 W=3.1E-07
M38 VSS S[2] 10 VSS DPNPDHVT L=7.0E-08 W=3.1E-07
M39 VSS S[2] 10 VSS DPNPDHVT L=7.0E-08 W=3.1E-07
.ENDS

************************************************************************
* Library Name:  SMIC_MEMORY
* Cell Name:    S55NLLGDPH_X512Y8D16_BW
* View Name:    schematic
************************************************************************

.SUBCKT S55NLLGDPH_X512Y8D16_BW AA[11] AA[10] AA[9] AA[8] AA[7] AA[6] AA[5] AA[4] AA[3] AA[2]
+AA[1] AA[0] AB[11] AB[10] AB[9] AB[8] AB[7] AB[6] AB[5] AB[4]
+AB[3] AB[2] AB[1] AB[0] BWENA[15] BWENA[14] BWENA[13] BWENA[12] BWENA[11] BWENA[10]
+BWENA[9] BWENA[8] BWENA[7] BWENA[6] BWENA[5] BWENA[4] BWENA[3] BWENA[2] BWENA[1] BWENA[0]
+BWENB[15] BWENB[14] BWENB[13] BWENB[12] BWENB[11] BWENB[10] BWENB[9] BWENB[8] BWENB[7] BWENB[6]
+BWENB[5] BWENB[4] BWENB[3] BWENB[2] BWENB[1] BWENB[0] CENA CENB CLKA CLKB
+DA[15] DA[14] DA[13] DA[12] DA[11] DA[10] DA[9] DA[8] DA[7] DA[6]
+DA[5] DA[4] DA[3] DA[2] DA[1] DA[0] DB[15] DB[14] DB[13] DB[12]
+DB[11] DB[10] DB[9] DB[8] DB[7] DB[6] DB[5] DB[4] DB[3] DB[2]
+DB[1] DB[0] QA[15] QA[14] QA[13] QA[12] QA[11] QA[10] QA[9] QA[8]
+QA[7] QA[6] QA[5] QA[4] QA[3] QA[2] QA[1] QA[0] QB[15] QB[14]
+QB[13] QB[12] QB[11] QB[10] QB[9] QB[8] QB[7] QB[6] QB[5] QB[4]
+QB[3] QB[2] QB[1] QB[0] VDD VSS WENA WENB
XI0 EMCLKA STWLA VDD VSS S55NLLGDPH_X512Y8D16_BW_STWL_DEC
XI1 EMCLKB STWLB VDD VSS S55NLLGDPH_X512Y8D16_BW_STWL_DEC
XI2 BWENA[7] BWENA[6] BWENA[5] BWENA[4] BWENA[3] BWENA[2] BWENA[1] BWENA[0] BWENB[7] BWENB[6]
+BWENB[5] BWENB[4] BWENB[3] BWENB[2] BWENB[1] BWENB[0] DCTRCLKA DCTRCLKB DCTRCLKXA DCTRCLKXB
+DA[7] DA[6] DA[5] DA[4] DA[3] DA[2] DA[1] DA[0] DB[7] DB[6]
+DB[5] DB[4] DB[3] DB[2] DB[1] DB[0] DBLA QA[7] QA[6] QA[5]
+QA[4] QA[3] QA[2] QA[1] QA[0] QB[7] QB[6] QB[5] QB[4] QB[3]
+QB[2] QB[1] QB[0] VSS RWLA VSS RWLB SACK1A SACK1B SACK4A
+SACK4B STWLA STWLB VDD VSS WEA WEB WLA[511] WLA[510] WLA[509]
+WLA[508] WLA[507] WLA[506] WLA[505] WLA[504] WLA[503] WLA[502] WLA[501] WLA[500] WLA[499]
+WLA[498] WLA[497] WLA[496] WLA[495] WLA[494] WLA[493] WLA[492] WLA[491] WLA[490] WLA[489]
+WLA[488] WLA[487] WLA[486] WLA[485] WLA[484] WLA[483] WLA[482] WLA[481] WLA[480] WLA[479]
+WLA[478] WLA[477] WLA[476] WLA[475] WLA[474] WLA[473] WLA[472] WLA[471] WLA[470] WLA[469]
+WLA[468] WLA[467] WLA[466] WLA[465] WLA[464] WLA[463] WLA[462] WLA[461] WLA[460] WLA[459]
+WLA[458] WLA[457] WLA[456] WLA[455] WLA[454] WLA[453] WLA[452] WLA[451] WLA[450] WLA[449]
+WLA[448] WLA[447] WLA[446] WLA[445] WLA[444] WLA[443] WLA[442] WLA[441] WLA[440] WLA[439]
+WLA[438] WLA[437] WLA[436] WLA[435] WLA[434] WLA[433] WLA[432] WLA[431] WLA[430] WLA[429]
+WLA[428] WLA[427] WLA[426] WLA[425] WLA[424] WLA[423] WLA[422] WLA[421] WLA[420] WLA[419]
+WLA[418] WLA[417] WLA[416] WLA[415] WLA[414] WLA[413] WLA[412] WLA[411] WLA[410] WLA[409]
+WLA[408] WLA[407] WLA[406] WLA[405] WLA[404] WLA[403] WLA[402] WLA[401] WLA[400] WLA[399]
+WLA[398] WLA[397] WLA[396] WLA[395] WLA[394] WLA[393] WLA[392] WLA[391] WLA[390] WLA[389]
+WLA[388] WLA[387] WLA[386] WLA[385] WLA[384] WLA[383] WLA[382] WLA[381] WLA[380] WLA[379]
+WLA[378] WLA[377] WLA[376] WLA[375] WLA[374] WLA[373] WLA[372] WLA[371] WLA[370] WLA[369]
+WLA[368] WLA[367] WLA[366] WLA[365] WLA[364] WLA[363] WLA[362] WLA[361] WLA[360] WLA[359]
+WLA[358] WLA[357] WLA[356] WLA[355] WLA[354] WLA[353] WLA[352] WLA[351] WLA[350] WLA[349]
+WLA[348] WLA[347] WLA[346] WLA[345] WLA[344] WLA[343] WLA[342] WLA[341] WLA[340] WLA[339]
+WLA[338] WLA[337] WLA[336] WLA[335] WLA[334] WLA[333] WLA[332] WLA[331] WLA[330] WLA[329]
+WLA[328] WLA[327] WLA[326] WLA[325] WLA[324] WLA[323] WLA[322] WLA[321] WLA[320] WLA[319]
+WLA[318] WLA[317] WLA[316] WLA[315] WLA[314] WLA[313] WLA[312] WLA[311] WLA[310] WLA[309]
+WLA[308] WLA[307] WLA[306] WLA[305] WLA[304] WLA[303] WLA[302] WLA[301] WLA[300] WLA[299]
+WLA[298] WLA[297] WLA[296] WLA[295] WLA[294] WLA[293] WLA[292] WLA[291] WLA[290] WLA[289]
+WLA[288] WLA[287] WLA[286] WLA[285] WLA[284] WLA[283] WLA[282] WLA[281] WLA[280] WLA[279]
+WLA[278] WLA[277] WLA[276] WLA[275] WLA[274] WLA[273] WLA[272] WLA[271] WLA[270] WLA[269]
+WLA[268] WLA[267] WLA[266] WLA[265] WLA[264] WLA[263] WLA[262] WLA[261] WLA[260] WLA[259]
+WLA[258] WLA[257] WLA[256] WLA[255] WLA[254] WLA[253] WLA[252] WLA[251] WLA[250] WLA[249]
+WLA[248] WLA[247] WLA[246] WLA[245] WLA[244] WLA[243] WLA[242] WLA[241] WLA[240] WLA[239]
+WLA[238] WLA[237] WLA[236] WLA[235] WLA[234] WLA[233] WLA[232] WLA[231] WLA[230] WLA[229]
+WLA[228] WLA[227] WLA[226] WLA[225] WLA[224] WLA[223] WLA[222] WLA[221] WLA[220] WLA[219]
+WLA[218] WLA[217] WLA[216] WLA[215] WLA[214] WLA[213] WLA[212] WLA[211] WLA[210] WLA[209]
+WLA[208] WLA[207] WLA[206] WLA[205] WLA[204] WLA[203] WLA[202] WLA[201] WLA[200] WLA[199]
+WLA[198] WLA[197] WLA[196] WLA[195] WLA[194] WLA[193] WLA[192] WLA[191] WLA[190] WLA[189]
+WLA[188] WLA[187] WLA[186] WLA[185] WLA[184] WLA[183] WLA[182] WLA[181] WLA[180] WLA[179]
+WLA[178] WLA[177] WLA[176] WLA[175] WLA[174] WLA[173] WLA[172] WLA[171] WLA[170] WLA[169]
+WLA[168] WLA[167] WLA[166] WLA[165] WLA[164] WLA[163] WLA[162] WLA[161] WLA[160] WLA[159]
+WLA[158] WLA[157] WLA[156] WLA[155] WLA[154] WLA[153] WLA[152] WLA[151] WLA[150] WLA[149]
+WLA[148] WLA[147] WLA[146] WLA[145] WLA[144] WLA[143] WLA[142] WLA[141] WLA[140] WLA[139]
+WLA[138] WLA[137] WLA[136] WLA[135] WLA[134] WLA[133] WLA[132] WLA[131] WLA[130] WLA[129]
+WLA[128] WLA[127] WLA[126] WLA[125] WLA[124] WLA[123] WLA[122] WLA[121] WLA[120] WLA[119]
+WLA[118] WLA[117] WLA[116] WLA[115] WLA[114] WLA[113] WLA[112] WLA[111] WLA[110] WLA[109]
+WLA[108] WLA[107] WLA[106] WLA[105] WLA[104] WLA[103] WLA[102] WLA[101] WLA[100] WLA[99]
+WLA[98] WLA[97] WLA[96] WLA[95] WLA[94] WLA[93] WLA[92] WLA[91] WLA[90] WLA[89]
+WLA[88] WLA[87] WLA[86] WLA[85] WLA[84] WLA[83] WLA[82] WLA[81] WLA[80] WLA[79]
+WLA[78] WLA[77] WLA[76] WLA[75] WLA[74] WLA[73] WLA[72] WLA[71] WLA[70] WLA[69]
+WLA[68] WLA[67] WLA[66] WLA[65] WLA[64] WLA[63] WLA[62] WLA[61] WLA[60] WLA[59]
+WLA[58] WLA[57] WLA[56] WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50] WLA[49]
+WLA[48] WLA[47] WLA[46] WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39]
+WLA[38] WLA[37] WLA[36] WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29]
+WLA[28] WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19]
+WLA[18] WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9]
+WLA[8] WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] WLB[511]
+WLB[510] WLB[509] WLB[508] WLB[507] WLB[506] WLB[505] WLB[504] WLB[503] WLB[502] WLB[501]
+WLB[500] WLB[499] WLB[498] WLB[497] WLB[496] WLB[495] WLB[494] WLB[493] WLB[492] WLB[491]
+WLB[490] WLB[489] WLB[488] WLB[487] WLB[486] WLB[485] WLB[484] WLB[483] WLB[482] WLB[481]
+WLB[480] WLB[479] WLB[478] WLB[477] WLB[476] WLB[475] WLB[474] WLB[473] WLB[472] WLB[471]
+WLB[470] WLB[469] WLB[468] WLB[467] WLB[466] WLB[465] WLB[464] WLB[463] WLB[462] WLB[461]
+WLB[460] WLB[459] WLB[458] WLB[457] WLB[456] WLB[455] WLB[454] WLB[453] WLB[452] WLB[451]
+WLB[450] WLB[449] WLB[448] WLB[447] WLB[446] WLB[445] WLB[444] WLB[443] WLB[442] WLB[441]
+WLB[440] WLB[439] WLB[438] WLB[437] WLB[436] WLB[435] WLB[434] WLB[433] WLB[432] WLB[431]
+WLB[430] WLB[429] WLB[428] WLB[427] WLB[426] WLB[425] WLB[424] WLB[423] WLB[422] WLB[421]
+WLB[420] WLB[419] WLB[418] WLB[417] WLB[416] WLB[415] WLB[414] WLB[413] WLB[412] WLB[411]
+WLB[410] WLB[409] WLB[408] WLB[407] WLB[406] WLB[405] WLB[404] WLB[403] WLB[402] WLB[401]
+WLB[400] WLB[399] WLB[398] WLB[397] WLB[396] WLB[395] WLB[394] WLB[393] WLB[392] WLB[391]
+WLB[390] WLB[389] WLB[388] WLB[387] WLB[386] WLB[385] WLB[384] WLB[383] WLB[382] WLB[381]
+WLB[380] WLB[379] WLB[378] WLB[377] WLB[376] WLB[375] WLB[374] WLB[373] WLB[372] WLB[371]
+WLB[370] WLB[369] WLB[368] WLB[367] WLB[366] WLB[365] WLB[364] WLB[363] WLB[362] WLB[361]
+WLB[360] WLB[359] WLB[358] WLB[357] WLB[356] WLB[355] WLB[354] WLB[353] WLB[352] WLB[351]
+WLB[350] WLB[349] WLB[348] WLB[347] WLB[346] WLB[345] WLB[344] WLB[343] WLB[342] WLB[341]
+WLB[340] WLB[339] WLB[338] WLB[337] WLB[336] WLB[335] WLB[334] WLB[333] WLB[332] WLB[331]
+WLB[330] WLB[329] WLB[328] WLB[327] WLB[326] WLB[325] WLB[324] WLB[323] WLB[322] WLB[321]
+WLB[320] WLB[319] WLB[318] WLB[317] WLB[316] WLB[315] WLB[314] WLB[313] WLB[312] WLB[311]
+WLB[310] WLB[309] WLB[308] WLB[307] WLB[306] WLB[305] WLB[304] WLB[303] WLB[302] WLB[301]
+WLB[300] WLB[299] WLB[298] WLB[297] WLB[296] WLB[295] WLB[294] WLB[293] WLB[292] WLB[291]
+WLB[290] WLB[289] WLB[288] WLB[287] WLB[286] WLB[285] WLB[284] WLB[283] WLB[282] WLB[281]
+WLB[280] WLB[279] WLB[278] WLB[277] WLB[276] WLB[275] WLB[274] WLB[273] WLB[272] WLB[271]
+WLB[270] WLB[269] WLB[268] WLB[267] WLB[266] WLB[265] WLB[264] WLB[263] WLB[262] WLB[261]
+WLB[260] WLB[259] WLB[258] WLB[257] WLB[256] WLB[255] WLB[254] WLB[253] WLB[252] WLB[251]
+WLB[250] WLB[249] WLB[248] WLB[247] WLB[246] WLB[245] WLB[244] WLB[243] WLB[242] WLB[241]
+WLB[240] WLB[239] WLB[238] WLB[237] WLB[236] WLB[235] WLB[234] WLB[233] WLB[232] WLB[231]
+WLB[230] WLB[229] WLB[228] WLB[227] WLB[226] WLB[225] WLB[224] WLB[223] WLB[222] WLB[221]
+WLB[220] WLB[219] WLB[218] WLB[217] WLB[216] WLB[215] WLB[214] WLB[213] WLB[212] WLB[211]
+WLB[210] WLB[209] WLB[208] WLB[207] WLB[206] WLB[205] WLB[204] WLB[203] WLB[202] WLB[201]
+WLB[200] WLB[199] WLB[198] WLB[197] WLB[196] WLB[195] WLB[194] WLB[193] WLB[192] WLB[191]
+WLB[190] WLB[189] WLB[188] WLB[187] WLB[186] WLB[185] WLB[184] WLB[183] WLB[182] WLB[181]
+WLB[180] WLB[179] WLB[178] WLB[177] WLB[176] WLB[175] WLB[174] WLB[173] WLB[172] WLB[171]
+WLB[170] WLB[169] WLB[168] WLB[167] WLB[166] WLB[165] WLB[164] WLB[163] WLB[162] WLB[161]
+WLB[160] WLB[159] WLB[158] WLB[157] WLB[156] WLB[155] WLB[154] WLB[153] WLB[152] WLB[151]
+WLB[150] WLB[149] WLB[148] WLB[147] WLB[146] WLB[145] WLB[144] WLB[143] WLB[142] WLB[141]
+WLB[140] WLB[139] WLB[138] WLB[137] WLB[136] WLB[135] WLB[134] WLB[133] WLB[132] WLB[131]
+WLB[130] WLB[129] WLB[128] WLB[127] WLB[126] WLB[125] WLB[124] WLB[123] WLB[122] WLB[121]
+WLB[120] WLB[119] WLB[118] WLB[117] WLB[116] WLB[115] WLB[114] WLB[113] WLB[112] WLB[111]
+WLB[110] WLB[109] WLB[108] WLB[107] WLB[106] WLB[105] WLB[104] WLB[103] WLB[102] WLB[101]
+WLB[100] WLB[99] WLB[98] WLB[97] WLB[96] WLB[95] WLB[94] WLB[93] WLB[92] WLB[91]
+WLB[90] WLB[89] WLB[88] WLB[87] WLB[86] WLB[85] WLB[84] WLB[83] WLB[82] WLB[81]
+WLB[80] WLB[79] WLB[78] WLB[77] WLB[76] WLB[75] WLB[74] WLB[73] WLB[72] WLB[71]
+WLB[70] WLB[69] WLB[68] WLB[67] WLB[66] WLB[65] WLB[64] WLB[63] WLB[62] WLB[61]
+WLB[60] WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54] WLB[53] WLB[52] WLB[51]
+WLB[50] WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44] WLB[43] WLB[42] WLB[41]
+WLB[40] WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34] WLB[33] WLB[32] WLB[31]
+WLB[30] WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24] WLB[23] WLB[22] WLB[21]
+WLB[20] WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14] WLB[13] WLB[12] WLB[11]
+WLB[10] WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4] WLB[3] WLB[2] WLB[1]
+WLB[0] YXA[7] YXA[6] YXA[5] YXA[4] YXA[3] YXA[2] YXA[1] YXA[0] YXB[7]
+YXB[6] YXB[5] YXB[4] YXB[3] YXB[2] YXB[1] YXB[0] S55NLLGDPH_X512Y8D16_BW_Y512X8CELLX8_BW_LEFT
XI3 BWENA[15] BWENA[14] BWENA[13] BWENA[12] BWENA[11] BWENA[10] BWENA[9] BWENA[8] BWENB[15] BWENB[14]
+BWENB[13] BWENB[12] BWENB[11] BWENB[10] BWENB[9] BWENB[8] DCTRCLKA DCTRCLKB DCTRCLKXA DCTRCLKXB
+DA[15] DA[14] DA[13] DA[12] DA[11] DA[10] DA[9] DA[8] DB[15] DB[14]
+DB[13] DB[12] DB[11] DB[10] DB[9] DB[8] DBLB QA[15] QA[14] QA[13]
+QA[12] QA[11] QA[10] QA[9] QA[8] QB[15] QB[14] QB[13] QB[12] QB[11]
+QB[10] QB[9] QB[8] VSS RWLA VSS RWLB SACK1A SACK1B SACK4A
+SACK4B STWLA STWLB VDD VSS WEA WEB WLA[511] WLA[510] WLA[509]
+WLA[508] WLA[507] WLA[506] WLA[505] WLA[504] WLA[503] WLA[502] WLA[501] WLA[500] WLA[499]
+WLA[498] WLA[497] WLA[496] WLA[495] WLA[494] WLA[493] WLA[492] WLA[491] WLA[490] WLA[489]
+WLA[488] WLA[487] WLA[486] WLA[485] WLA[484] WLA[483] WLA[482] WLA[481] WLA[480] WLA[479]
+WLA[478] WLA[477] WLA[476] WLA[475] WLA[474] WLA[473] WLA[472] WLA[471] WLA[470] WLA[469]
+WLA[468] WLA[467] WLA[466] WLA[465] WLA[464] WLA[463] WLA[462] WLA[461] WLA[460] WLA[459]
+WLA[458] WLA[457] WLA[456] WLA[455] WLA[454] WLA[453] WLA[452] WLA[451] WLA[450] WLA[449]
+WLA[448] WLA[447] WLA[446] WLA[445] WLA[444] WLA[443] WLA[442] WLA[441] WLA[440] WLA[439]
+WLA[438] WLA[437] WLA[436] WLA[435] WLA[434] WLA[433] WLA[432] WLA[431] WLA[430] WLA[429]
+WLA[428] WLA[427] WLA[426] WLA[425] WLA[424] WLA[423] WLA[422] WLA[421] WLA[420] WLA[419]
+WLA[418] WLA[417] WLA[416] WLA[415] WLA[414] WLA[413] WLA[412] WLA[411] WLA[410] WLA[409]
+WLA[408] WLA[407] WLA[406] WLA[405] WLA[404] WLA[403] WLA[402] WLA[401] WLA[400] WLA[399]
+WLA[398] WLA[397] WLA[396] WLA[395] WLA[394] WLA[393] WLA[392] WLA[391] WLA[390] WLA[389]
+WLA[388] WLA[387] WLA[386] WLA[385] WLA[384] WLA[383] WLA[382] WLA[381] WLA[380] WLA[379]
+WLA[378] WLA[377] WLA[376] WLA[375] WLA[374] WLA[373] WLA[372] WLA[371] WLA[370] WLA[369]
+WLA[368] WLA[367] WLA[366] WLA[365] WLA[364] WLA[363] WLA[362] WLA[361] WLA[360] WLA[359]
+WLA[358] WLA[357] WLA[356] WLA[355] WLA[354] WLA[353] WLA[352] WLA[351] WLA[350] WLA[349]
+WLA[348] WLA[347] WLA[346] WLA[345] WLA[344] WLA[343] WLA[342] WLA[341] WLA[340] WLA[339]
+WLA[338] WLA[337] WLA[336] WLA[335] WLA[334] WLA[333] WLA[332] WLA[331] WLA[330] WLA[329]
+WLA[328] WLA[327] WLA[326] WLA[325] WLA[324] WLA[323] WLA[322] WLA[321] WLA[320] WLA[319]
+WLA[318] WLA[317] WLA[316] WLA[315] WLA[314] WLA[313] WLA[312] WLA[311] WLA[310] WLA[309]
+WLA[308] WLA[307] WLA[306] WLA[305] WLA[304] WLA[303] WLA[302] WLA[301] WLA[300] WLA[299]
+WLA[298] WLA[297] WLA[296] WLA[295] WLA[294] WLA[293] WLA[292] WLA[291] WLA[290] WLA[289]
+WLA[288] WLA[287] WLA[286] WLA[285] WLA[284] WLA[283] WLA[282] WLA[281] WLA[280] WLA[279]
+WLA[278] WLA[277] WLA[276] WLA[275] WLA[274] WLA[273] WLA[272] WLA[271] WLA[270] WLA[269]
+WLA[268] WLA[267] WLA[266] WLA[265] WLA[264] WLA[263] WLA[262] WLA[261] WLA[260] WLA[259]
+WLA[258] WLA[257] WLA[256] WLA[255] WLA[254] WLA[253] WLA[252] WLA[251] WLA[250] WLA[249]
+WLA[248] WLA[247] WLA[246] WLA[245] WLA[244] WLA[243] WLA[242] WLA[241] WLA[240] WLA[239]
+WLA[238] WLA[237] WLA[236] WLA[235] WLA[234] WLA[233] WLA[232] WLA[231] WLA[230] WLA[229]
+WLA[228] WLA[227] WLA[226] WLA[225] WLA[224] WLA[223] WLA[222] WLA[221] WLA[220] WLA[219]
+WLA[218] WLA[217] WLA[216] WLA[215] WLA[214] WLA[213] WLA[212] WLA[211] WLA[210] WLA[209]
+WLA[208] WLA[207] WLA[206] WLA[205] WLA[204] WLA[203] WLA[202] WLA[201] WLA[200] WLA[199]
+WLA[198] WLA[197] WLA[196] WLA[195] WLA[194] WLA[193] WLA[192] WLA[191] WLA[190] WLA[189]
+WLA[188] WLA[187] WLA[186] WLA[185] WLA[184] WLA[183] WLA[182] WLA[181] WLA[180] WLA[179]
+WLA[178] WLA[177] WLA[176] WLA[175] WLA[174] WLA[173] WLA[172] WLA[171] WLA[170] WLA[169]
+WLA[168] WLA[167] WLA[166] WLA[165] WLA[164] WLA[163] WLA[162] WLA[161] WLA[160] WLA[159]
+WLA[158] WLA[157] WLA[156] WLA[155] WLA[154] WLA[153] WLA[152] WLA[151] WLA[150] WLA[149]
+WLA[148] WLA[147] WLA[146] WLA[145] WLA[144] WLA[143] WLA[142] WLA[141] WLA[140] WLA[139]
+WLA[138] WLA[137] WLA[136] WLA[135] WLA[134] WLA[133] WLA[132] WLA[131] WLA[130] WLA[129]
+WLA[128] WLA[127] WLA[126] WLA[125] WLA[124] WLA[123] WLA[122] WLA[121] WLA[120] WLA[119]
+WLA[118] WLA[117] WLA[116] WLA[115] WLA[114] WLA[113] WLA[112] WLA[111] WLA[110] WLA[109]
+WLA[108] WLA[107] WLA[106] WLA[105] WLA[104] WLA[103] WLA[102] WLA[101] WLA[100] WLA[99]
+WLA[98] WLA[97] WLA[96] WLA[95] WLA[94] WLA[93] WLA[92] WLA[91] WLA[90] WLA[89]
+WLA[88] WLA[87] WLA[86] WLA[85] WLA[84] WLA[83] WLA[82] WLA[81] WLA[80] WLA[79]
+WLA[78] WLA[77] WLA[76] WLA[75] WLA[74] WLA[73] WLA[72] WLA[71] WLA[70] WLA[69]
+WLA[68] WLA[67] WLA[66] WLA[65] WLA[64] WLA[63] WLA[62] WLA[61] WLA[60] WLA[59]
+WLA[58] WLA[57] WLA[56] WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50] WLA[49]
+WLA[48] WLA[47] WLA[46] WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39]
+WLA[38] WLA[37] WLA[36] WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29]
+WLA[28] WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19]
+WLA[18] WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9]
+WLA[8] WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] WLB[511]
+WLB[510] WLB[509] WLB[508] WLB[507] WLB[506] WLB[505] WLB[504] WLB[503] WLB[502] WLB[501]
+WLB[500] WLB[499] WLB[498] WLB[497] WLB[496] WLB[495] WLB[494] WLB[493] WLB[492] WLB[491]
+WLB[490] WLB[489] WLB[488] WLB[487] WLB[486] WLB[485] WLB[484] WLB[483] WLB[482] WLB[481]
+WLB[480] WLB[479] WLB[478] WLB[477] WLB[476] WLB[475] WLB[474] WLB[473] WLB[472] WLB[471]
+WLB[470] WLB[469] WLB[468] WLB[467] WLB[466] WLB[465] WLB[464] WLB[463] WLB[462] WLB[461]
+WLB[460] WLB[459] WLB[458] WLB[457] WLB[456] WLB[455] WLB[454] WLB[453] WLB[452] WLB[451]
+WLB[450] WLB[449] WLB[448] WLB[447] WLB[446] WLB[445] WLB[444] WLB[443] WLB[442] WLB[441]
+WLB[440] WLB[439] WLB[438] WLB[437] WLB[436] WLB[435] WLB[434] WLB[433] WLB[432] WLB[431]
+WLB[430] WLB[429] WLB[428] WLB[427] WLB[426] WLB[425] WLB[424] WLB[423] WLB[422] WLB[421]
+WLB[420] WLB[419] WLB[418] WLB[417] WLB[416] WLB[415] WLB[414] WLB[413] WLB[412] WLB[411]
+WLB[410] WLB[409] WLB[408] WLB[407] WLB[406] WLB[405] WLB[404] WLB[403] WLB[402] WLB[401]
+WLB[400] WLB[399] WLB[398] WLB[397] WLB[396] WLB[395] WLB[394] WLB[393] WLB[392] WLB[391]
+WLB[390] WLB[389] WLB[388] WLB[387] WLB[386] WLB[385] WLB[384] WLB[383] WLB[382] WLB[381]
+WLB[380] WLB[379] WLB[378] WLB[377] WLB[376] WLB[375] WLB[374] WLB[373] WLB[372] WLB[371]
+WLB[370] WLB[369] WLB[368] WLB[367] WLB[366] WLB[365] WLB[364] WLB[363] WLB[362] WLB[361]
+WLB[360] WLB[359] WLB[358] WLB[357] WLB[356] WLB[355] WLB[354] WLB[353] WLB[352] WLB[351]
+WLB[350] WLB[349] WLB[348] WLB[347] WLB[346] WLB[345] WLB[344] WLB[343] WLB[342] WLB[341]
+WLB[340] WLB[339] WLB[338] WLB[337] WLB[336] WLB[335] WLB[334] WLB[333] WLB[332] WLB[331]
+WLB[330] WLB[329] WLB[328] WLB[327] WLB[326] WLB[325] WLB[324] WLB[323] WLB[322] WLB[321]
+WLB[320] WLB[319] WLB[318] WLB[317] WLB[316] WLB[315] WLB[314] WLB[313] WLB[312] WLB[311]
+WLB[310] WLB[309] WLB[308] WLB[307] WLB[306] WLB[305] WLB[304] WLB[303] WLB[302] WLB[301]
+WLB[300] WLB[299] WLB[298] WLB[297] WLB[296] WLB[295] WLB[294] WLB[293] WLB[292] WLB[291]
+WLB[290] WLB[289] WLB[288] WLB[287] WLB[286] WLB[285] WLB[284] WLB[283] WLB[282] WLB[281]
+WLB[280] WLB[279] WLB[278] WLB[277] WLB[276] WLB[275] WLB[274] WLB[273] WLB[272] WLB[271]
+WLB[270] WLB[269] WLB[268] WLB[267] WLB[266] WLB[265] WLB[264] WLB[263] WLB[262] WLB[261]
+WLB[260] WLB[259] WLB[258] WLB[257] WLB[256] WLB[255] WLB[254] WLB[253] WLB[252] WLB[251]
+WLB[250] WLB[249] WLB[248] WLB[247] WLB[246] WLB[245] WLB[244] WLB[243] WLB[242] WLB[241]
+WLB[240] WLB[239] WLB[238] WLB[237] WLB[236] WLB[235] WLB[234] WLB[233] WLB[232] WLB[231]
+WLB[230] WLB[229] WLB[228] WLB[227] WLB[226] WLB[225] WLB[224] WLB[223] WLB[222] WLB[221]
+WLB[220] WLB[219] WLB[218] WLB[217] WLB[216] WLB[215] WLB[214] WLB[213] WLB[212] WLB[211]
+WLB[210] WLB[209] WLB[208] WLB[207] WLB[206] WLB[205] WLB[204] WLB[203] WLB[202] WLB[201]
+WLB[200] WLB[199] WLB[198] WLB[197] WLB[196] WLB[195] WLB[194] WLB[193] WLB[192] WLB[191]
+WLB[190] WLB[189] WLB[188] WLB[187] WLB[186] WLB[185] WLB[184] WLB[183] WLB[182] WLB[181]
+WLB[180] WLB[179] WLB[178] WLB[177] WLB[176] WLB[175] WLB[174] WLB[173] WLB[172] WLB[171]
+WLB[170] WLB[169] WLB[168] WLB[167] WLB[166] WLB[165] WLB[164] WLB[163] WLB[162] WLB[161]
+WLB[160] WLB[159] WLB[158] WLB[157] WLB[156] WLB[155] WLB[154] WLB[153] WLB[152] WLB[151]
+WLB[150] WLB[149] WLB[148] WLB[147] WLB[146] WLB[145] WLB[144] WLB[143] WLB[142] WLB[141]
+WLB[140] WLB[139] WLB[138] WLB[137] WLB[136] WLB[135] WLB[134] WLB[133] WLB[132] WLB[131]
+WLB[130] WLB[129] WLB[128] WLB[127] WLB[126] WLB[125] WLB[124] WLB[123] WLB[122] WLB[121]
+WLB[120] WLB[119] WLB[118] WLB[117] WLB[116] WLB[115] WLB[114] WLB[113] WLB[112] WLB[111]
+WLB[110] WLB[109] WLB[108] WLB[107] WLB[106] WLB[105] WLB[104] WLB[103] WLB[102] WLB[101]
+WLB[100] WLB[99] WLB[98] WLB[97] WLB[96] WLB[95] WLB[94] WLB[93] WLB[92] WLB[91]
+WLB[90] WLB[89] WLB[88] WLB[87] WLB[86] WLB[85] WLB[84] WLB[83] WLB[82] WLB[81]
+WLB[80] WLB[79] WLB[78] WLB[77] WLB[76] WLB[75] WLB[74] WLB[73] WLB[72] WLB[71]
+WLB[70] WLB[69] WLB[68] WLB[67] WLB[66] WLB[65] WLB[64] WLB[63] WLB[62] WLB[61]
+WLB[60] WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54] WLB[53] WLB[52] WLB[51]
+WLB[50] WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44] WLB[43] WLB[42] WLB[41]
+WLB[40] WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34] WLB[33] WLB[32] WLB[31]
+WLB[30] WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24] WLB[23] WLB[22] WLB[21]
+WLB[20] WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14] WLB[13] WLB[12] WLB[11]
+WLB[10] WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4] WLB[3] WLB[2] WLB[1]
+WLB[0] YXA[7] YXA[6] YXA[5] YXA[4] YXA[3] YXA[2] YXA[1] YXA[0] YXB[7]
+YXB[6] YXB[5] YXB[4] YXB[3] YXB[2] YXB[1] YXB[0] S55NLLGDPH_X512Y8D16_BW_Y512X8CELLX8_BW_RIGHT
XI4 FCKXA[7] FCKXA[6] FCKXA[5] FCKXA[4] FCKXA[3] FCKXA[2] FCKXA[1] FCKXA[0] PXAA[3] PXAA[2]
+PXAA[1] PXAA[0] PXBA[3] PXBA[2] PXBA[1] PXBA[0] PXCA[3] PXCA[2] PXCA[1] PXCA[0]
+VDD VSS WLA[511] WLA[510] WLA[509] WLA[508] WLA[507] WLA[506] WLA[505] WLA[504]
+WLA[503] WLA[502] WLA[501] WLA[500] WLA[499] WLA[498] WLA[497] WLA[496] WLA[495] WLA[494]
+WLA[493] WLA[492] WLA[491] WLA[490] WLA[489] WLA[488] WLA[487] WLA[486] WLA[485] WLA[484]
+WLA[483] WLA[482] WLA[481] WLA[480] WLA[479] WLA[478] WLA[477] WLA[476] WLA[475] WLA[474]
+WLA[473] WLA[472] WLA[471] WLA[470] WLA[469] WLA[468] WLA[467] WLA[466] WLA[465] WLA[464]
+WLA[463] WLA[462] WLA[461] WLA[460] WLA[459] WLA[458] WLA[457] WLA[456] WLA[455] WLA[454]
+WLA[453] WLA[452] WLA[451] WLA[450] WLA[449] WLA[448] WLA[447] WLA[446] WLA[445] WLA[444]
+WLA[443] WLA[442] WLA[441] WLA[440] WLA[439] WLA[438] WLA[437] WLA[436] WLA[435] WLA[434]
+WLA[433] WLA[432] WLA[431] WLA[430] WLA[429] WLA[428] WLA[427] WLA[426] WLA[425] WLA[424]
+WLA[423] WLA[422] WLA[421] WLA[420] WLA[419] WLA[418] WLA[417] WLA[416] WLA[415] WLA[414]
+WLA[413] WLA[412] WLA[411] WLA[410] WLA[409] WLA[408] WLA[407] WLA[406] WLA[405] WLA[404]
+WLA[403] WLA[402] WLA[401] WLA[400] WLA[399] WLA[398] WLA[397] WLA[396] WLA[395] WLA[394]
+WLA[393] WLA[392] WLA[391] WLA[390] WLA[389] WLA[388] WLA[387] WLA[386] WLA[385] WLA[384]
+WLA[383] WLA[382] WLA[381] WLA[380] WLA[379] WLA[378] WLA[377] WLA[376] WLA[375] WLA[374]
+WLA[373] WLA[372] WLA[371] WLA[370] WLA[369] WLA[368] WLA[367] WLA[366] WLA[365] WLA[364]
+WLA[363] WLA[362] WLA[361] WLA[360] WLA[359] WLA[358] WLA[357] WLA[356] WLA[355] WLA[354]
+WLA[353] WLA[352] WLA[351] WLA[350] WLA[349] WLA[348] WLA[347] WLA[346] WLA[345] WLA[344]
+WLA[343] WLA[342] WLA[341] WLA[340] WLA[339] WLA[338] WLA[337] WLA[336] WLA[335] WLA[334]
+WLA[333] WLA[332] WLA[331] WLA[330] WLA[329] WLA[328] WLA[327] WLA[326] WLA[325] WLA[324]
+WLA[323] WLA[322] WLA[321] WLA[320] WLA[319] WLA[318] WLA[317] WLA[316] WLA[315] WLA[314]
+WLA[313] WLA[312] WLA[311] WLA[310] WLA[309] WLA[308] WLA[307] WLA[306] WLA[305] WLA[304]
+WLA[303] WLA[302] WLA[301] WLA[300] WLA[299] WLA[298] WLA[297] WLA[296] WLA[295] WLA[294]
+WLA[293] WLA[292] WLA[291] WLA[290] WLA[289] WLA[288] WLA[287] WLA[286] WLA[285] WLA[284]
+WLA[283] WLA[282] WLA[281] WLA[280] WLA[279] WLA[278] WLA[277] WLA[276] WLA[275] WLA[274]
+WLA[273] WLA[272] WLA[271] WLA[270] WLA[269] WLA[268] WLA[267] WLA[266] WLA[265] WLA[264]
+WLA[263] WLA[262] WLA[261] WLA[260] WLA[259] WLA[258] WLA[257] WLA[256] WLA[255] WLA[254]
+WLA[253] WLA[252] WLA[251] WLA[250] WLA[249] WLA[248] WLA[247] WLA[246] WLA[245] WLA[244]
+WLA[243] WLA[242] WLA[241] WLA[240] WLA[239] WLA[238] WLA[237] WLA[236] WLA[235] WLA[234]
+WLA[233] WLA[232] WLA[231] WLA[230] WLA[229] WLA[228] WLA[227] WLA[226] WLA[225] WLA[224]
+WLA[223] WLA[222] WLA[221] WLA[220] WLA[219] WLA[218] WLA[217] WLA[216] WLA[215] WLA[214]
+WLA[213] WLA[212] WLA[211] WLA[210] WLA[209] WLA[208] WLA[207] WLA[206] WLA[205] WLA[204]
+WLA[203] WLA[202] WLA[201] WLA[200] WLA[199] WLA[198] WLA[197] WLA[196] WLA[195] WLA[194]
+WLA[193] WLA[192] WLA[191] WLA[190] WLA[189] WLA[188] WLA[187] WLA[186] WLA[185] WLA[184]
+WLA[183] WLA[182] WLA[181] WLA[180] WLA[179] WLA[178] WLA[177] WLA[176] WLA[175] WLA[174]
+WLA[173] WLA[172] WLA[171] WLA[170] WLA[169] WLA[168] WLA[167] WLA[166] WLA[165] WLA[164]
+WLA[163] WLA[162] WLA[161] WLA[160] WLA[159] WLA[158] WLA[157] WLA[156] WLA[155] WLA[154]
+WLA[153] WLA[152] WLA[151] WLA[150] WLA[149] WLA[148] WLA[147] WLA[146] WLA[145] WLA[144]
+WLA[143] WLA[142] WLA[141] WLA[140] WLA[139] WLA[138] WLA[137] WLA[136] WLA[135] WLA[134]
+WLA[133] WLA[132] WLA[131] WLA[130] WLA[129] WLA[128] WLA[127] WLA[126] WLA[125] WLA[124]
+WLA[123] WLA[122] WLA[121] WLA[120] WLA[119] WLA[118] WLA[117] WLA[116] WLA[115] WLA[114]
+WLA[113] WLA[112] WLA[111] WLA[110] WLA[109] WLA[108] WLA[107] WLA[106] WLA[105] WLA[104]
+WLA[103] WLA[102] WLA[101] WLA[100] WLA[99] WLA[98] WLA[97] WLA[96] WLA[95] WLA[94]
+WLA[93] WLA[92] WLA[91] WLA[90] WLA[89] WLA[88] WLA[87] WLA[86] WLA[85] WLA[84]
+WLA[83] WLA[82] WLA[81] WLA[80] WLA[79] WLA[78] WLA[77] WLA[76] WLA[75] WLA[74]
+WLA[73] WLA[72] WLA[71] WLA[70] WLA[69] WLA[68] WLA[67] WLA[66] WLA[65] WLA[64]
+WLA[63] WLA[62] WLA[61] WLA[60] WLA[59] WLA[58] WLA[57] WLA[56] WLA[55] WLA[54]
+WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48] WLA[47] WLA[46] WLA[45] WLA[44]
+WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38] WLA[37] WLA[36] WLA[35] WLA[34]
+WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28] WLA[27] WLA[26] WLA[25] WLA[24]
+WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18] WLA[17] WLA[16] WLA[15] WLA[14]
+WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8] WLA[7] WLA[6] WLA[5] WLA[4]
+WLA[3] WLA[2] WLA[1] WLA[0] S55NLLGDPH_X512Y8D16_BW_XDEC64
XI5 FCKXB[7] FCKXB[6] FCKXB[5] FCKXB[4] FCKXB[3] FCKXB[2] FCKXB[1] FCKXB[0] PXAB[3] PXAB[2]
+PXAB[1] PXAB[0] PXBB[3] PXBB[2] PXBB[1] PXBB[0] PXCB[3] PXCB[2] PXCB[1] PXCB[0]
+VDD VSS WLB[511] WLB[510] WLB[509] WLB[508] WLB[507] WLB[506] WLB[505] WLB[504]
+WLB[503] WLB[502] WLB[501] WLB[500] WLB[499] WLB[498] WLB[497] WLB[496] WLB[495] WLB[494]
+WLB[493] WLB[492] WLB[491] WLB[490] WLB[489] WLB[488] WLB[487] WLB[486] WLB[485] WLB[484]
+WLB[483] WLB[482] WLB[481] WLB[480] WLB[479] WLB[478] WLB[477] WLB[476] WLB[475] WLB[474]
+WLB[473] WLB[472] WLB[471] WLB[470] WLB[469] WLB[468] WLB[467] WLB[466] WLB[465] WLB[464]
+WLB[463] WLB[462] WLB[461] WLB[460] WLB[459] WLB[458] WLB[457] WLB[456] WLB[455] WLB[454]
+WLB[453] WLB[452] WLB[451] WLB[450] WLB[449] WLB[448] WLB[447] WLB[446] WLB[445] WLB[444]
+WLB[443] WLB[442] WLB[441] WLB[440] WLB[439] WLB[438] WLB[437] WLB[436] WLB[435] WLB[434]
+WLB[433] WLB[432] WLB[431] WLB[430] WLB[429] WLB[428] WLB[427] WLB[426] WLB[425] WLB[424]
+WLB[423] WLB[422] WLB[421] WLB[420] WLB[419] WLB[418] WLB[417] WLB[416] WLB[415] WLB[414]
+WLB[413] WLB[412] WLB[411] WLB[410] WLB[409] WLB[408] WLB[407] WLB[406] WLB[405] WLB[404]
+WLB[403] WLB[402] WLB[401] WLB[400] WLB[399] WLB[398] WLB[397] WLB[396] WLB[395] WLB[394]
+WLB[393] WLB[392] WLB[391] WLB[390] WLB[389] WLB[388] WLB[387] WLB[386] WLB[385] WLB[384]
+WLB[383] WLB[382] WLB[381] WLB[380] WLB[379] WLB[378] WLB[377] WLB[376] WLB[375] WLB[374]
+WLB[373] WLB[372] WLB[371] WLB[370] WLB[369] WLB[368] WLB[367] WLB[366] WLB[365] WLB[364]
+WLB[363] WLB[362] WLB[361] WLB[360] WLB[359] WLB[358] WLB[357] WLB[356] WLB[355] WLB[354]
+WLB[353] WLB[352] WLB[351] WLB[350] WLB[349] WLB[348] WLB[347] WLB[346] WLB[345] WLB[344]
+WLB[343] WLB[342] WLB[341] WLB[340] WLB[339] WLB[338] WLB[337] WLB[336] WLB[335] WLB[334]
+WLB[333] WLB[332] WLB[331] WLB[330] WLB[329] WLB[328] WLB[327] WLB[326] WLB[325] WLB[324]
+WLB[323] WLB[322] WLB[321] WLB[320] WLB[319] WLB[318] WLB[317] WLB[316] WLB[315] WLB[314]
+WLB[313] WLB[312] WLB[311] WLB[310] WLB[309] WLB[308] WLB[307] WLB[306] WLB[305] WLB[304]
+WLB[303] WLB[302] WLB[301] WLB[300] WLB[299] WLB[298] WLB[297] WLB[296] WLB[295] WLB[294]
+WLB[293] WLB[292] WLB[291] WLB[290] WLB[289] WLB[288] WLB[287] WLB[286] WLB[285] WLB[284]
+WLB[283] WLB[282] WLB[281] WLB[280] WLB[279] WLB[278] WLB[277] WLB[276] WLB[275] WLB[274]
+WLB[273] WLB[272] WLB[271] WLB[270] WLB[269] WLB[268] WLB[267] WLB[266] WLB[265] WLB[264]
+WLB[263] WLB[262] WLB[261] WLB[260] WLB[259] WLB[258] WLB[257] WLB[256] WLB[255] WLB[254]
+WLB[253] WLB[252] WLB[251] WLB[250] WLB[249] WLB[248] WLB[247] WLB[246] WLB[245] WLB[244]
+WLB[243] WLB[242] WLB[241] WLB[240] WLB[239] WLB[238] WLB[237] WLB[236] WLB[235] WLB[234]
+WLB[233] WLB[232] WLB[231] WLB[230] WLB[229] WLB[228] WLB[227] WLB[226] WLB[225] WLB[224]
+WLB[223] WLB[222] WLB[221] WLB[220] WLB[219] WLB[218] WLB[217] WLB[216] WLB[215] WLB[214]
+WLB[213] WLB[212] WLB[211] WLB[210] WLB[209] WLB[208] WLB[207] WLB[206] WLB[205] WLB[204]
+WLB[203] WLB[202] WLB[201] WLB[200] WLB[199] WLB[198] WLB[197] WLB[196] WLB[195] WLB[194]
+WLB[193] WLB[192] WLB[191] WLB[190] WLB[189] WLB[188] WLB[187] WLB[186] WLB[185] WLB[184]
+WLB[183] WLB[182] WLB[181] WLB[180] WLB[179] WLB[178] WLB[177] WLB[176] WLB[175] WLB[174]
+WLB[173] WLB[172] WLB[171] WLB[170] WLB[169] WLB[168] WLB[167] WLB[166] WLB[165] WLB[164]
+WLB[163] WLB[162] WLB[161] WLB[160] WLB[159] WLB[158] WLB[157] WLB[156] WLB[155] WLB[154]
+WLB[153] WLB[152] WLB[151] WLB[150] WLB[149] WLB[148] WLB[147] WLB[146] WLB[145] WLB[144]
+WLB[143] WLB[142] WLB[141] WLB[140] WLB[139] WLB[138] WLB[137] WLB[136] WLB[135] WLB[134]
+WLB[133] WLB[132] WLB[131] WLB[130] WLB[129] WLB[128] WLB[127] WLB[126] WLB[125] WLB[124]
+WLB[123] WLB[122] WLB[121] WLB[120] WLB[119] WLB[118] WLB[117] WLB[116] WLB[115] WLB[114]
+WLB[113] WLB[112] WLB[111] WLB[110] WLB[109] WLB[108] WLB[107] WLB[106] WLB[105] WLB[104]
+WLB[103] WLB[102] WLB[101] WLB[100] WLB[99] WLB[98] WLB[97] WLB[96] WLB[95] WLB[94]
+WLB[93] WLB[92] WLB[91] WLB[90] WLB[89] WLB[88] WLB[87] WLB[86] WLB[85] WLB[84]
+WLB[83] WLB[82] WLB[81] WLB[80] WLB[79] WLB[78] WLB[77] WLB[76] WLB[75] WLB[74]
+WLB[73] WLB[72] WLB[71] WLB[70] WLB[69] WLB[68] WLB[67] WLB[66] WLB[65] WLB[64]
+WLB[63] WLB[62] WLB[61] WLB[60] WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54]
+WLB[53] WLB[52] WLB[51] WLB[50] WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44]
+WLB[43] WLB[42] WLB[41] WLB[40] WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34]
+WLB[33] WLB[32] WLB[31] WLB[30] WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24]
+WLB[23] WLB[22] WLB[21] WLB[20] WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14]
+WLB[13] WLB[12] WLB[11] WLB[10] WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4]
+WLB[3] WLB[2] WLB[1] WLB[0] S55NLLGDPH_X512Y8D16_BW_XDEC64
XI6 AB[10] AB[11] ACTRCLKB ACTRCLKXB PXCB[3] PXCB[2] PXCB[1] PXCB[0] VDD VSS S55NLLGDPH_X512Y8D16_BW_PX4
XI7 AA[10] AA[11] ACTRCLKA ACTRCLKXA PXCA[3] PXCA[2] PXCA[1] PXCA[0] VDD VSS S55NLLGDPH_X512Y8D16_BW_PX4
XI8 AB[8] AB[9] ACTRCLKB ACTRCLKXB PXBB[3] PXBB[2] PXBB[1] PXBB[0] VDD VSS S55NLLGDPH_X512Y8D16_BW_PX4
XI9 AA[8] AA[9] ACTRCLKA ACTRCLKXA PXBA[3] PXBA[2] PXBA[1] PXBA[0] VDD VSS S55NLLGDPH_X512Y8D16_BW_PX4
XI10 AA[7] AA[6] AA[5] AA[4] AA[3] AA[2] AA[1] AA[0] ACTRCLKA ACTRCLKXA
+CENA CLKA DCTRCLKA DCTRCLKXA EMCLKA DBLA FCKXA[7] FCKXA[6] FCKXA[5] FCKXA[4]
+FCKXA[3] FCKXA[2] FCKXA[1] FCKXA[0] PXAA[3] PXAA[2] PXAA[1] PXAA[0] RDE RWLA
+TIE_LOW TIE_LOW SACK1A SACK4A VDD VSS WEA WENA YXA[7] YXA[6]
+YXA[5] YXA[4] YXA[3] YXA[2] YXA[1] YXA[0] S55NLLGDPH_X512Y8D16_BW_LOGIC_BASE_Y8
XI11 AB[7] AB[6] AB[5] AB[4] AB[3] AB[2] AB[1] AB[0] ACTRCLKB ACTRCLKXB
+CENB CLKB DCTRCLKB DCTRCLKXB EMCLKB DBLB FCKXB[7] FCKXB[6] FCKXB[5] FCKXB[4]
+FCKXB[3] FCKXB[2] FCKXB[1] FCKXB[0] PXAB[3] PXAB[2] PXAB[1] PXAB[0] RDE RWLB
+TIE_LOW TIE_LOW SACK1B SACK4B VDD VSS WEB WENB YXB[7] YXB[6]
+YXB[5] YXB[4] YXB[3] YXB[2] YXB[1] YXB[0] S55NLLGDPH_X512Y8D16_BW_LOGIC_BASE_Y8
XI12 AA[11] AA[10] AA[9] AA[8] AA[7] AA[6] AA[5] AA[4] AA[3] AA[2]
+AA[1] AA[0] CENA CLKA WENA VDD VSS S55NLLGDPH_X512Y8D16_BW_ESDA11
XI13 AB[11] AB[10] AB[9] AB[8] AB[7] AB[6] AB[5] AB[4] AB[3] AB[2]
+AB[1] AB[0] CENB CLKB WENB VDD VSS S55NLLGDPH_X512Y8D16_BW_ESDA11
XI14 TIE_LOW VSS VDD S55NLLGDPH_X512Y8D16_BW_TIE_LOW_S
XI15 TIE_HIGH VSS VDD S55NLLGDPH_X512Y8D16_BW_TIE_HIGH_S
XI16 TIE_LOW TIE_LOW SOPB[2] SOPB[1] SOPB[0] VDD VSS S55NLLGDPH_X512Y8D16_BW_OPDEC
XI17 TIE_LOW TIE_LOW SOPA[2] SOPA[1] SOPA[0] VDD VSS S55NLLGDPH_X512Y8D16_BW_OPDEC
XI18 RDE VSS VDD S55NLLGDPH_X512Y8D16_BW_TIE_LOW_X2
XI19 DBLB STWLB SOPB[2] SOPB[1] SOPB[0] VDD VSS S55NLLGDPH_X512Y8D16_BW_DISCHARGECELLS
XI20 DBLA STWLA SOPA[2] SOPA[1] SOPA[0] VDD VSS S55NLLGDPH_X512Y8D16_BW_DISCHARGECELLS
.ENDS
