// removed module with interface ports: DcpSwitchUnit
