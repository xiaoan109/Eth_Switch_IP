// removed module with interface ports: DcpRouteUnit
