// removed module with interface ports: RdCtrlTop16Ch
