// removed module with interface ports: RdDstLock
