// removed module with interface ports: DcpRdCmd16x16
