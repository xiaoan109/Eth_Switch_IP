// removed module with interface ports: PortCtrl
