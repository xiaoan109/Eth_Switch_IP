module RdScheTopWrapper (
	iClk,
	iRst_n,
	oPkgRdy0,
	iPkgPri0,
	iPkgDstPort0,
	iPkgFirAddr0,
	iPkgLen0,
	iPkgTagVld0,
	oPkgRdy1,
	iPkgPri1,
	iPkgDstPort1,
	iPkgFirAddr1,
	iPkgLen1,
	iPkgTagVld1,
	oPkgRdy2,
	iPkgPri2,
	iPkgDstPort2,
	iPkgFirAddr2,
	iPkgLen2,
	iPkgTagVld2,
	oPkgRdy3,
	iPkgPri3,
	iPkgDstPort3,
	iPkgFirAddr3,
	iPkgLen3,
	iPkgTagVld3,
	oPkgRdy4,
	iPkgPri4,
	iPkgDstPort4,
	iPkgFirAddr4,
	iPkgLen4,
	iPkgTagVld4,
	oPkgRdy5,
	iPkgPri5,
	iPkgDstPort5,
	iPkgFirAddr5,
	iPkgLen5,
	iPkgTagVld5,
	oPkgRdy6,
	iPkgPri6,
	iPkgDstPort6,
	iPkgFirAddr6,
	iPkgLen6,
	iPkgTagVld6,
	oPkgRdy7,
	iPkgPri7,
	iPkgDstPort7,
	iPkgFirAddr7,
	iPkgLen7,
	iPkgTagVld7,
	oPkgRdy8,
	iPkgPri8,
	iPkgDstPort8,
	iPkgFirAddr8,
	iPkgLen8,
	iPkgTagVld8,
	oPkgRdy9,
	iPkgPri9,
	iPkgDstPort9,
	iPkgFirAddr9,
	iPkgLen9,
	iPkgTagVld9,
	oPkgRdy10,
	iPkgPri10,
	iPkgDstPort10,
	iPkgFirAddr10,
	iPkgLen10,
	iPkgTagVld10,
	oPkgRdy11,
	iPkgPri11,
	iPkgDstPort11,
	iPkgFirAddr11,
	iPkgLen11,
	iPkgTagVld11,
	oPkgRdy12,
	iPkgPri12,
	iPkgDstPort12,
	iPkgFirAddr12,
	iPkgLen12,
	iPkgTagVld12,
	oPkgRdy13,
	iPkgPri13,
	iPkgDstPort13,
	iPkgFirAddr13,
	iPkgLen13,
	iPkgTagVld13,
	oPkgRdy14,
	iPkgPri14,
	iPkgDstPort14,
	iPkgFirAddr14,
	iPkgLen14,
	iPkgTagVld14,
	oPkgRdy15,
	iPkgPri15,
	iPkgDstPort15,
	iPkgFirAddr15,
	iPkgLen15,
	iPkgTagVld15,
	oPkgFirAddr0,
	oPkgFirAddrVld0,
	oPkgBlockNum0,
	oPkgDrop0,
	iPkgFirAddrRdy0,
	oPkgFirAddr1,
	oPkgFirAddrVld1,
	oPkgBlockNum1,
	oPkgDrop1,
	iPkgFirAddrRdy1,
	oPkgFirAddr2,
	oPkgFirAddrVld2,
	oPkgBlockNum2,
	oPkgDrop2,
	iPkgFirAddrRdy2,
	oPkgFirAddr3,
	oPkgFirAddrVld3,
	oPkgBlockNum3,
	oPkgDrop3,
	iPkgFirAddrRdy3,
	oPkgFirAddr4,
	oPkgFirAddrVld4,
	oPkgBlockNum4,
	oPkgDrop4,
	iPkgFirAddrRdy4,
	oPkgFirAddr5,
	oPkgFirAddrVld5,
	oPkgBlockNum5,
	oPkgDrop5,
	iPkgFirAddrRdy5,
	oPkgFirAddr6,
	oPkgFirAddrVld6,
	oPkgBlockNum6,
	oPkgDrop6,
	iPkgFirAddrRdy6,
	oPkgFirAddr7,
	oPkgFirAddrVld7,
	oPkgBlockNum7,
	oPkgDrop7,
	iPkgFirAddrRdy7,
	oPkgFirAddr8,
	oPkgFirAddrVld8,
	oPkgBlockNum8,
	oPkgDrop8,
	iPkgFirAddrRdy8,
	oPkgFirAddr9,
	oPkgFirAddrVld9,
	oPkgBlockNum9,
	oPkgDrop9,
	iPkgFirAddrRdy9,
	oPkgFirAddr10,
	oPkgFirAddrVld10,
	oPkgBlockNum10,
	oPkgDrop10,
	iPkgFirAddrRdy10,
	oPkgFirAddr11,
	oPkgFirAddrVld11,
	oPkgBlockNum11,
	oPkgDrop11,
	iPkgFirAddrRdy11,
	oPkgFirAddr12,
	oPkgFirAddrVld12,
	oPkgBlockNum12,
	oPkgDrop12,
	iPkgFirAddrRdy12,
	oPkgFirAddr13,
	oPkgFirAddrVld13,
	oPkgBlockNum13,
	oPkgDrop13,
	iPkgFirAddrRdy13,
	oPkgFirAddr14,
	oPkgFirAddrVld14,
	oPkgBlockNum14,
	oPkgDrop14,
	iPkgFirAddrRdy14,
	oPkgFirAddr15,
	oPkgFirAddrVld15,
	oPkgBlockNum15,
	oPkgDrop15,
	iPkgFirAddrRdy15,
	iWrrData0,
	iWrrVld0,
	iWrrLast0,
	oWrrRdy0,
	iWrrData1,
	iWrrVld1,
	iWrrLast1,
	oWrrRdy1,
	iWrrData2,
	iWrrVld2,
	iWrrLast2,
	oWrrRdy2,
	iWrrData3,
	iWrrVld3,
	iWrrLast3,
	oWrrRdy3,
	iWrrData4,
	iWrrVld4,
	iWrrLast4,
	oWrrRdy4,
	iWrrData5,
	iWrrVld5,
	iWrrLast5,
	oWrrRdy5,
	iWrrData6,
	iWrrVld6,
	iWrrLast6,
	oWrrRdy6,
	iWrrData7,
	iWrrVld7,
	iWrrLast7,
	oWrrRdy7,
	iWrrData8,
	iWrrVld8,
	iWrrLast8,
	oWrrRdy8,
	iWrrData9,
	iWrrVld9,
	iWrrLast9,
	oWrrRdy9,
	iWrrData10,
	iWrrVld10,
	iWrrLast10,
	oWrrRdy10,
	iWrrData11,
	iWrrVld11,
	iWrrLast11,
	oWrrRdy11,
	iWrrData12,
	iWrrVld12,
	iWrrLast12,
	oWrrRdy12,
	iWrrData13,
	iWrrVld13,
	iWrrLast13,
	oWrrRdy13,
	iWrrData14,
	iWrrVld14,
	iWrrLast14,
	oWrrRdy14,
	iWrrData15,
	iWrrVld15,
	iWrrLast15,
	oWrrRdy15,
	oRdSop0,
	oRdEop0,
	oRdVld0,
	oRdData0,
	iRdRdy0,
	oRdLast0,
	oRdSop1,
	oRdEop1,
	oRdVld1,
	oRdData1,
	iRdRdy1,
	oRdLast1,
	oRdSop2,
	oRdEop2,
	oRdVld2,
	oRdData2,
	iRdRdy2,
	oRdLast2,
	oRdSop3,
	oRdEop3,
	oRdVld3,
	oRdData3,
	iRdRdy3,
	oRdLast3,
	oRdSop4,
	oRdEop4,
	oRdVld4,
	oRdData4,
	iRdRdy4,
	oRdLast4,
	oRdSop5,
	oRdEop5,
	oRdVld5,
	oRdData5,
	iRdRdy5,
	oRdLast5,
	oRdSop6,
	oRdEop6,
	oRdVld6,
	oRdData6,
	iRdRdy6,
	oRdLast6,
	oRdSop7,
	oRdEop7,
	oRdVld7,
	oRdData7,
	iRdRdy7,
	oRdLast7,
	oRdSop8,
	oRdEop8,
	oRdVld8,
	oRdData8,
	iRdRdy8,
	oRdLast8,
	oRdSop9,
	oRdEop9,
	oRdVld9,
	oRdData9,
	iRdRdy9,
	oRdLast9,
	oRdSop10,
	oRdEop10,
	oRdVld10,
	oRdData10,
	iRdRdy10,
	oRdLast10,
	oRdSop11,
	oRdEop11,
	oRdVld11,
	oRdData11,
	iRdRdy11,
	oRdLast11,
	oRdSop12,
	oRdEop12,
	oRdVld12,
	oRdData12,
	iRdRdy12,
	oRdLast12,
	oRdSop13,
	oRdEop13,
	oRdVld13,
	oRdData13,
	iRdRdy13,
	oRdLast13,
	oRdSop14,
	oRdEop14,
	oRdVld14,
	oRdData14,
	iRdRdy14,
	oRdLast14,
	oRdSop15,
	oRdEop15,
	oRdVld15,
	oRdData15,
	iRdRdy15,
	oRdLast15,
	iWrrWeightPld0,
	iWrrWeightPld1,
	iWrrWeightPld2,
	iWrrWeightPld3,
	iWrrWeightPld4,
	iWrrWeightPld5,
	iWrrWeightPld6,
	iWrrWeightPld7,
	iWrrWeightIdx,
	iWrrWeightLoad
);
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:3:13
	parameter PRI_DEPTH = 8;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:4:13
	parameter WRR_WEIGHT_NUM = 8;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:6:3
	input wire iClk;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:7:3
	input wire iRst_n;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:10:3
	output wire oPkgRdy0;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:11:3
	input wire [2:0] iPkgPri0;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:12:3
	input wire [3:0] iPkgDstPort0;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:13:3
	input wire [11:0] iPkgFirAddr0;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:14:3
	input wire [3:0] iPkgLen0;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:15:3
	input wire iPkgTagVld0;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:17:3
	output wire oPkgRdy1;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:18:3
	input wire [2:0] iPkgPri1;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:19:3
	input wire [3:0] iPkgDstPort1;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:20:3
	input wire [11:0] iPkgFirAddr1;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:21:3
	input wire [3:0] iPkgLen1;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:22:3
	input wire iPkgTagVld1;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:24:3
	output wire oPkgRdy2;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:25:3
	input wire [2:0] iPkgPri2;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:26:3
	input wire [3:0] iPkgDstPort2;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:27:3
	input wire [11:0] iPkgFirAddr2;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:28:3
	input wire [3:0] iPkgLen2;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:29:3
	input wire iPkgTagVld2;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:31:3
	output wire oPkgRdy3;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:32:3
	input wire [2:0] iPkgPri3;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:33:3
	input wire [3:0] iPkgDstPort3;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:34:3
	input wire [11:0] iPkgFirAddr3;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:35:3
	input wire [3:0] iPkgLen3;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:36:3
	input wire iPkgTagVld3;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:38:3
	output wire oPkgRdy4;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:39:3
	input wire [2:0] iPkgPri4;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:40:3
	input wire [3:0] iPkgDstPort4;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:41:3
	input wire [11:0] iPkgFirAddr4;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:42:3
	input wire [3:0] iPkgLen4;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:43:3
	input wire iPkgTagVld4;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:45:3
	output wire oPkgRdy5;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:46:3
	input wire [2:0] iPkgPri5;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:47:3
	input wire [3:0] iPkgDstPort5;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:48:3
	input wire [11:0] iPkgFirAddr5;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:49:3
	input wire [3:0] iPkgLen5;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:50:3
	input wire iPkgTagVld5;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:52:3
	output wire oPkgRdy6;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:53:3
	input wire [2:0] iPkgPri6;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:54:3
	input wire [3:0] iPkgDstPort6;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:55:3
	input wire [11:0] iPkgFirAddr6;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:56:3
	input wire [3:0] iPkgLen6;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:57:3
	input wire iPkgTagVld6;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:59:3
	output wire oPkgRdy7;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:60:3
	input wire [2:0] iPkgPri7;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:61:3
	input wire [3:0] iPkgDstPort7;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:62:3
	input wire [11:0] iPkgFirAddr7;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:63:3
	input wire [3:0] iPkgLen7;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:64:3
	input wire iPkgTagVld7;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:66:3
	output wire oPkgRdy8;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:67:3
	input wire [2:0] iPkgPri8;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:68:3
	input wire [3:0] iPkgDstPort8;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:69:3
	input wire [11:0] iPkgFirAddr8;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:70:3
	input wire [3:0] iPkgLen8;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:71:3
	input wire iPkgTagVld8;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:73:3
	output wire oPkgRdy9;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:74:3
	input wire [2:0] iPkgPri9;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:75:3
	input wire [3:0] iPkgDstPort9;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:76:3
	input wire [11:0] iPkgFirAddr9;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:77:3
	input wire [3:0] iPkgLen9;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:78:3
	input wire iPkgTagVld9;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:80:3
	output wire oPkgRdy10;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:81:3
	input wire [2:0] iPkgPri10;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:82:3
	input wire [3:0] iPkgDstPort10;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:83:3
	input wire [11:0] iPkgFirAddr10;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:84:3
	input wire [3:0] iPkgLen10;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:85:3
	input wire iPkgTagVld10;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:87:3
	output wire oPkgRdy11;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:88:3
	input wire [2:0] iPkgPri11;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:89:3
	input wire [3:0] iPkgDstPort11;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:90:3
	input wire [11:0] iPkgFirAddr11;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:91:3
	input wire [3:0] iPkgLen11;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:92:3
	input wire iPkgTagVld11;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:94:3
	output wire oPkgRdy12;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:95:3
	input wire [2:0] iPkgPri12;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:96:3
	input wire [3:0] iPkgDstPort12;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:97:3
	input wire [11:0] iPkgFirAddr12;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:98:3
	input wire [3:0] iPkgLen12;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:99:3
	input wire iPkgTagVld12;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:101:3
	output wire oPkgRdy13;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:102:3
	input wire [2:0] iPkgPri13;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:103:3
	input wire [3:0] iPkgDstPort13;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:104:3
	input wire [11:0] iPkgFirAddr13;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:105:3
	input wire [3:0] iPkgLen13;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:106:3
	input wire iPkgTagVld13;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:108:3
	output wire oPkgRdy14;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:109:3
	input wire [2:0] iPkgPri14;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:110:3
	input wire [3:0] iPkgDstPort14;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:111:3
	input wire [11:0] iPkgFirAddr14;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:112:3
	input wire [3:0] iPkgLen14;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:113:3
	input wire iPkgTagVld14;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:115:3
	output wire oPkgRdy15;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:116:3
	input wire [2:0] iPkgPri15;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:117:3
	input wire [3:0] iPkgDstPort15;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:118:3
	input wire [11:0] iPkgFirAddr15;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:119:3
	input wire [3:0] iPkgLen15;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:120:3
	input wire iPkgTagVld15;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:123:3
	output wire [11:0] oPkgFirAddr0;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:124:3
	output wire oPkgFirAddrVld0;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:125:3
	output wire [3:0] oPkgBlockNum0;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:126:3
	output wire oPkgDrop0;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:127:3
	input wire iPkgFirAddrRdy0;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:129:3
	output wire [11:0] oPkgFirAddr1;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:130:3
	output wire oPkgFirAddrVld1;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:131:3
	output wire [3:0] oPkgBlockNum1;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:132:3
	output wire oPkgDrop1;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:133:3
	input wire iPkgFirAddrRdy1;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:135:3
	output wire [11:0] oPkgFirAddr2;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:136:3
	output wire oPkgFirAddrVld2;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:137:3
	output wire [3:0] oPkgBlockNum2;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:138:3
	output wire oPkgDrop2;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:139:3
	input wire iPkgFirAddrRdy2;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:141:3
	output wire [11:0] oPkgFirAddr3;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:142:3
	output wire oPkgFirAddrVld3;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:143:3
	output wire [3:0] oPkgBlockNum3;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:144:3
	output wire oPkgDrop3;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:145:3
	input wire iPkgFirAddrRdy3;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:147:3
	output wire [11:0] oPkgFirAddr4;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:148:3
	output wire oPkgFirAddrVld4;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:149:3
	output wire [3:0] oPkgBlockNum4;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:150:3
	output wire oPkgDrop4;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:151:3
	input wire iPkgFirAddrRdy4;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:153:3
	output wire [11:0] oPkgFirAddr5;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:154:3
	output wire oPkgFirAddrVld5;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:155:3
	output wire [3:0] oPkgBlockNum5;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:156:3
	output wire oPkgDrop5;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:157:3
	input wire iPkgFirAddrRdy5;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:159:3
	output wire [11:0] oPkgFirAddr6;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:160:3
	output wire oPkgFirAddrVld6;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:161:3
	output wire [3:0] oPkgBlockNum6;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:162:3
	output wire oPkgDrop6;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:163:3
	input wire iPkgFirAddrRdy6;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:165:3
	output wire [11:0] oPkgFirAddr7;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:166:3
	output wire oPkgFirAddrVld7;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:167:3
	output wire [3:0] oPkgBlockNum7;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:168:3
	output wire oPkgDrop7;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:169:3
	input wire iPkgFirAddrRdy7;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:171:3
	output wire [11:0] oPkgFirAddr8;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:172:3
	output wire oPkgFirAddrVld8;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:173:3
	output wire [3:0] oPkgBlockNum8;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:174:3
	output wire oPkgDrop8;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:175:3
	input wire iPkgFirAddrRdy8;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:177:3
	output wire [11:0] oPkgFirAddr9;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:178:3
	output wire oPkgFirAddrVld9;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:179:3
	output wire [3:0] oPkgBlockNum9;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:180:3
	output wire oPkgDrop9;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:181:3
	input wire iPkgFirAddrRdy9;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:183:3
	output wire [11:0] oPkgFirAddr10;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:184:3
	output wire oPkgFirAddrVld10;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:185:3
	output wire [3:0] oPkgBlockNum10;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:186:3
	output wire oPkgDrop10;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:187:3
	input wire iPkgFirAddrRdy10;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:189:3
	output wire [11:0] oPkgFirAddr11;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:190:3
	output wire oPkgFirAddrVld11;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:191:3
	output wire [3:0] oPkgBlockNum11;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:192:3
	output wire oPkgDrop11;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:193:3
	input wire iPkgFirAddrRdy11;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:195:3
	output wire [11:0] oPkgFirAddr12;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:196:3
	output wire oPkgFirAddrVld12;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:197:3
	output wire [3:0] oPkgBlockNum12;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:198:3
	output wire oPkgDrop12;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:199:3
	input wire iPkgFirAddrRdy12;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:201:3
	output wire [11:0] oPkgFirAddr13;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:202:3
	output wire oPkgFirAddrVld13;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:203:3
	output wire [3:0] oPkgBlockNum13;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:204:3
	output wire oPkgDrop13;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:205:3
	input wire iPkgFirAddrRdy13;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:207:3
	output wire [11:0] oPkgFirAddr14;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:208:3
	output wire oPkgFirAddrVld14;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:209:3
	output wire [3:0] oPkgBlockNum14;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:210:3
	output wire oPkgDrop14;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:211:3
	input wire iPkgFirAddrRdy14;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:213:3
	output wire [11:0] oPkgFirAddr15;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:214:3
	output wire oPkgFirAddrVld15;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:215:3
	output wire [3:0] oPkgBlockNum15;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:216:3
	output wire oPkgDrop15;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:217:3
	input wire iPkgFirAddrRdy15;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:220:3
	input wire [31:0] iWrrData0;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:221:3
	input wire iWrrVld0;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:222:3
	input wire iWrrLast0;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:223:3
	output wire oWrrRdy0;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:225:3
	input wire [31:0] iWrrData1;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:226:3
	input wire iWrrVld1;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:227:3
	input wire iWrrLast1;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:228:3
	output wire oWrrRdy1;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:230:3
	input wire [31:0] iWrrData2;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:231:3
	input wire iWrrVld2;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:232:3
	input wire iWrrLast2;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:233:3
	output wire oWrrRdy2;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:235:3
	input wire [31:0] iWrrData3;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:236:3
	input wire iWrrVld3;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:237:3
	input wire iWrrLast3;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:238:3
	output wire oWrrRdy3;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:240:3
	input wire [31:0] iWrrData4;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:241:3
	input wire iWrrVld4;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:242:3
	input wire iWrrLast4;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:243:3
	output wire oWrrRdy4;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:245:3
	input wire [31:0] iWrrData5;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:246:3
	input wire iWrrVld5;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:247:3
	input wire iWrrLast5;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:248:3
	output wire oWrrRdy5;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:250:3
	input wire [31:0] iWrrData6;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:251:3
	input wire iWrrVld6;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:252:3
	input wire iWrrLast6;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:253:3
	output wire oWrrRdy6;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:255:3
	input wire [31:0] iWrrData7;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:256:3
	input wire iWrrVld7;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:257:3
	input wire iWrrLast7;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:258:3
	output wire oWrrRdy7;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:260:3
	input wire [31:0] iWrrData8;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:261:3
	input wire iWrrVld8;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:262:3
	input wire iWrrLast8;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:263:3
	output wire oWrrRdy8;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:265:3
	input wire [31:0] iWrrData9;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:266:3
	input wire iWrrVld9;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:267:3
	input wire iWrrLast9;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:268:3
	output wire oWrrRdy9;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:270:3
	input wire [31:0] iWrrData10;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:271:3
	input wire iWrrVld10;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:272:3
	input wire iWrrLast10;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:273:3
	output wire oWrrRdy10;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:275:3
	input wire [31:0] iWrrData11;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:276:3
	input wire iWrrVld11;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:277:3
	input wire iWrrLast11;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:278:3
	output wire oWrrRdy11;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:280:3
	input wire [31:0] iWrrData12;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:281:3
	input wire iWrrVld12;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:282:3
	input wire iWrrLast12;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:283:3
	output wire oWrrRdy12;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:285:3
	input wire [31:0] iWrrData13;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:286:3
	input wire iWrrVld13;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:287:3
	input wire iWrrLast13;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:288:3
	output wire oWrrRdy13;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:290:3
	input wire [31:0] iWrrData14;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:291:3
	input wire iWrrVld14;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:292:3
	input wire iWrrLast14;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:293:3
	output wire oWrrRdy14;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:295:3
	input wire [31:0] iWrrData15;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:296:3
	input wire iWrrVld15;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:297:3
	input wire iWrrLast15;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:298:3
	output wire oWrrRdy15;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:301:3
	output wire oRdSop0;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:302:3
	output wire oRdEop0;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:303:3
	output wire oRdVld0;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:304:3
	output wire [31:0] oRdData0;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:305:3
	input wire iRdRdy0;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:306:3
	output wire oRdLast0;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:308:3
	output wire oRdSop1;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:309:3
	output wire oRdEop1;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:310:3
	output wire oRdVld1;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:311:3
	output wire [31:0] oRdData1;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:312:3
	input wire iRdRdy1;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:313:3
	output wire oRdLast1;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:315:3
	output wire oRdSop2;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:316:3
	output wire oRdEop2;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:317:3
	output wire oRdVld2;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:318:3
	output wire [31:0] oRdData2;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:319:3
	input wire iRdRdy2;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:320:3
	output wire oRdLast2;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:322:3
	output wire oRdSop3;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:323:3
	output wire oRdEop3;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:324:3
	output wire oRdVld3;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:325:3
	output wire [31:0] oRdData3;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:326:3
	input wire iRdRdy3;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:327:3
	output wire oRdLast3;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:329:3
	output wire oRdSop4;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:330:3
	output wire oRdEop4;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:331:3
	output wire oRdVld4;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:332:3
	output wire [31:0] oRdData4;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:333:3
	input wire iRdRdy4;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:334:3
	output wire oRdLast4;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:336:3
	output wire oRdSop5;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:337:3
	output wire oRdEop5;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:338:3
	output wire oRdVld5;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:339:3
	output wire [31:0] oRdData5;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:340:3
	input wire iRdRdy5;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:341:3
	output wire oRdLast5;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:343:3
	output wire oRdSop6;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:344:3
	output wire oRdEop6;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:345:3
	output wire oRdVld6;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:346:3
	output wire [31:0] oRdData6;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:347:3
	input wire iRdRdy6;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:348:3
	output wire oRdLast6;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:350:3
	output wire oRdSop7;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:351:3
	output wire oRdEop7;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:352:3
	output wire oRdVld7;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:353:3
	output wire [31:0] oRdData7;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:354:3
	input wire iRdRdy7;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:355:3
	output wire oRdLast7;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:357:3
	output wire oRdSop8;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:358:3
	output wire oRdEop8;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:359:3
	output wire oRdVld8;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:360:3
	output wire [31:0] oRdData8;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:361:3
	input wire iRdRdy8;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:362:3
	output wire oRdLast8;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:364:3
	output wire oRdSop9;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:365:3
	output wire oRdEop9;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:366:3
	output wire oRdVld9;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:367:3
	output wire [31:0] oRdData9;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:368:3
	input wire iRdRdy9;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:369:3
	output wire oRdLast9;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:371:3
	output wire oRdSop10;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:372:3
	output wire oRdEop10;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:373:3
	output wire oRdVld10;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:374:3
	output wire [31:0] oRdData10;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:375:3
	input wire iRdRdy10;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:376:3
	output wire oRdLast10;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:378:3
	output wire oRdSop11;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:379:3
	output wire oRdEop11;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:380:3
	output wire oRdVld11;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:381:3
	output wire [31:0] oRdData11;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:382:3
	input wire iRdRdy11;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:383:3
	output wire oRdLast11;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:385:3
	output wire oRdSop12;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:386:3
	output wire oRdEop12;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:387:3
	output wire oRdVld12;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:388:3
	output wire [31:0] oRdData12;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:389:3
	input wire iRdRdy12;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:390:3
	output wire oRdLast12;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:392:3
	output wire oRdSop13;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:393:3
	output wire oRdEop13;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:394:3
	output wire oRdVld13;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:395:3
	output wire [31:0] oRdData13;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:396:3
	input wire iRdRdy13;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:397:3
	output wire oRdLast13;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:399:3
	output wire oRdSop14;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:400:3
	output wire oRdEop14;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:401:3
	output wire oRdVld14;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:402:3
	output wire [31:0] oRdData14;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:403:3
	input wire iRdRdy14;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:404:3
	output wire oRdLast14;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:406:3
	output wire oRdSop15;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:407:3
	output wire oRdEop15;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:408:3
	output wire oRdVld15;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:409:3
	output wire [31:0] oRdData15;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:410:3
	input wire iRdRdy15;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:411:3
	output wire oRdLast15;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:414:3
	input wire [$clog2(WRR_WEIGHT_NUM):0] iWrrWeightPld0;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:415:3
	input wire [$clog2(WRR_WEIGHT_NUM):0] iWrrWeightPld1;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:416:3
	input wire [$clog2(WRR_WEIGHT_NUM):0] iWrrWeightPld2;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:417:3
	input wire [$clog2(WRR_WEIGHT_NUM):0] iWrrWeightPld3;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:418:3
	input wire [$clog2(WRR_WEIGHT_NUM):0] iWrrWeightPld4;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:419:3
	input wire [$clog2(WRR_WEIGHT_NUM):0] iWrrWeightPld5;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:420:3
	input wire [$clog2(WRR_WEIGHT_NUM):0] iWrrWeightPld6;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:421:3
	input wire [$clog2(WRR_WEIGHT_NUM):0] iWrrWeightPld7;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:422:3
	input wire [3:0] iWrrWeightIdx;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:423:3
	input wire iWrrWeightLoad;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:426:3
	localparam TAG_WIDTH = 23;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:427:3
	localparam RDCMD_WIDTH = 21;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:428:3
	localparam RDDATA_WIDTH = 33;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:431:3
	// expanded interface instance: intTag
	localparam _param_83F1A_DW = TAG_WIDTH;
	localparam _param_83F1A_AW = 4;
	genvar _arr_83F1A;
	generate
		for (_arr_83F1A = 0; _arr_83F1A <= 15; _arr_83F1A = _arr_83F1A + 1) begin : intTag
			// Trace: src/src/rtl/design/svsrc/interface_list.sv:64:33
			localparam DW = _param_83F1A_DW;
			// Trace: src/src/rtl/design/svsrc/interface_list.sv:64:52
			localparam AW = _param_83F1A_AW;
			// Trace: src/src/rtl/design/svsrc/interface_list.sv:65:3
			wire [22:0] Pld;
			// Trace: src/src/rtl/design/svsrc/interface_list.sv:66:3
			wire [3:0] Dst;
			// Trace: src/src/rtl/design/svsrc/interface_list.sv:67:3
			wire Vld;
			// Trace: src/src/rtl/design/svsrc/interface_list.sv:68:3
			wire Rdy;
			// Trace: src/src/rtl/design/svsrc/interface_list.sv:69:3
			// Trace: src/src/rtl/design/svsrc/interface_list.sv:75:3
		end
	endgenerate
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:432:3
	// expanded interface instance: intRdCmd
	localparam _param_F36BA_DW = RDCMD_WIDTH;
	localparam _param_F36BA_AW = 4;
	genvar _arr_F36BA;
	generate
		for (_arr_F36BA = 0; _arr_F36BA <= 15; _arr_F36BA = _arr_F36BA + 1) begin : intRdCmd
			// Trace: src/src/rtl/design/svsrc/interface_list.sv:64:33
			localparam DW = _param_F36BA_DW;
			// Trace: src/src/rtl/design/svsrc/interface_list.sv:64:52
			localparam AW = _param_F36BA_AW;
			// Trace: src/src/rtl/design/svsrc/interface_list.sv:65:3
			wire [20:0] Pld;
			// Trace: src/src/rtl/design/svsrc/interface_list.sv:66:3
			wire [3:0] Dst;
			// Trace: src/src/rtl/design/svsrc/interface_list.sv:67:3
			wire Vld;
			// Trace: src/src/rtl/design/svsrc/interface_list.sv:68:3
			wire Rdy;
			// Trace: src/src/rtl/design/svsrc/interface_list.sv:69:3
			// Trace: src/src/rtl/design/svsrc/interface_list.sv:75:3
		end
	endgenerate
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:433:3
	// expanded interface instance: intRdData
	localparam _param_8CEC1_DW = RDDATA_WIDTH;
	localparam _param_8CEC1_AW = 4;
	genvar _arr_8CEC1;
	generate
		for (_arr_8CEC1 = 0; _arr_8CEC1 <= 15; _arr_8CEC1 = _arr_8CEC1 + 1) begin : intRdData
			// Trace: src/src/rtl/design/svsrc/interface_list.sv:64:33
			localparam DW = _param_8CEC1_DW;
			// Trace: src/src/rtl/design/svsrc/interface_list.sv:64:52
			localparam AW = _param_8CEC1_AW;
			// Trace: src/src/rtl/design/svsrc/interface_list.sv:65:3
			wire [32:0] Pld;
			// Trace: src/src/rtl/design/svsrc/interface_list.sv:66:3
			wire [3:0] Dst;
			// Trace: src/src/rtl/design/svsrc/interface_list.sv:67:3
			wire Vld;
			// Trace: src/src/rtl/design/svsrc/interface_list.sv:68:3
			wire Rdy;
			// Trace: src/src/rtl/design/svsrc/interface_list.sv:69:3
			// Trace: src/src/rtl/design/svsrc/interface_list.sv:75:3
		end
	endgenerate
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:436:3
	assign intTag[0].Vld = iPkgTagVld0;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:437:3
	assign intTag[0].Dst = iPkgDstPort0;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:438:3
	assign intTag[0].Pld = {iPkgPri0, iPkgFirAddr0, iPkgLen0, 4'h0};
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:439:3
	assign oPkgRdy0 = intTag[0].Rdy;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:441:3
	assign intTag[1].Vld = iPkgTagVld1;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:442:3
	assign intTag[1].Dst = iPkgDstPort1;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:443:3
	assign intTag[1].Pld = {iPkgPri1, iPkgFirAddr1, iPkgLen1, 4'h1};
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:444:3
	assign oPkgRdy1 = intTag[1].Rdy;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:446:3
	assign intTag[2].Vld = iPkgTagVld2;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:447:3
	assign intTag[2].Dst = iPkgDstPort2;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:448:3
	assign intTag[2].Pld = {iPkgPri2, iPkgFirAddr2, iPkgLen2, 4'h2};
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:449:3
	assign oPkgRdy2 = intTag[2].Rdy;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:451:3
	assign intTag[3].Vld = iPkgTagVld3;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:452:3
	assign intTag[3].Dst = iPkgDstPort3;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:453:3
	assign intTag[3].Pld = {iPkgPri3, iPkgFirAddr3, iPkgLen3, 4'h3};
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:454:3
	assign oPkgRdy3 = intTag[3].Rdy;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:456:3
	assign intTag[4].Vld = iPkgTagVld4;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:457:3
	assign intTag[4].Dst = iPkgDstPort4;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:458:3
	assign intTag[4].Pld = {iPkgPri4, iPkgFirAddr4, iPkgLen4, 4'h4};
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:459:3
	assign oPkgRdy4 = intTag[4].Rdy;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:461:3
	assign intTag[5].Vld = iPkgTagVld5;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:462:3
	assign intTag[5].Dst = iPkgDstPort5;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:463:3
	assign intTag[5].Pld = {iPkgPri5, iPkgFirAddr5, iPkgLen5, 4'h5};
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:464:3
	assign oPkgRdy5 = intTag[5].Rdy;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:466:3
	assign intTag[6].Vld = iPkgTagVld6;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:467:3
	assign intTag[6].Dst = iPkgDstPort6;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:468:3
	assign intTag[6].Pld = {iPkgPri6, iPkgFirAddr6, iPkgLen6, 4'h6};
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:469:3
	assign oPkgRdy6 = intTag[6].Rdy;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:471:3
	assign intTag[7].Vld = iPkgTagVld7;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:472:3
	assign intTag[7].Dst = iPkgDstPort7;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:473:3
	assign intTag[7].Pld = {iPkgPri7, iPkgFirAddr7, iPkgLen7, 4'h7};
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:474:3
	assign oPkgRdy7 = intTag[7].Rdy;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:476:3
	assign intTag[8].Vld = iPkgTagVld8;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:477:3
	assign intTag[8].Dst = iPkgDstPort8;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:478:3
	assign intTag[8].Pld = {iPkgPri8, iPkgFirAddr8, iPkgLen8, 4'h8};
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:479:3
	assign oPkgRdy8 = intTag[8].Rdy;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:481:3
	assign intTag[9].Vld = iPkgTagVld9;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:482:3
	assign intTag[9].Dst = iPkgDstPort9;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:483:3
	assign intTag[9].Pld = {iPkgPri9, iPkgFirAddr9, iPkgLen9, 4'h9};
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:484:3
	assign oPkgRdy9 = intTag[9].Rdy;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:486:3
	assign intTag[10].Vld = iPkgTagVld10;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:487:3
	assign intTag[10].Dst = iPkgDstPort10;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:488:3
	assign intTag[10].Pld = {iPkgPri10, iPkgFirAddr10, iPkgLen10, 4'ha};
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:489:3
	assign oPkgRdy10 = intTag[10].Rdy;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:491:3
	assign intTag[11].Vld = iPkgTagVld11;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:492:3
	assign intTag[11].Dst = iPkgDstPort11;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:493:3
	assign intTag[11].Pld = {iPkgPri11, iPkgFirAddr11, iPkgLen11, 4'hb};
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:494:3
	assign oPkgRdy11 = intTag[11].Rdy;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:496:3
	assign intTag[12].Vld = iPkgTagVld12;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:497:3
	assign intTag[12].Dst = iPkgDstPort12;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:498:3
	assign intTag[12].Pld = {iPkgPri12, iPkgFirAddr12, iPkgLen12, 4'hc};
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:499:3
	assign oPkgRdy12 = intTag[12].Rdy;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:501:3
	assign intTag[13].Vld = iPkgTagVld13;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:502:3
	assign intTag[13].Dst = iPkgDstPort13;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:503:3
	assign intTag[13].Pld = {iPkgPri13, iPkgFirAddr13, iPkgLen13, 4'hd};
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:504:3
	assign oPkgRdy13 = intTag[13].Rdy;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:506:3
	assign intTag[14].Vld = iPkgTagVld14;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:507:3
	assign intTag[14].Dst = iPkgDstPort14;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:508:3
	assign intTag[14].Pld = {iPkgPri14, iPkgFirAddr14, iPkgLen14, 4'he};
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:509:3
	assign oPkgRdy14 = intTag[14].Rdy;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:511:3
	assign intTag[15].Vld = iPkgTagVld15;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:512:3
	assign intTag[15].Dst = iPkgDstPort15;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:513:3
	assign intTag[15].Pld = {iPkgPri15, iPkgFirAddr15, iPkgLen15, 4'hf};
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:514:3
	assign oPkgRdy15 = intTag[15].Rdy;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:518:3
	wire [63:0] rdCmdDstPort;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:520:3
	assign oPkgFirAddrVld0 = intRdCmd[0].Vld;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:521:3
	assign intRdCmd[0].Rdy = iPkgFirAddrRdy0;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:522:3
	assign {oPkgFirAddr0, oPkgBlockNum0, rdCmdDstPort[60+:4], oPkgDrop0} = intRdCmd[0].Pld;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:524:3
	assign oPkgFirAddrVld1 = intRdCmd[1].Vld;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:525:3
	assign intRdCmd[1].Rdy = iPkgFirAddrRdy1;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:526:3
	assign {oPkgFirAddr1, oPkgBlockNum1, rdCmdDstPort[56+:4], oPkgDrop1} = intRdCmd[1].Pld;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:528:3
	assign oPkgFirAddrVld2 = intRdCmd[2].Vld;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:529:3
	assign intRdCmd[2].Rdy = iPkgFirAddrRdy2;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:530:3
	assign {oPkgFirAddr2, oPkgBlockNum2, rdCmdDstPort[52+:4], oPkgDrop2} = intRdCmd[2].Pld;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:532:3
	assign oPkgFirAddrVld3 = intRdCmd[3].Vld;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:533:3
	assign intRdCmd[3].Rdy = iPkgFirAddrRdy3;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:534:3
	assign {oPkgFirAddr3, oPkgBlockNum3, rdCmdDstPort[48+:4], oPkgDrop3} = intRdCmd[3].Pld;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:536:3
	assign oPkgFirAddrVld4 = intRdCmd[4].Vld;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:537:3
	assign intRdCmd[4].Rdy = iPkgFirAddrRdy4;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:538:3
	assign {oPkgFirAddr4, oPkgBlockNum4, rdCmdDstPort[44+:4], oPkgDrop4} = intRdCmd[4].Pld;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:540:3
	assign oPkgFirAddrVld5 = intRdCmd[5].Vld;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:541:3
	assign intRdCmd[5].Rdy = iPkgFirAddrRdy5;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:542:3
	assign {oPkgFirAddr5, oPkgBlockNum5, rdCmdDstPort[40+:4], oPkgDrop5} = intRdCmd[5].Pld;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:544:3
	assign oPkgFirAddrVld6 = intRdCmd[6].Vld;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:545:3
	assign intRdCmd[6].Rdy = iPkgFirAddrRdy6;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:546:3
	assign {oPkgFirAddr6, oPkgBlockNum6, rdCmdDstPort[36+:4], oPkgDrop6} = intRdCmd[6].Pld;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:548:3
	assign oPkgFirAddrVld7 = intRdCmd[7].Vld;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:549:3
	assign intRdCmd[7].Rdy = iPkgFirAddrRdy7;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:550:3
	assign {oPkgFirAddr7, oPkgBlockNum7, rdCmdDstPort[32+:4], oPkgDrop7} = intRdCmd[7].Pld;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:552:3
	assign oPkgFirAddrVld8 = intRdCmd[8].Vld;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:553:3
	assign intRdCmd[8].Rdy = iPkgFirAddrRdy8;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:554:3
	assign {oPkgFirAddr8, oPkgBlockNum8, rdCmdDstPort[28+:4], oPkgDrop8} = intRdCmd[8].Pld;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:556:3
	assign oPkgFirAddrVld9 = intRdCmd[9].Vld;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:557:3
	assign intRdCmd[9].Rdy = iPkgFirAddrRdy9;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:558:3
	assign {oPkgFirAddr9, oPkgBlockNum9, rdCmdDstPort[24+:4], oPkgDrop9} = intRdCmd[9].Pld;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:560:3
	assign oPkgFirAddrVld10 = intRdCmd[10].Vld;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:561:3
	assign intRdCmd[10].Rdy = iPkgFirAddrRdy10;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:562:3
	assign {oPkgFirAddr10, oPkgBlockNum10, rdCmdDstPort[20+:4], oPkgDrop10} = intRdCmd[10].Pld;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:564:3
	assign oPkgFirAddrVld11 = intRdCmd[11].Vld;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:565:3
	assign intRdCmd[11].Rdy = iPkgFirAddrRdy11;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:566:3
	assign {oPkgFirAddr11, oPkgBlockNum11, rdCmdDstPort[16+:4], oPkgDrop11} = intRdCmd[11].Pld;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:568:3
	assign oPkgFirAddrVld12 = intRdCmd[12].Vld;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:569:3
	assign intRdCmd[12].Rdy = iPkgFirAddrRdy12;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:570:3
	assign {oPkgFirAddr12, oPkgBlockNum12, rdCmdDstPort[12+:4], oPkgDrop12} = intRdCmd[12].Pld;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:572:3
	assign oPkgFirAddrVld13 = intRdCmd[13].Vld;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:573:3
	assign intRdCmd[13].Rdy = iPkgFirAddrRdy13;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:574:3
	assign {oPkgFirAddr13, oPkgBlockNum13, rdCmdDstPort[8+:4], oPkgDrop13} = intRdCmd[13].Pld;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:576:3
	assign oPkgFirAddrVld14 = intRdCmd[14].Vld;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:577:3
	assign intRdCmd[14].Rdy = iPkgFirAddrRdy14;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:578:3
	assign {oPkgFirAddr14, oPkgBlockNum14, rdCmdDstPort[4+:4], oPkgDrop14} = intRdCmd[14].Pld;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:580:3
	assign oPkgFirAddrVld15 = intRdCmd[15].Vld;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:581:3
	assign intRdCmd[15].Rdy = iPkgFirAddrRdy15;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:582:3
	assign {oPkgFirAddr15, oPkgBlockNum15, rdCmdDstPort[0+:4], oPkgDrop15} = intRdCmd[15].Pld;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:586:3
	assign intRdData[0].Vld = iWrrVld0;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:587:3
	assign intRdData[0].Pld = {iWrrData0, iWrrLast0};
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:588:3
	assign oWrrRdy0 = intRdData[0].Rdy;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:590:3
	assign intRdData[1].Vld = iWrrVld1;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:591:3
	assign intRdData[1].Pld = {iWrrData1, iWrrLast1};
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:592:3
	assign oWrrRdy1 = intRdData[1].Rdy;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:594:3
	assign intRdData[2].Vld = iWrrVld2;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:595:3
	assign intRdData[2].Pld = {iWrrData2, iWrrLast2};
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:596:3
	assign oWrrRdy2 = intRdData[2].Rdy;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:598:3
	assign intRdData[3].Vld = iWrrVld3;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:599:3
	assign intRdData[3].Pld = {iWrrData3, iWrrLast3};
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:600:3
	assign oWrrRdy3 = intRdData[3].Rdy;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:602:3
	assign intRdData[4].Vld = iWrrVld4;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:603:3
	assign intRdData[4].Pld = {iWrrData4, iWrrLast4};
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:604:3
	assign oWrrRdy4 = intRdData[4].Rdy;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:606:3
	assign intRdData[5].Vld = iWrrVld5;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:607:3
	assign intRdData[5].Pld = {iWrrData5, iWrrLast5};
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:608:3
	assign oWrrRdy5 = intRdData[5].Rdy;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:610:3
	assign intRdData[6].Vld = iWrrVld6;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:611:3
	assign intRdData[6].Pld = {iWrrData6, iWrrLast6};
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:612:3
	assign oWrrRdy6 = intRdData[6].Rdy;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:614:3
	assign intRdData[7].Vld = iWrrVld7;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:615:3
	assign intRdData[7].Pld = {iWrrData7, iWrrLast7};
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:616:3
	assign oWrrRdy7 = intRdData[7].Rdy;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:618:3
	assign intRdData[8].Vld = iWrrVld8;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:619:3
	assign intRdData[8].Pld = {iWrrData8, iWrrLast8};
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:620:3
	assign oWrrRdy8 = intRdData[8].Rdy;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:622:3
	assign intRdData[9].Vld = iWrrVld9;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:623:3
	assign intRdData[9].Pld = {iWrrData9, iWrrLast9};
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:624:3
	assign oWrrRdy9 = intRdData[9].Rdy;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:626:3
	assign intRdData[10].Vld = iWrrVld10;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:627:3
	assign intRdData[10].Pld = {iWrrData10, iWrrLast10};
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:628:3
	assign oWrrRdy10 = intRdData[10].Rdy;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:630:3
	assign intRdData[11].Vld = iWrrVld11;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:631:3
	assign intRdData[11].Pld = {iWrrData11, iWrrLast11};
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:632:3
	assign oWrrRdy11 = intRdData[11].Rdy;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:634:3
	assign intRdData[12].Vld = iWrrVld12;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:635:3
	assign intRdData[12].Pld = {iWrrData12, iWrrLast12};
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:636:3
	assign oWrrRdy12 = intRdData[12].Rdy;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:638:3
	assign intRdData[13].Vld = iWrrVld13;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:639:3
	assign intRdData[13].Pld = {iWrrData13, iWrrLast13};
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:640:3
	assign oWrrRdy13 = intRdData[13].Rdy;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:642:3
	assign intRdData[14].Vld = iWrrVld14;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:643:3
	assign intRdData[14].Pld = {iWrrData14, iWrrLast14};
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:644:3
	assign oWrrRdy14 = intRdData[14].Rdy;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:646:3
	assign intRdData[15].Vld = iWrrVld15;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:647:3
	assign intRdData[15].Pld = {iWrrData15, iWrrLast15};
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:648:3
	assign oWrrRdy15 = intRdData[15].Rdy;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:652:3
	wire [0:15] rdSop;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:653:3
	wire [0:15] rdEop;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:654:3
	wire [0:15] rdVld;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:655:3
	wire [511:0] rdData;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:656:3
	wire [0:15] rdRdy;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:657:3
	wire [0:15] rdLast;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:659:3
	assign oRdSop0 = rdSop[0];
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:660:3
	assign oRdEop0 = rdEop[0];
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:661:3
	assign oRdVld0 = rdVld[0];
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:662:3
	assign oRdData0 = rdData[480+:32];
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:663:3
	assign rdRdy[0] = iRdRdy0;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:664:3
	assign oRdLast0 = rdLast[0];
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:666:3
	assign oRdSop1 = rdSop[1];
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:667:3
	assign oRdEop1 = rdEop[1];
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:668:3
	assign oRdVld1 = rdVld[1];
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:669:3
	assign oRdData1 = rdData[448+:32];
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:670:3
	assign rdRdy[1] = iRdRdy1;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:671:3
	assign oRdLast1 = rdLast[1];
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:673:3
	assign oRdSop2 = rdSop[2];
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:674:3
	assign oRdEop2 = rdEop[2];
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:675:3
	assign oRdVld2 = rdVld[2];
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:676:3
	assign oRdData2 = rdData[416+:32];
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:677:3
	assign rdRdy[2] = iRdRdy2;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:678:3
	assign oRdLast2 = rdLast[2];
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:680:3
	assign oRdSop3 = rdSop[3];
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:681:3
	assign oRdEop3 = rdEop[3];
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:682:3
	assign oRdVld3 = rdVld[3];
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:683:3
	assign oRdData3 = rdData[384+:32];
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:684:3
	assign rdRdy[3] = iRdRdy3;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:685:3
	assign oRdLast3 = rdLast[3];
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:687:3
	assign oRdSop4 = rdSop[4];
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:688:3
	assign oRdEop4 = rdEop[4];
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:689:3
	assign oRdVld4 = rdVld[4];
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:690:3
	assign oRdData4 = rdData[352+:32];
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:691:3
	assign rdRdy[4] = iRdRdy4;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:692:3
	assign oRdLast4 = rdLast[4];
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:694:3
	assign oRdSop5 = rdSop[5];
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:695:3
	assign oRdEop5 = rdEop[5];
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:696:3
	assign oRdVld5 = rdVld[5];
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:697:3
	assign oRdData5 = rdData[320+:32];
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:698:3
	assign rdRdy[5] = iRdRdy5;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:699:3
	assign oRdLast5 = rdLast[5];
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:701:3
	assign oRdSop6 = rdSop[6];
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:702:3
	assign oRdEop6 = rdEop[6];
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:703:3
	assign oRdVld6 = rdVld[6];
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:704:3
	assign oRdData6 = rdData[288+:32];
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:705:3
	assign rdRdy[6] = iRdRdy6;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:706:3
	assign oRdLast6 = rdLast[6];
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:708:3
	assign oRdSop7 = rdSop[7];
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:709:3
	assign oRdEop7 = rdEop[7];
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:710:3
	assign oRdVld7 = rdVld[7];
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:711:3
	assign oRdData7 = rdData[256+:32];
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:712:3
	assign rdRdy[7] = iRdRdy7;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:713:3
	assign oRdLast7 = rdLast[7];
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:715:3
	assign oRdSop8 = rdSop[8];
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:716:3
	assign oRdEop8 = rdEop[8];
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:717:3
	assign oRdVld8 = rdVld[8];
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:718:3
	assign oRdData8 = rdData[224+:32];
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:719:3
	assign rdRdy[8] = iRdRdy8;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:720:3
	assign oRdLast8 = rdLast[8];
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:722:3
	assign oRdSop9 = rdSop[9];
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:723:3
	assign oRdEop9 = rdEop[9];
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:724:3
	assign oRdVld9 = rdVld[9];
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:725:3
	assign oRdData9 = rdData[192+:32];
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:726:3
	assign rdRdy[9] = iRdRdy9;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:727:3
	assign oRdLast9 = rdLast[9];
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:729:3
	assign oRdSop10 = rdSop[10];
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:730:3
	assign oRdEop10 = rdEop[10];
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:731:3
	assign oRdVld10 = rdVld[10];
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:732:3
	assign oRdData10 = rdData[160+:32];
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:733:3
	assign rdRdy[10] = iRdRdy10;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:734:3
	assign oRdLast10 = rdLast[10];
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:736:3
	assign oRdSop11 = rdSop[11];
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:737:3
	assign oRdEop11 = rdEop[11];
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:738:3
	assign oRdVld11 = rdVld[11];
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:739:3
	assign oRdData11 = rdData[128+:32];
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:740:3
	assign rdRdy[11] = iRdRdy11;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:741:3
	assign oRdLast11 = rdLast[11];
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:743:3
	assign oRdSop12 = rdSop[12];
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:744:3
	assign oRdEop12 = rdEop[12];
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:745:3
	assign oRdVld12 = rdVld[12];
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:746:3
	assign oRdData12 = rdData[96+:32];
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:747:3
	assign rdRdy[12] = iRdRdy12;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:748:3
	assign oRdLast12 = rdLast[12];
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:750:3
	assign oRdSop13 = rdSop[13];
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:751:3
	assign oRdEop13 = rdEop[13];
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:752:3
	assign oRdVld13 = rdVld[13];
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:753:3
	assign oRdData13 = rdData[64+:32];
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:754:3
	assign rdRdy[13] = iRdRdy13;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:755:3
	assign oRdLast13 = rdLast[13];
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:757:3
	assign oRdSop14 = rdSop[14];
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:758:3
	assign oRdEop14 = rdEop[14];
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:759:3
	assign oRdVld14 = rdVld[14];
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:760:3
	assign oRdData14 = rdData[32+:32];
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:761:3
	assign rdRdy[14] = iRdRdy14;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:762:3
	assign oRdLast14 = rdLast[14];
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:764:3
	assign oRdSop15 = rdSop[15];
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:765:3
	assign oRdEop15 = rdEop[15];
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:766:3
	assign oRdVld15 = rdVld[15];
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:767:3
	assign oRdData15 = rdData[0+:32];
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:768:3
	assign rdRdy[15] = iRdRdy15;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:769:3
	assign oRdLast15 = rdLast[15];
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:773:3
	wire [($clog2(WRR_WEIGHT_NUM) >= 0 ? (8 * ($clog2(WRR_WEIGHT_NUM) + 1)) - 1 : (8 * (1 - $clog2(WRR_WEIGHT_NUM))) + ($clog2(WRR_WEIGHT_NUM) - 1)):($clog2(WRR_WEIGHT_NUM) >= 0 ? 0 : $clog2(WRR_WEIGHT_NUM) + 0)] weightPld;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:775:3
	assign weightPld[($clog2(WRR_WEIGHT_NUM) >= 0 ? 0 : $clog2(WRR_WEIGHT_NUM)) + (7 * ($clog2(WRR_WEIGHT_NUM) >= 0 ? $clog2(WRR_WEIGHT_NUM) + 1 : 1 - $clog2(WRR_WEIGHT_NUM)))+:($clog2(WRR_WEIGHT_NUM) >= 0 ? $clog2(WRR_WEIGHT_NUM) + 1 : 1 - $clog2(WRR_WEIGHT_NUM))] = iWrrWeightPld0;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:776:3
	assign weightPld[($clog2(WRR_WEIGHT_NUM) >= 0 ? 0 : $clog2(WRR_WEIGHT_NUM)) + (6 * ($clog2(WRR_WEIGHT_NUM) >= 0 ? $clog2(WRR_WEIGHT_NUM) + 1 : 1 - $clog2(WRR_WEIGHT_NUM)))+:($clog2(WRR_WEIGHT_NUM) >= 0 ? $clog2(WRR_WEIGHT_NUM) + 1 : 1 - $clog2(WRR_WEIGHT_NUM))] = iWrrWeightPld1;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:777:3
	assign weightPld[($clog2(WRR_WEIGHT_NUM) >= 0 ? 0 : $clog2(WRR_WEIGHT_NUM)) + (5 * ($clog2(WRR_WEIGHT_NUM) >= 0 ? $clog2(WRR_WEIGHT_NUM) + 1 : 1 - $clog2(WRR_WEIGHT_NUM)))+:($clog2(WRR_WEIGHT_NUM) >= 0 ? $clog2(WRR_WEIGHT_NUM) + 1 : 1 - $clog2(WRR_WEIGHT_NUM))] = iWrrWeightPld2;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:778:3
	assign weightPld[($clog2(WRR_WEIGHT_NUM) >= 0 ? 0 : $clog2(WRR_WEIGHT_NUM)) + (4 * ($clog2(WRR_WEIGHT_NUM) >= 0 ? $clog2(WRR_WEIGHT_NUM) + 1 : 1 - $clog2(WRR_WEIGHT_NUM)))+:($clog2(WRR_WEIGHT_NUM) >= 0 ? $clog2(WRR_WEIGHT_NUM) + 1 : 1 - $clog2(WRR_WEIGHT_NUM))] = iWrrWeightPld3;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:779:3
	assign weightPld[($clog2(WRR_WEIGHT_NUM) >= 0 ? 0 : $clog2(WRR_WEIGHT_NUM)) + (3 * ($clog2(WRR_WEIGHT_NUM) >= 0 ? $clog2(WRR_WEIGHT_NUM) + 1 : 1 - $clog2(WRR_WEIGHT_NUM)))+:($clog2(WRR_WEIGHT_NUM) >= 0 ? $clog2(WRR_WEIGHT_NUM) + 1 : 1 - $clog2(WRR_WEIGHT_NUM))] = iWrrWeightPld4;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:780:3
	assign weightPld[($clog2(WRR_WEIGHT_NUM) >= 0 ? 0 : $clog2(WRR_WEIGHT_NUM)) + (2 * ($clog2(WRR_WEIGHT_NUM) >= 0 ? $clog2(WRR_WEIGHT_NUM) + 1 : 1 - $clog2(WRR_WEIGHT_NUM)))+:($clog2(WRR_WEIGHT_NUM) >= 0 ? $clog2(WRR_WEIGHT_NUM) + 1 : 1 - $clog2(WRR_WEIGHT_NUM))] = iWrrWeightPld5;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:781:3
	assign weightPld[($clog2(WRR_WEIGHT_NUM) >= 0 ? 0 : $clog2(WRR_WEIGHT_NUM)) + ($clog2(WRR_WEIGHT_NUM) >= 0 ? $clog2(WRR_WEIGHT_NUM) + 1 : 1 - $clog2(WRR_WEIGHT_NUM))+:($clog2(WRR_WEIGHT_NUM) >= 0 ? $clog2(WRR_WEIGHT_NUM) + 1 : 1 - $clog2(WRR_WEIGHT_NUM))] = iWrrWeightPld6;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:782:3
	assign weightPld[($clog2(WRR_WEIGHT_NUM) >= 0 ? 0 : $clog2(WRR_WEIGHT_NUM)) + 0+:($clog2(WRR_WEIGHT_NUM) >= 0 ? $clog2(WRR_WEIGHT_NUM) + 1 : 1 - $clog2(WRR_WEIGHT_NUM))] = iWrrWeightPld7;
	// Trace: src/src/rtl/design/svsrc/RdScheTopWrapper.sv:785:1
	// expanded module instance: U_RD_SCHE_TOP_SV
	localparam _bbase_F00F8_iTagIn = 0;
	localparam _bbase_F00F8_iRdDataIn = 0;
	localparam _bbase_F00F8_oRdCmdOut = 0;
	localparam _param_F00F8_PRI_DEPTH = PRI_DEPTH;
	localparam _param_F00F8_WRR_WEIGHT_NUM = WRR_WEIGHT_NUM;
	generate
		if (1) begin : U_RD_SCHE_TOP_SV
			// Trace: src/src/rtl/design/svsrc/RdScheTop.sv:3:13
			localparam PRI_DEPTH = _param_F00F8_PRI_DEPTH;
			// Trace: src/src/rtl/design/svsrc/RdScheTop.sv:4:13
			localparam WRR_WEIGHT_NUM = _param_F00F8_WRR_WEIGHT_NUM;
			// Trace: src/src/rtl/design/svsrc/RdScheTop.sv:6:13
			localparam PRI_NUM = 8;
			// Trace: src/src/rtl/design/svsrc/RdScheTop.sv:8:3
			wire iClk;
			// Trace: src/src/rtl/design/svsrc/RdScheTop.sv:9:3
			wire iRst_n;
			// Trace: src/src/rtl/design/svsrc/RdScheTop.sv:11:3
			localparam _mbase_iTagIn = 0;
			// Trace: src/src/rtl/design/svsrc/RdScheTop.sv:12:3
			localparam _mbase_iRdDataIn = 0;
			// Trace: src/src/rtl/design/svsrc/RdScheTop.sv:13:3
			localparam _mbase_oRdCmdOut = 0;
			// Trace: src/src/rtl/design/svsrc/RdScheTop.sv:15:3
			wire [0:15] oRdSop;
			// Trace: src/src/rtl/design/svsrc/RdScheTop.sv:16:3
			wire [0:15] oRdEop;
			// Trace: src/src/rtl/design/svsrc/RdScheTop.sv:17:3
			wire [0:15] oRdVld;
			// Trace: src/src/rtl/design/svsrc/RdScheTop.sv:18:3
			wire [511:0] oRdData;
			// Trace: src/src/rtl/design/svsrc/RdScheTop.sv:19:3
			wire [0:15] iRdRdy;
			// Trace: src/src/rtl/design/svsrc/RdScheTop.sv:20:3
			wire [0:15] oRdLast;
			// Trace: src/src/rtl/design/svsrc/RdScheTop.sv:22:3
			wire [($clog2(WRR_WEIGHT_NUM) >= 0 ? (8 * ($clog2(WRR_WEIGHT_NUM) + 1)) - 1 : (8 * (1 - $clog2(WRR_WEIGHT_NUM))) + ($clog2(WRR_WEIGHT_NUM) - 1)):($clog2(WRR_WEIGHT_NUM) >= 0 ? 0 : $clog2(WRR_WEIGHT_NUM) + 0)] iWeightPld;
			// Trace: src/src/rtl/design/svsrc/RdScheTop.sv:23:3
			wire [3:0] iWeightIdx;
			// Trace: src/src/rtl/design/svsrc/RdScheTop.sv:24:3
			wire iWeightLoad;
			// Trace: src/src/rtl/design/svsrc/RdScheTop.sv:26:3
			genvar _gv_i_9;
			// Trace: src/src/rtl/design/svsrc/RdScheTop.sv:28:3
			localparam TAG_WIDTH = 23;
			// Trace: src/src/rtl/design/svsrc/RdScheTop.sv:29:3
			localparam RDCMD_WIDTH = 21;
			// Trace: src/src/rtl/design/svsrc/RdScheTop.sv:30:3
			localparam RDDATA_WIDTH = 33;
			// Trace: src/src/rtl/design/svsrc/RdScheTop.sv:32:3
			// expanded interface instance: tagCrsbarOut
			localparam _param_BA01E_DW = TAG_WIDTH;
			localparam _param_BA01E_AW = 4;
			genvar _arr_BA01E;
			for (_arr_BA01E = 0; _arr_BA01E <= 15; _arr_BA01E = _arr_BA01E + 1) begin : tagCrsbarOut
				// Trace: src/src/rtl/design/svsrc/interface_list.sv:64:33
				localparam DW = _param_BA01E_DW;
				// Trace: src/src/rtl/design/svsrc/interface_list.sv:64:52
				localparam AW = _param_BA01E_AW;
				// Trace: src/src/rtl/design/svsrc/interface_list.sv:65:3
				wire [22:0] Pld;
				// Trace: src/src/rtl/design/svsrc/interface_list.sv:66:3
				wire [3:0] Dst;
				// Trace: src/src/rtl/design/svsrc/interface_list.sv:67:3
				wire Vld;
				// Trace: src/src/rtl/design/svsrc/interface_list.sv:68:3
				wire Rdy;
				// Trace: src/src/rtl/design/svsrc/interface_list.sv:69:3
				// Trace: src/src/rtl/design/svsrc/interface_list.sv:75:3
			end
			// Trace: src/src/rtl/design/svsrc/RdScheTop.sv:34:3
			// expanded interface instance: rdcmdCrsbarIn
			localparam _param_4DE78_DW = RDCMD_WIDTH;
			localparam _param_4DE78_AW = 4;
			genvar _arr_4DE78;
			for (_arr_4DE78 = 0; _arr_4DE78 <= 15; _arr_4DE78 = _arr_4DE78 + 1) begin : rdcmdCrsbarIn
				// Trace: src/src/rtl/design/svsrc/interface_list.sv:64:33
				localparam DW = _param_4DE78_DW;
				// Trace: src/src/rtl/design/svsrc/interface_list.sv:64:52
				localparam AW = _param_4DE78_AW;
				// Trace: src/src/rtl/design/svsrc/interface_list.sv:65:3
				wire [20:0] Pld;
				// Trace: src/src/rtl/design/svsrc/interface_list.sv:66:3
				wire [3:0] Dst;
				// Trace: src/src/rtl/design/svsrc/interface_list.sv:67:3
				wire Vld;
				// Trace: src/src/rtl/design/svsrc/interface_list.sv:68:3
				wire Rdy;
				// Trace: src/src/rtl/design/svsrc/interface_list.sv:69:3
				// Trace: src/src/rtl/design/svsrc/interface_list.sv:75:3
			end
			// Trace: src/src/rtl/design/svsrc/RdScheTop.sv:35:3
			// expanded interface instance: rdcmdCrsbarOut
			localparam _param_E7892_DW = RDCMD_WIDTH;
			localparam _param_E7892_AW = 4;
			genvar _arr_E7892;
			for (_arr_E7892 = 0; _arr_E7892 <= 15; _arr_E7892 = _arr_E7892 + 1) begin : rdcmdCrsbarOut
				// Trace: src/src/rtl/design/svsrc/interface_list.sv:64:33
				localparam DW = _param_E7892_DW;
				// Trace: src/src/rtl/design/svsrc/interface_list.sv:64:52
				localparam AW = _param_E7892_AW;
				// Trace: src/src/rtl/design/svsrc/interface_list.sv:65:3
				wire [20:0] Pld;
				// Trace: src/src/rtl/design/svsrc/interface_list.sv:66:3
				wire [3:0] Dst;
				// Trace: src/src/rtl/design/svsrc/interface_list.sv:67:3
				wire Vld;
				// Trace: src/src/rtl/design/svsrc/interface_list.sv:68:3
				wire Rdy;
				// Trace: src/src/rtl/design/svsrc/interface_list.sv:69:3
				// Trace: src/src/rtl/design/svsrc/interface_list.sv:75:3
			end
			// Trace: src/src/rtl/design/svsrc/RdScheTop.sv:37:3
			// expanded interface instance: rddataCrsbarIn
			localparam _param_CA251_DW = RDDATA_WIDTH;
			localparam _param_CA251_AW = 4;
			genvar _arr_CA251;
			for (_arr_CA251 = 0; _arr_CA251 <= 15; _arr_CA251 = _arr_CA251 + 1) begin : rddataCrsbarIn
				// Trace: src/src/rtl/design/svsrc/interface_list.sv:64:33
				localparam DW = _param_CA251_DW;
				// Trace: src/src/rtl/design/svsrc/interface_list.sv:64:52
				localparam AW = _param_CA251_AW;
				// Trace: src/src/rtl/design/svsrc/interface_list.sv:65:3
				wire [32:0] Pld;
				// Trace: src/src/rtl/design/svsrc/interface_list.sv:66:3
				wire [3:0] Dst;
				// Trace: src/src/rtl/design/svsrc/interface_list.sv:67:3
				wire Vld;
				// Trace: src/src/rtl/design/svsrc/interface_list.sv:68:3
				wire Rdy;
				// Trace: src/src/rtl/design/svsrc/interface_list.sv:69:3
				// Trace: src/src/rtl/design/svsrc/interface_list.sv:75:3
			end
			// Trace: src/src/rtl/design/svsrc/RdScheTop.sv:38:3
			// expanded interface instance: rddataCrsbarOut
			localparam _param_D6959_DW = RDDATA_WIDTH;
			localparam _param_D6959_AW = 4;
			genvar _arr_D6959;
			for (_arr_D6959 = 0; _arr_D6959 <= 15; _arr_D6959 = _arr_D6959 + 1) begin : rddataCrsbarOut
				// Trace: src/src/rtl/design/svsrc/interface_list.sv:64:33
				localparam DW = _param_D6959_DW;
				// Trace: src/src/rtl/design/svsrc/interface_list.sv:64:52
				localparam AW = _param_D6959_AW;
				// Trace: src/src/rtl/design/svsrc/interface_list.sv:65:3
				wire [32:0] Pld;
				// Trace: src/src/rtl/design/svsrc/interface_list.sv:66:3
				wire [3:0] Dst;
				// Trace: src/src/rtl/design/svsrc/interface_list.sv:67:3
				wire Vld;
				// Trace: src/src/rtl/design/svsrc/interface_list.sv:68:3
				wire Rdy;
				// Trace: src/src/rtl/design/svsrc/interface_list.sv:69:3
				// Trace: src/src/rtl/design/svsrc/interface_list.sv:75:3
			end
			// Trace: src/src/rtl/design/svsrc/RdScheTop.sv:40:3
			for (_gv_i_9 = 0; _gv_i_9 < 16; _gv_i_9 = _gv_i_9 + 1) begin : GEN_RDDST_LOCK
				localparam i = _gv_i_9;
				// Trace: src/src/rtl/design/svsrc/RdScheTop.sv:42:7
				// expanded module instance: U_RDDST_LOCK
				localparam _bbase_30E91_iRdCmdIn = _gv_i_9;
				localparam _bbase_30E91_iRdDataIn = _gv_i_9 + _mbase_iRdDataIn;
				localparam _bbase_30E91_oRdDataOut = _gv_i_9;
				if (1) begin : U_RDDST_LOCK
					// Trace: src/src/rtl/design/svsrc/RdDstLock.sv:27:3
					wire iClk;
					// Trace: src/src/rtl/design/svsrc/RdDstLock.sv:28:3
					wire iRst_n;
					// Trace: src/src/rtl/design/svsrc/RdDstLock.sv:30:3
					localparam _mbase_iRdDataIn = _bbase_30E91_iRdDataIn;
					// Trace: src/src/rtl/design/svsrc/RdDstLock.sv:31:3
					localparam _mbase_oRdDataOut = _bbase_30E91_oRdDataOut;
					// Trace: src/src/rtl/design/svsrc/RdDstLock.sv:32:3
					localparam _mbase_iRdCmdIn = _bbase_30E91_iRdCmdIn;
					// Trace: src/src/rtl/design/svsrc/RdDstLock.sv:35:3
					wire [3:0] rdCmdDstPort;
					// Trace: src/src/rtl/design/svsrc/RdDstLock.sv:36:3
					wire [15:0] rdCmdMsg;
					// Trace: src/src/rtl/design/svsrc/RdDstLock.sv:37:3
					wire rdCmdDrop;
					// Trace: src/src/rtl/design/svsrc/RdDstLock.sv:39:3
					reg [3:0] lockedDst;
					// Trace: src/src/rtl/design/svsrc/RdDstLock.sv:41:3
					assign {rdCmdMsg, rdCmdDstPort, rdCmdDrop} = RdScheTopWrapper.U_RD_SCHE_TOP_SV.rdcmdCrsbarOut[_mbase_iRdCmdIn].Pld;
					// Trace: src/src/rtl/design/svsrc/RdDstLock.sv:43:3
					always @(posedge iClk or negedge iRst_n)
						// Trace: src/src/rtl/design/svsrc/RdDstLock.sv:44:5
						if (!iRst_n)
							// Trace: src/src/rtl/design/svsrc/RdDstLock.sv:45:7
							lockedDst <= 'b0;
						else if ((RdScheTopWrapper.U_RD_SCHE_TOP_SV.rdcmdCrsbarOut[_mbase_iRdCmdIn].Vld && RdScheTopWrapper.U_RD_SCHE_TOP_SV.rdcmdCrsbarOut[_mbase_iRdCmdIn].Rdy) && !rdCmdDrop)
							// Trace: src/src/rtl/design/svsrc/RdDstLock.sv:47:7
							lockedDst <= rdCmdDstPort;
						else
							// Trace: src/src/rtl/design/svsrc/RdDstLock.sv:49:7
							lockedDst <= lockedDst;
					// Trace: src/src/rtl/design/svsrc/RdDstLock.sv:53:3
					assign RdScheTopWrapper.U_RD_SCHE_TOP_SV.rddataCrsbarIn[_mbase_oRdDataOut].Dst = lockedDst;
					// Trace: src/src/rtl/design/svsrc/RdDstLock.sv:54:3
					assign RdScheTopWrapper.U_RD_SCHE_TOP_SV.rddataCrsbarIn[_mbase_oRdDataOut].Pld = RdScheTopWrapper.intRdData[_mbase_iRdDataIn].Pld;
					// Trace: src/src/rtl/design/svsrc/RdDstLock.sv:55:3
					assign RdScheTopWrapper.U_RD_SCHE_TOP_SV.rddataCrsbarIn[_mbase_oRdDataOut].Vld = RdScheTopWrapper.intRdData[_mbase_iRdDataIn].Vld;
					// Trace: src/src/rtl/design/svsrc/RdDstLock.sv:56:3
					assign RdScheTopWrapper.intRdData[_mbase_iRdDataIn].Rdy = RdScheTopWrapper.U_RD_SCHE_TOP_SV.rddataCrsbarIn[_mbase_oRdDataOut].Rdy;
				end
				assign U_RDDST_LOCK.iClk = iClk;
				assign U_RDDST_LOCK.iRst_n = iRst_n;
				// Trace: src/src/rtl/design/svsrc/RdScheTop.sv:50:7
				assign rdcmdCrsbarOut[i].Rdy = RdScheTopWrapper.intRdCmd[i + _mbase_oRdCmdOut].Rdy;
				// Trace: src/src/rtl/design/svsrc/RdScheTop.sv:51:7
				assign RdScheTopWrapper.intRdCmd[i + _mbase_oRdCmdOut].Vld = rdcmdCrsbarOut[i].Vld;
				// Trace: src/src/rtl/design/svsrc/RdScheTop.sv:52:7
				assign RdScheTopWrapper.intRdCmd[i + _mbase_oRdCmdOut].Pld = rdcmdCrsbarOut[i].Pld;
				// Trace: src/src/rtl/design/svsrc/RdScheTop.sv:53:7
				assign RdScheTopWrapper.intRdCmd[i + _mbase_oRdCmdOut].Dst = rdcmdCrsbarOut[i].Dst;
			end
			// Trace: src/src/rtl/design/svsrc/RdScheTop.sv:58:3
			// expanded module instance: U_TAG_CRSBAR
			localparam _bbase_7E85F_iTagIn = 0;
			localparam _bbase_7E85F_oTagOut = 0;
			if (1) begin : U_TAG_CRSBAR
				// Trace: src/src/rtl/design/svsrc/DcpTag16x16.sv:27:3
				wire iClk;
				// Trace: src/src/rtl/design/svsrc/DcpTag16x16.sv:28:3
				wire iRst_n;
				// Trace: src/src/rtl/design/svsrc/DcpTag16x16.sv:30:3
				localparam _mbase_iTagIn = 0;
				// Trace: src/src/rtl/design/svsrc/DcpTag16x16.sv:31:3
				localparam _mbase_oTagOut = 0;
				// Trace: src/src/rtl/design/svsrc/DcpTag16x16.sv:33:3
				localparam CRSBAR_N = 4;
				// Trace: src/src/rtl/design/svsrc/DcpTag16x16.sv:34:3
				localparam CRSBAR_WIDTH = 23;
				// Trace: src/src/rtl/design/svsrc/DcpTag16x16.sv:36:3
				// expanded interface instance: switchOut
				localparam _param_CF9F8_DW = CRSBAR_WIDTH;
				localparam _param_CF9F8_AW = 4;
				genvar _arr_CF9F8;
				for (_arr_CF9F8 = 0; _arr_CF9F8 <= 3; _arr_CF9F8 = _arr_CF9F8 + 1) begin : switchOut
					// Trace: src/src/rtl/design/svsrc/interface_list.sv:64:33
					localparam DW = _param_CF9F8_DW;
					// Trace: src/src/rtl/design/svsrc/interface_list.sv:64:52
					localparam AW = _param_CF9F8_AW;
					// Trace: src/src/rtl/design/svsrc/interface_list.sv:65:3
					wire [22:0] Pld;
					// Trace: src/src/rtl/design/svsrc/interface_list.sv:66:3
					wire [3:0] Dst;
					// Trace: src/src/rtl/design/svsrc/interface_list.sv:67:3
					wire Vld;
					// Trace: src/src/rtl/design/svsrc/interface_list.sv:68:3
					wire Rdy;
					// Trace: src/src/rtl/design/svsrc/interface_list.sv:69:3
					// Trace: src/src/rtl/design/svsrc/interface_list.sv:75:3
				end
				// Trace: src/src/rtl/design/svsrc/DcpTag16x16.sv:37:3
				// expanded interface instance: routeIn
				localparam _param_37094_DW = CRSBAR_WIDTH;
				localparam _param_37094_AW = 4;
				genvar _arr_37094;
				for (_arr_37094 = 0; _arr_37094 <= 3; _arr_37094 = _arr_37094 + 1) begin : routeIn
					// Trace: src/src/rtl/design/svsrc/interface_list.sv:64:33
					localparam DW = _param_37094_DW;
					// Trace: src/src/rtl/design/svsrc/interface_list.sv:64:52
					localparam AW = _param_37094_AW;
					// Trace: src/src/rtl/design/svsrc/interface_list.sv:65:3
					wire [22:0] Pld;
					// Trace: src/src/rtl/design/svsrc/interface_list.sv:66:3
					wire [3:0] Dst;
					// Trace: src/src/rtl/design/svsrc/interface_list.sv:67:3
					wire Vld;
					// Trace: src/src/rtl/design/svsrc/interface_list.sv:68:3
					wire Rdy;
					// Trace: src/src/rtl/design/svsrc/interface_list.sv:69:3
					// Trace: src/src/rtl/design/svsrc/interface_list.sv:75:3
				end
				// Trace: src/src/rtl/design/svsrc/DcpTag16x16.sv:39:3
				// expanded interface instance: tagIn
				localparam _param_455CD_DW = CRSBAR_WIDTH;
				localparam _param_455CD_AW = 4;
				genvar _arr_455CD;
				for (_arr_455CD = 0; _arr_455CD <= 15; _arr_455CD = _arr_455CD + 1) begin : tagIn
					// Trace: src/src/rtl/design/svsrc/interface_list.sv:64:33
					localparam DW = _param_455CD_DW;
					// Trace: src/src/rtl/design/svsrc/interface_list.sv:64:52
					localparam AW = _param_455CD_AW;
					// Trace: src/src/rtl/design/svsrc/interface_list.sv:65:3
					wire [22:0] Pld;
					// Trace: src/src/rtl/design/svsrc/interface_list.sv:66:3
					wire [3:0] Dst;
					// Trace: src/src/rtl/design/svsrc/interface_list.sv:67:3
					wire Vld;
					// Trace: src/src/rtl/design/svsrc/interface_list.sv:68:3
					wire Rdy;
					// Trace: src/src/rtl/design/svsrc/interface_list.sv:69:3
					// Trace: src/src/rtl/design/svsrc/interface_list.sv:75:3
				end
				// Trace: src/src/rtl/design/svsrc/DcpTag16x16.sv:40:3
				// expanded interface instance: tagOut
				localparam _param_D8E37_DW = CRSBAR_WIDTH;
				localparam _param_D8E37_AW = 4;
				genvar _arr_D8E37;
				for (_arr_D8E37 = 0; _arr_D8E37 <= 15; _arr_D8E37 = _arr_D8E37 + 1) begin : tagOut
					// Trace: src/src/rtl/design/svsrc/interface_list.sv:64:33
					localparam DW = _param_D8E37_DW;
					// Trace: src/src/rtl/design/svsrc/interface_list.sv:64:52
					localparam AW = _param_D8E37_AW;
					// Trace: src/src/rtl/design/svsrc/interface_list.sv:65:3
					wire [22:0] Pld;
					// Trace: src/src/rtl/design/svsrc/interface_list.sv:66:3
					wire [3:0] Dst;
					// Trace: src/src/rtl/design/svsrc/interface_list.sv:67:3
					wire Vld;
					// Trace: src/src/rtl/design/svsrc/interface_list.sv:68:3
					wire Rdy;
					// Trace: src/src/rtl/design/svsrc/interface_list.sv:69:3
					// Trace: src/src/rtl/design/svsrc/interface_list.sv:75:3
				end
				// Trace: src/src/rtl/design/svsrc/DcpTag16x16.sv:42:3
				genvar _gv_i_5;
				// Trace: src/src/rtl/design/svsrc/DcpTag16x16.sv:44:3
				for (_gv_i_5 = 0; _gv_i_5 < 4; _gv_i_5 = _gv_i_5 + 1) begin : GEN_INPUT_SWITCH
					localparam i = _gv_i_5;
					// Trace: src/src/rtl/design/svsrc/DcpTag16x16.sv:46:7
					// expanded module instance: U_INPUT_SWITCH
					localparam _bbase_66B98_iDcpIn = 4 * _gv_i_5;
					localparam _bbase_66B98_oDcpOut = _gv_i_5;
					localparam _param_66B98_DW = CRSBAR_WIDTH;
					localparam _param_66B98_AW = 4;
					localparam _param_66B98_SNUM = 4;
					if (1) begin : U_INPUT_SWITCH
						// Trace: src/src/rtl/design/svsrc/DcpSwitchUnit.sv:28:13
						localparam DW = _param_66B98_DW;
						// Trace: src/src/rtl/design/svsrc/DcpSwitchUnit.sv:29:13
						localparam AW = _param_66B98_AW;
						// Trace: src/src/rtl/design/svsrc/DcpSwitchUnit.sv:30:13
						localparam SNUM = _param_66B98_SNUM;
						// Trace: src/src/rtl/design/svsrc/DcpSwitchUnit.sv:32:3
						wire iClk;
						// Trace: src/src/rtl/design/svsrc/DcpSwitchUnit.sv:33:3
						wire iRst_n;
						// Trace: src/src/rtl/design/svsrc/DcpSwitchUnit.sv:35:3
						localparam _mbase_iDcpIn = _bbase_66B98_iDcpIn;
						// Trace: src/src/rtl/design/svsrc/DcpSwitchUnit.sv:36:3
						localparam _mbase_oDcpOut = _bbase_66B98_oDcpOut;
						// Trace: src/src/rtl/design/svsrc/DcpSwitchUnit.sv:38:3
						wire [3:0] arbInReqArray;
						// Trace: src/src/rtl/design/svsrc/DcpSwitchUnit.sv:39:3
						wire [3:0] arbInGntArray;
						// Trace: src/src/rtl/design/svsrc/DcpSwitchUnit.sv:40:3
						wire [107:0] arbInPldArray;
						// Trace: src/src/rtl/design/svsrc/DcpSwitchUnit.sv:42:3
						wire arbOutReq;
						// Trace: src/src/rtl/design/svsrc/DcpSwitchUnit.sv:43:3
						wire arbOutGnt;
						// Trace: src/src/rtl/design/svsrc/DcpSwitchUnit.sv:44:3
						wire [26:0] arbOutPld;
						// Trace: src/src/rtl/design/svsrc/DcpSwitchUnit.sv:46:3
						genvar _gv_i_4;
						// Trace: src/src/rtl/design/svsrc/DcpSwitchUnit.sv:48:3
						for (_gv_i_4 = 0; _gv_i_4 < SNUM; _gv_i_4 = _gv_i_4 + 1) begin : GEN_INBUF
							localparam i = _gv_i_4;
							// Trace: src/src/rtl/design/svsrc/DcpSwitchUnit.sv:50:7
							gnrl_buf #(
								.DW(27),
								.CUT_RDY(1)
							) U_INBUF(
								.clk_i(iClk),
								.rst_n_i(iRst_n),
								.din_i({RdScheTopWrapper.U_RD_SCHE_TOP_SV.U_TAG_CRSBAR.tagIn[i + _mbase_iDcpIn].Dst, RdScheTopWrapper.U_RD_SCHE_TOP_SV.U_TAG_CRSBAR.tagIn[i + _mbase_iDcpIn].Pld}),
								.din_vld_i(RdScheTopWrapper.U_RD_SCHE_TOP_SV.U_TAG_CRSBAR.tagIn[i + _mbase_iDcpIn].Vld),
								.din_rdy_o(RdScheTopWrapper.U_RD_SCHE_TOP_SV.U_TAG_CRSBAR.tagIn[i + _mbase_iDcpIn].Rdy),
								.dout_o(arbInPldArray[i * 27+:27]),
								.dout_vld_o(arbInReqArray[i]),
								.dout_rdy_i(arbInGntArray[i])
							);
						end
						// Trace: src/src/rtl/design/svsrc/DcpSwitchUnit.sv:67:3
						rr_arb_tree #(
							.NumIn(SNUM),
							.DataWidth(27),
							.AxiVldRdy(1),
							.LockIn(0)
						) U_RR_ARB(
							.rst_ni(iRst_n),
							.clk_i(iClk),
							.req_i(arbInReqArray),
							.gnt_o(arbInGntArray),
							.data_i(arbInPldArray),
							.req_o(arbOutReq),
							.gnt_i(arbOutGnt),
							.data_o(arbOutPld)
						);
						// Trace: src/src/rtl/design/svsrc/DcpSwitchUnit.sv:86:3
						gnrl_buf #(
							.DW(27),
							.CUT_RDY(1)
						) U_INBUF(
							.clk_i(iClk),
							.rst_n_i(iRst_n),
							.din_i(arbOutPld),
							.din_vld_i(arbOutReq),
							.din_rdy_o(arbOutGnt),
							.dout_o({RdScheTopWrapper.U_RD_SCHE_TOP_SV.U_TAG_CRSBAR.switchOut[_mbase_oDcpOut].Dst, RdScheTopWrapper.U_RD_SCHE_TOP_SV.U_TAG_CRSBAR.switchOut[_mbase_oDcpOut].Pld}),
							.dout_vld_o(RdScheTopWrapper.U_RD_SCHE_TOP_SV.U_TAG_CRSBAR.switchOut[_mbase_oDcpOut].Vld),
							.dout_rdy_i(RdScheTopWrapper.U_RD_SCHE_TOP_SV.U_TAG_CRSBAR.switchOut[_mbase_oDcpOut].Rdy)
						);
					end
					assign U_INPUT_SWITCH.iClk = iClk;
					assign U_INPUT_SWITCH.iRst_n = iRst_n;
				end
				// Trace: src/src/rtl/design/svsrc/DcpTag16x16.sv:59:3
				// expanded module instance: U_CRSBAR
				localparam _bbase_509DC_iDcpIn = 0;
				localparam _bbase_509DC_oDcpOut = 0;
				localparam _param_509DC_DW = CRSBAR_WIDTH;
				localparam _param_509DC_AW = 4;
				localparam _param_509DC_N = 4;
				if (1) begin : U_CRSBAR
					// Trace: src/src/rtl/design/svsrc/DcpCrossbarNxN.sv:26:13
					localparam DW = _param_509DC_DW;
					// Trace: src/src/rtl/design/svsrc/DcpCrossbarNxN.sv:27:13
					localparam AW = _param_509DC_AW;
					// Trace: src/src/rtl/design/svsrc/DcpCrossbarNxN.sv:28:13
					localparam N = _param_509DC_N;
					// Trace: src/src/rtl/design/svsrc/DcpCrossbarNxN.sv:30:3
					wire iClk;
					// Trace: src/src/rtl/design/svsrc/DcpCrossbarNxN.sv:31:3
					wire iRst_n;
					// Trace: src/src/rtl/design/svsrc/DcpCrossbarNxN.sv:32:3
					localparam _mbase_iDcpIn = 0;
					// Trace: src/src/rtl/design/svsrc/DcpCrossbarNxN.sv:33:3
					localparam _mbase_oDcpOut = 0;
					// Trace: src/src/rtl/design/svsrc/DcpCrossbarNxN.sv:35:3
					// Trace: src/src/rtl/design/svsrc/DcpCrossbarNxN.sv:41:3
					// expanded interface instance: xbarCon
					localparam _param_7FFE1_DW = DW;
					localparam _param_7FFE1_AW = AW;
					genvar _arr_7FFE1;
					for (_arr_7FFE1 = 0; _arr_7FFE1 <= 15; _arr_7FFE1 = _arr_7FFE1 + 1) begin : xbarCon
						// Trace: src/src/rtl/design/svsrc/interface_list.sv:64:33
						localparam DW = _param_7FFE1_DW;
						// Trace: src/src/rtl/design/svsrc/interface_list.sv:64:52
						localparam AW = _param_7FFE1_AW;
						// Trace: src/src/rtl/design/svsrc/interface_list.sv:65:3
						wire [22:0] Pld;
						// Trace: src/src/rtl/design/svsrc/interface_list.sv:66:3
						wire [3:0] Dst;
						// Trace: src/src/rtl/design/svsrc/interface_list.sv:67:3
						wire Vld;
						// Trace: src/src/rtl/design/svsrc/interface_list.sv:68:3
						wire Rdy;
						// Trace: src/src/rtl/design/svsrc/interface_list.sv:69:3
						// Trace: src/src/rtl/design/svsrc/interface_list.sv:75:3
					end
					// Trace: src/src/rtl/design/svsrc/DcpCrossbarNxN.sv:42:3
					// expanded interface instance: xbarConT
					localparam _param_46BCA_DW = DW;
					localparam _param_46BCA_AW = AW;
					genvar _arr_46BCA;
					for (_arr_46BCA = 0; _arr_46BCA <= 15; _arr_46BCA = _arr_46BCA + 1) begin : xbarConT
						// Trace: src/src/rtl/design/svsrc/interface_list.sv:64:33
						localparam DW = _param_46BCA_DW;
						// Trace: src/src/rtl/design/svsrc/interface_list.sv:64:52
						localparam AW = _param_46BCA_AW;
						// Trace: src/src/rtl/design/svsrc/interface_list.sv:65:3
						wire [22:0] Pld;
						// Trace: src/src/rtl/design/svsrc/interface_list.sv:66:3
						wire [3:0] Dst;
						// Trace: src/src/rtl/design/svsrc/interface_list.sv:67:3
						wire Vld;
						// Trace: src/src/rtl/design/svsrc/interface_list.sv:68:3
						wire Rdy;
						// Trace: src/src/rtl/design/svsrc/interface_list.sv:69:3
						// Trace: src/src/rtl/design/svsrc/interface_list.sv:75:3
					end
					// Trace: src/src/rtl/design/svsrc/DcpCrossbarNxN.sv:44:3
					genvar _gv_i_1;
					// Trace: src/src/rtl/design/svsrc/DcpCrossbarNxN.sv:45:3
					genvar _gv_j_1;
					// Trace: src/src/rtl/design/svsrc/DcpCrossbarNxN.sv:46:3
					for (_gv_i_1 = 0; _gv_i_1 < N; _gv_i_1 = _gv_i_1 + 1) begin : GEN_XBAR_CON_TRANS_ROW
						localparam i = _gv_i_1;
						for (_gv_j_1 = 0; _gv_j_1 < N; _gv_j_1 = _gv_j_1 + 1) begin : GEN_XBAR_CON_TRANS_COL
							localparam j = _gv_j_1;
							// Trace: src/src/rtl/design/svsrc/DcpCrossbarNxN.sv:52:9
							assign xbarConT[(i * N) + j].Vld = xbarCon[(j * N) + i].Vld;
							// Trace: src/src/rtl/design/svsrc/DcpCrossbarNxN.sv:53:9
							assign xbarConT[(i * N) + j].Pld = xbarCon[(j * N) + i].Pld;
							// Trace: src/src/rtl/design/svsrc/DcpCrossbarNxN.sv:54:9
							assign xbarConT[(i * N) + j].Dst = xbarCon[(j * N) + i].Dst;
							// Trace: src/src/rtl/design/svsrc/DcpCrossbarNxN.sv:55:9
							assign xbarCon[(j * N) + i].Rdy = xbarConT[(i * N) + j].Rdy;
						end
					end
					// Trace: src/src/rtl/design/svsrc/DcpCrossbarNxN.sv:60:3
					for (_gv_i_1 = 0; _gv_i_1 < N; _gv_i_1 = _gv_i_1 + 1) begin : GEN_CON
						localparam i = _gv_i_1;
						// Trace: src/src/rtl/design/svsrc/DcpCrossbarNxN.sv:62:7
						// expanded module instance: U_ROUTEUNIT
						localparam _bbase_08BCB_iDcpIn = _gv_i_1 + _mbase_iDcpIn;
						localparam _bbase_08BCB_oDcpOut = N * _gv_i_1;
						localparam _param_08BCB_DW = DW;
						localparam _param_08BCB_AW = AW;
						localparam _param_08BCB_RNUM = N;
						if (1) begin : U_ROUTEUNIT
							reg _sv2v_0;
							// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:3:13
							localparam DW = _param_08BCB_DW;
							// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:4:13
							localparam AW = _param_08BCB_AW;
							// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:5:13
							localparam RNUM = _param_08BCB_RNUM;
							// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:7:3
							wire iClk;
							// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:8:3
							wire iRst_n;
							// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:10:3
							localparam _mbase_iDcpIn = _bbase_08BCB_iDcpIn;
							// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:11:3
							localparam _mbase_oDcpOut = _bbase_08BCB_oDcpOut;
							// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:14:3
							reg swiInRdy;
							// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:15:3
							wire swiInVld;
							// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:16:3
							wire [22:0] swiInPld;
							// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:17:3
							wire [3:0] swiInDst;
							// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:19:3
							reg [3:0] swiOutVld;
							// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:20:3
							wire [3:0] swiOutRdy;
							// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:22:3
							localparam IDLE = 1'b0;
							// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:23:3
							localparam GRANT = 1'b1;
							// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:25:3
							gnrl_buf #(
								.DW(27),
								.CUT_RDY(1)
							) U_INBUF(
								.clk_i(iClk),
								.rst_n_i(iRst_n),
								.din_i({RdScheTopWrapper.U_RD_SCHE_TOP_SV.U_TAG_CRSBAR.switchOut[_mbase_iDcpIn].Dst[3:0], RdScheTopWrapper.U_RD_SCHE_TOP_SV.U_TAG_CRSBAR.switchOut[_mbase_iDcpIn].Pld}),
								.din_vld_i(RdScheTopWrapper.U_RD_SCHE_TOP_SV.U_TAG_CRSBAR.switchOut[_mbase_iDcpIn].Vld),
								.din_rdy_o(RdScheTopWrapper.U_RD_SCHE_TOP_SV.U_TAG_CRSBAR.switchOut[_mbase_iDcpIn].Rdy),
								.dout_o({swiInDst, swiInPld}),
								.dout_vld_o(swiInVld),
								.dout_rdy_i(swiInRdy)
							);
							// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:39:3
							genvar _gv_i_3;
							// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:40:3
							for (_gv_i_3 = 0; _gv_i_3 < RNUM; _gv_i_3 = _gv_i_3 + 1) begin : GEN_ROUTE
								localparam i = _gv_i_3;
								// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:42:7
								always @(*) begin
									if (_sv2v_0)
										;
									// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:44:9
									if (swiInVld && (swiInDst[3-:2] == i))
										// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:45:11
										swiOutVld[i] = swiInVld;
									else
										// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:47:11
										swiOutVld[i] = 1'b0;
								end
							end
							// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:53:3
							reg signed [31:0] j;
							// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:54:3
							always @(*) begin
								if (_sv2v_0)
									;
								// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:55:5
								if (swiInVld) begin
									begin
										// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:56:7
										for (j = 0; j < RNUM; j = j + 1)
											begin
												// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:58:9
												if (swiInDst[3-:2] == j)
													// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:59:11
													swiInRdy = swiOutRdy[j];
											end
									end
								end
								else
									// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:63:7
									swiInRdy = 1'b0;
							end
							// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:67:3
							for (_gv_i_3 = 0; _gv_i_3 < RNUM; _gv_i_3 = _gv_i_3 + 1) begin : GEN_OUTBUF
								localparam i = _gv_i_3;
								// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:69:7
								gnrl_buf #(
									.DW(27),
									.CUT_RDY(1)
								) U_OUTBUF(
									.clk_i(iClk),
									.rst_n_i(iRst_n),
									.din_i({swiInDst, swiInPld}),
									.din_vld_i(swiOutVld[i]),
									.din_rdy_o(swiOutRdy[i]),
									.dout_o({RdScheTopWrapper.U_RD_SCHE_TOP_SV.U_TAG_CRSBAR.U_CRSBAR.xbarCon[i + _mbase_oDcpOut].Dst[3:0], RdScheTopWrapper.U_RD_SCHE_TOP_SV.U_TAG_CRSBAR.U_CRSBAR.xbarCon[i + _mbase_oDcpOut].Pld}),
									.dout_vld_o(RdScheTopWrapper.U_RD_SCHE_TOP_SV.U_TAG_CRSBAR.U_CRSBAR.xbarCon[i + _mbase_oDcpOut].Vld),
									.dout_rdy_i(RdScheTopWrapper.U_RD_SCHE_TOP_SV.U_TAG_CRSBAR.U_CRSBAR.xbarCon[i + _mbase_oDcpOut].Rdy)
								);
							end
							initial _sv2v_0 = 0;
						end
						assign U_ROUTEUNIT.iClk = iClk;
						assign U_ROUTEUNIT.iRst_n = iRst_n;
						// Trace: src/src/rtl/design/svsrc/DcpCrossbarNxN.sv:72:7
						// expanded module instance: U_SWITCHUNIT
						localparam _bbase_C87B5_iDcpIn = N * _gv_i_1;
						localparam _bbase_C87B5_oDcpOut = _gv_i_1 + _mbase_oDcpOut;
						localparam _param_C87B5_DW = DW;
						localparam _param_C87B5_AW = AW;
						localparam _param_C87B5_SNUM = N;
						if (1) begin : U_SWITCHUNIT
							// Trace: src/src/rtl/design/svsrc/DcpSwitchUnit.sv:28:13
							localparam DW = _param_C87B5_DW;
							// Trace: src/src/rtl/design/svsrc/DcpSwitchUnit.sv:29:13
							localparam AW = _param_C87B5_AW;
							// Trace: src/src/rtl/design/svsrc/DcpSwitchUnit.sv:30:13
							localparam SNUM = _param_C87B5_SNUM;
							// Trace: src/src/rtl/design/svsrc/DcpSwitchUnit.sv:32:3
							wire iClk;
							// Trace: src/src/rtl/design/svsrc/DcpSwitchUnit.sv:33:3
							wire iRst_n;
							// Trace: src/src/rtl/design/svsrc/DcpSwitchUnit.sv:35:3
							localparam _mbase_iDcpIn = _bbase_C87B5_iDcpIn;
							// Trace: src/src/rtl/design/svsrc/DcpSwitchUnit.sv:36:3
							localparam _mbase_oDcpOut = _bbase_C87B5_oDcpOut;
							// Trace: src/src/rtl/design/svsrc/DcpSwitchUnit.sv:38:3
							wire [3:0] arbInReqArray;
							// Trace: src/src/rtl/design/svsrc/DcpSwitchUnit.sv:39:3
							wire [3:0] arbInGntArray;
							// Trace: src/src/rtl/design/svsrc/DcpSwitchUnit.sv:40:3
							wire [107:0] arbInPldArray;
							// Trace: src/src/rtl/design/svsrc/DcpSwitchUnit.sv:42:3
							wire arbOutReq;
							// Trace: src/src/rtl/design/svsrc/DcpSwitchUnit.sv:43:3
							wire arbOutGnt;
							// Trace: src/src/rtl/design/svsrc/DcpSwitchUnit.sv:44:3
							wire [26:0] arbOutPld;
							// Trace: src/src/rtl/design/svsrc/DcpSwitchUnit.sv:46:3
							genvar _gv_i_4;
							// Trace: src/src/rtl/design/svsrc/DcpSwitchUnit.sv:48:3
							for (_gv_i_4 = 0; _gv_i_4 < SNUM; _gv_i_4 = _gv_i_4 + 1) begin : GEN_INBUF
								localparam i = _gv_i_4;
								// Trace: src/src/rtl/design/svsrc/DcpSwitchUnit.sv:50:7
								gnrl_buf #(
									.DW(27),
									.CUT_RDY(1)
								) U_INBUF(
									.clk_i(iClk),
									.rst_n_i(iRst_n),
									.din_i({RdScheTopWrapper.U_RD_SCHE_TOP_SV.U_TAG_CRSBAR.U_CRSBAR.xbarConT[i + _mbase_iDcpIn].Dst, RdScheTopWrapper.U_RD_SCHE_TOP_SV.U_TAG_CRSBAR.U_CRSBAR.xbarConT[i + _mbase_iDcpIn].Pld}),
									.din_vld_i(RdScheTopWrapper.U_RD_SCHE_TOP_SV.U_TAG_CRSBAR.U_CRSBAR.xbarConT[i + _mbase_iDcpIn].Vld),
									.din_rdy_o(RdScheTopWrapper.U_RD_SCHE_TOP_SV.U_TAG_CRSBAR.U_CRSBAR.xbarConT[i + _mbase_iDcpIn].Rdy),
									.dout_o(arbInPldArray[i * 27+:27]),
									.dout_vld_o(arbInReqArray[i]),
									.dout_rdy_i(arbInGntArray[i])
								);
							end
							// Trace: src/src/rtl/design/svsrc/DcpSwitchUnit.sv:67:3
							rr_arb_tree #(
								.NumIn(SNUM),
								.DataWidth(27),
								.AxiVldRdy(1),
								.LockIn(0)
							) U_RR_ARB(
								.rst_ni(iRst_n),
								.clk_i(iClk),
								.req_i(arbInReqArray),
								.gnt_o(arbInGntArray),
								.data_i(arbInPldArray),
								.req_o(arbOutReq),
								.gnt_i(arbOutGnt),
								.data_o(arbOutPld)
							);
							// Trace: src/src/rtl/design/svsrc/DcpSwitchUnit.sv:86:3
							gnrl_buf #(
								.DW(27),
								.CUT_RDY(1)
							) U_INBUF(
								.clk_i(iClk),
								.rst_n_i(iRst_n),
								.din_i(arbOutPld),
								.din_vld_i(arbOutReq),
								.din_rdy_o(arbOutGnt),
								.dout_o({RdScheTopWrapper.U_RD_SCHE_TOP_SV.U_TAG_CRSBAR.routeIn[_mbase_oDcpOut].Dst, RdScheTopWrapper.U_RD_SCHE_TOP_SV.U_TAG_CRSBAR.routeIn[_mbase_oDcpOut].Pld}),
								.dout_vld_o(RdScheTopWrapper.U_RD_SCHE_TOP_SV.U_TAG_CRSBAR.routeIn[_mbase_oDcpOut].Vld),
								.dout_rdy_i(RdScheTopWrapper.U_RD_SCHE_TOP_SV.U_TAG_CRSBAR.routeIn[_mbase_oDcpOut].Rdy)
							);
						end
						assign U_SWITCHUNIT.iClk = iClk;
						assign U_SWITCHUNIT.iRst_n = iRst_n;
					end
				end
				assign U_CRSBAR.iClk = iClk;
				assign U_CRSBAR.iRst_n = iRst_n;
				// Trace: src/src/rtl/design/svsrc/DcpTag16x16.sv:70:3
				for (_gv_i_5 = 0; _gv_i_5 < 4; _gv_i_5 = _gv_i_5 + 1) begin : GEN_OUTPUT_ROUTE
					localparam i = _gv_i_5;
					// Trace: src/src/rtl/design/svsrc/DcpTag16x16.sv:72:7
					// expanded module instance: U_OUTPUT_ROUTE
					localparam _bbase_37972_iDcpIn = _gv_i_5;
					localparam _bbase_37972_oDcpOut = 4 * _gv_i_5;
					localparam _param_37972_DW = CRSBAR_WIDTH;
					localparam _param_37972_AW = 2;
					localparam _param_37972_RNUM = 4;
					if (1) begin : U_OUTPUT_ROUTE
						reg _sv2v_0;
						// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:3:13
						localparam DW = _param_37972_DW;
						// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:4:13
						localparam AW = _param_37972_AW;
						// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:5:13
						localparam RNUM = _param_37972_RNUM;
						// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:7:3
						wire iClk;
						// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:8:3
						wire iRst_n;
						// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:10:3
						localparam _mbase_iDcpIn = _bbase_37972_iDcpIn;
						// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:11:3
						localparam _mbase_oDcpOut = _bbase_37972_oDcpOut;
						// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:14:3
						reg swiInRdy;
						// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:15:3
						wire swiInVld;
						// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:16:3
						wire [22:0] swiInPld;
						// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:17:3
						wire [1:0] swiInDst;
						// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:19:3
						reg [3:0] swiOutVld;
						// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:20:3
						wire [3:0] swiOutRdy;
						// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:22:3
						localparam IDLE = 1'b0;
						// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:23:3
						localparam GRANT = 1'b1;
						// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:25:3
						gnrl_buf #(
							.DW(25),
							.CUT_RDY(1)
						) U_INBUF(
							.clk_i(iClk),
							.rst_n_i(iRst_n),
							.din_i({RdScheTopWrapper.U_RD_SCHE_TOP_SV.U_TAG_CRSBAR.routeIn[_mbase_iDcpIn].Dst[1:0], RdScheTopWrapper.U_RD_SCHE_TOP_SV.U_TAG_CRSBAR.routeIn[_mbase_iDcpIn].Pld}),
							.din_vld_i(RdScheTopWrapper.U_RD_SCHE_TOP_SV.U_TAG_CRSBAR.routeIn[_mbase_iDcpIn].Vld),
							.din_rdy_o(RdScheTopWrapper.U_RD_SCHE_TOP_SV.U_TAG_CRSBAR.routeIn[_mbase_iDcpIn].Rdy),
							.dout_o({swiInDst, swiInPld}),
							.dout_vld_o(swiInVld),
							.dout_rdy_i(swiInRdy)
						);
						// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:39:3
						genvar _gv_i_3;
						// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:40:3
						for (_gv_i_3 = 0; _gv_i_3 < RNUM; _gv_i_3 = _gv_i_3 + 1) begin : GEN_ROUTE
							localparam i = _gv_i_3;
							// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:42:7
							always @(*) begin
								if (_sv2v_0)
									;
								// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:44:9
								if (swiInVld && (swiInDst[1-:2] == i))
									// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:45:11
									swiOutVld[i] = swiInVld;
								else
									// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:47:11
									swiOutVld[i] = 1'b0;
							end
						end
						// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:53:3
						reg signed [31:0] j;
						// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:54:3
						always @(*) begin
							if (_sv2v_0)
								;
							// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:55:5
							if (swiInVld) begin
								begin
									// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:56:7
									for (j = 0; j < RNUM; j = j + 1)
										begin
											// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:58:9
											if (swiInDst[1-:2] == j)
												// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:59:11
												swiInRdy = swiOutRdy[j];
										end
								end
							end
							else
								// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:63:7
								swiInRdy = 1'b0;
						end
						// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:67:3
						for (_gv_i_3 = 0; _gv_i_3 < RNUM; _gv_i_3 = _gv_i_3 + 1) begin : GEN_OUTBUF
							localparam i = _gv_i_3;
							// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:69:7
							gnrl_buf #(
								.DW(25),
								.CUT_RDY(1)
							) U_OUTBUF(
								.clk_i(iClk),
								.rst_n_i(iRst_n),
								.din_i({swiInDst, swiInPld}),
								.din_vld_i(swiOutVld[i]),
								.din_rdy_o(swiOutRdy[i]),
								.dout_o({RdScheTopWrapper.U_RD_SCHE_TOP_SV.U_TAG_CRSBAR.tagOut[i + _mbase_oDcpOut].Dst[1:0], RdScheTopWrapper.U_RD_SCHE_TOP_SV.U_TAG_CRSBAR.tagOut[i + _mbase_oDcpOut].Pld}),
								.dout_vld_o(RdScheTopWrapper.U_RD_SCHE_TOP_SV.U_TAG_CRSBAR.tagOut[i + _mbase_oDcpOut].Vld),
								.dout_rdy_i(RdScheTopWrapper.U_RD_SCHE_TOP_SV.U_TAG_CRSBAR.tagOut[i + _mbase_oDcpOut].Rdy)
							);
						end
						initial _sv2v_0 = 0;
					end
					assign U_OUTPUT_ROUTE.iClk = iClk;
					assign U_OUTPUT_ROUTE.iRst_n = iRst_n;
				end
				// Trace: src/src/rtl/design/svsrc/DcpTag16x16.sv:86:3
				for (_gv_i_5 = 0; _gv_i_5 < 16; _gv_i_5 = _gv_i_5 + 1) begin : GENCON
					localparam i = _gv_i_5;
					// Trace: src/src/rtl/design/svsrc/DcpTag16x16.sv:88:7
					assign tagOut[i].Rdy = RdScheTopWrapper.U_RD_SCHE_TOP_SV.tagCrsbarOut[i + _mbase_oTagOut].Rdy;
					// Trace: src/src/rtl/design/svsrc/DcpTag16x16.sv:89:7
					assign RdScheTopWrapper.U_RD_SCHE_TOP_SV.tagCrsbarOut[i + _mbase_oTagOut].Pld = tagOut[i].Pld;
					// Trace: src/src/rtl/design/svsrc/DcpTag16x16.sv:90:7
					assign RdScheTopWrapper.U_RD_SCHE_TOP_SV.tagCrsbarOut[i + _mbase_oTagOut].Vld = tagOut[i].Vld;
					// Trace: src/src/rtl/design/svsrc/DcpTag16x16.sv:91:7
					assign RdScheTopWrapper.U_RD_SCHE_TOP_SV.tagCrsbarOut[i + _mbase_oTagOut].Dst = tagOut[i].Dst;
					// Trace: src/src/rtl/design/svsrc/DcpTag16x16.sv:93:7
					assign RdScheTopWrapper.intTag[i + _mbase_iTagIn].Rdy = tagIn[i].Rdy;
					// Trace: src/src/rtl/design/svsrc/DcpTag16x16.sv:94:7
					assign tagIn[i].Pld = RdScheTopWrapper.intTag[i + _mbase_iTagIn].Pld;
					// Trace: src/src/rtl/design/svsrc/DcpTag16x16.sv:95:7
					assign tagIn[i].Vld = RdScheTopWrapper.intTag[i + _mbase_iTagIn].Vld;
					// Trace: src/src/rtl/design/svsrc/DcpTag16x16.sv:96:7
					assign tagIn[i].Dst = RdScheTopWrapper.intTag[i + _mbase_iTagIn].Dst;
				end
			end
			assign U_TAG_CRSBAR.iClk = iClk;
			assign U_TAG_CRSBAR.iRst_n = iRst_n;
			// Trace: src/src/rtl/design/svsrc/RdScheTop.sv:65:3
			// expanded module instance: U_RDDATA_CRSBAR
			localparam _bbase_3A305_iRdDataIn = 0;
			localparam _bbase_3A305_oRdDataOut = 0;
			if (1) begin : U_RDDATA_CRSBAR
				// Trace: src/src/rtl/design/svsrc/DcpRdData16x16.sv:4:3
				wire iClk;
				// Trace: src/src/rtl/design/svsrc/DcpRdData16x16.sv:5:3
				wire iRst_n;
				// Trace: src/src/rtl/design/svsrc/DcpRdData16x16.sv:7:3
				localparam _mbase_iRdDataIn = 0;
				// Trace: src/src/rtl/design/svsrc/DcpRdData16x16.sv:8:3
				localparam _mbase_oRdDataOut = 0;
				// Trace: src/src/rtl/design/svsrc/DcpRdData16x16.sv:11:3
				localparam CRSBAR_WIDTH = 33;
				// Trace: src/src/rtl/design/svsrc/DcpRdData16x16.sv:78:3
				// expanded module instance: U_CRSBAR
				localparam _bbase_509DC_iDcpIn = 0;
				localparam _bbase_509DC_oDcpOut = 0;
				localparam _param_509DC_DW = CRSBAR_WIDTH;
				localparam _param_509DC_AW = 4;
				localparam _param_509DC_N = 16;
				if (1) begin : U_CRSBAR
					// Trace: src/src/rtl/design/svsrc/DcpCrossbarNxN.sv:26:13
					localparam DW = _param_509DC_DW;
					// Trace: src/src/rtl/design/svsrc/DcpCrossbarNxN.sv:27:13
					localparam AW = _param_509DC_AW;
					// Trace: src/src/rtl/design/svsrc/DcpCrossbarNxN.sv:28:13
					localparam N = _param_509DC_N;
					// Trace: src/src/rtl/design/svsrc/DcpCrossbarNxN.sv:30:3
					wire iClk;
					// Trace: src/src/rtl/design/svsrc/DcpCrossbarNxN.sv:31:3
					wire iRst_n;
					// Trace: src/src/rtl/design/svsrc/DcpCrossbarNxN.sv:32:3
					localparam _mbase_iDcpIn = 0;
					// Trace: src/src/rtl/design/svsrc/DcpCrossbarNxN.sv:33:3
					localparam _mbase_oDcpOut = 0;
					// Trace: src/src/rtl/design/svsrc/DcpCrossbarNxN.sv:35:3
					// Trace: src/src/rtl/design/svsrc/DcpCrossbarNxN.sv:41:3
					// expanded interface instance: xbarCon
					localparam _param_7FFE1_DW = DW;
					localparam _param_7FFE1_AW = AW;
					genvar _arr_7FFE1;
					for (_arr_7FFE1 = 0; _arr_7FFE1 <= 255; _arr_7FFE1 = _arr_7FFE1 + 1) begin : xbarCon
						// Trace: src/src/rtl/design/svsrc/interface_list.sv:64:33
						localparam DW = _param_7FFE1_DW;
						// Trace: src/src/rtl/design/svsrc/interface_list.sv:64:52
						localparam AW = _param_7FFE1_AW;
						// Trace: src/src/rtl/design/svsrc/interface_list.sv:65:3
						wire [32:0] Pld;
						// Trace: src/src/rtl/design/svsrc/interface_list.sv:66:3
						wire [3:0] Dst;
						// Trace: src/src/rtl/design/svsrc/interface_list.sv:67:3
						wire Vld;
						// Trace: src/src/rtl/design/svsrc/interface_list.sv:68:3
						wire Rdy;
						// Trace: src/src/rtl/design/svsrc/interface_list.sv:69:3
						// Trace: src/src/rtl/design/svsrc/interface_list.sv:75:3
					end
					// Trace: src/src/rtl/design/svsrc/DcpCrossbarNxN.sv:42:3
					// expanded interface instance: xbarConT
					localparam _param_46BCA_DW = DW;
					localparam _param_46BCA_AW = AW;
					genvar _arr_46BCA;
					for (_arr_46BCA = 0; _arr_46BCA <= 255; _arr_46BCA = _arr_46BCA + 1) begin : xbarConT
						// Trace: src/src/rtl/design/svsrc/interface_list.sv:64:33
						localparam DW = _param_46BCA_DW;
						// Trace: src/src/rtl/design/svsrc/interface_list.sv:64:52
						localparam AW = _param_46BCA_AW;
						// Trace: src/src/rtl/design/svsrc/interface_list.sv:65:3
						wire [32:0] Pld;
						// Trace: src/src/rtl/design/svsrc/interface_list.sv:66:3
						wire [3:0] Dst;
						// Trace: src/src/rtl/design/svsrc/interface_list.sv:67:3
						wire Vld;
						// Trace: src/src/rtl/design/svsrc/interface_list.sv:68:3
						wire Rdy;
						// Trace: src/src/rtl/design/svsrc/interface_list.sv:69:3
						// Trace: src/src/rtl/design/svsrc/interface_list.sv:75:3
					end
					// Trace: src/src/rtl/design/svsrc/DcpCrossbarNxN.sv:44:3
					genvar _gv_i_1;
					// Trace: src/src/rtl/design/svsrc/DcpCrossbarNxN.sv:45:3
					genvar _gv_j_1;
					// Trace: src/src/rtl/design/svsrc/DcpCrossbarNxN.sv:46:3
					for (_gv_i_1 = 0; _gv_i_1 < N; _gv_i_1 = _gv_i_1 + 1) begin : GEN_XBAR_CON_TRANS_ROW
						localparam i = _gv_i_1;
						for (_gv_j_1 = 0; _gv_j_1 < N; _gv_j_1 = _gv_j_1 + 1) begin : GEN_XBAR_CON_TRANS_COL
							localparam j = _gv_j_1;
							// Trace: src/src/rtl/design/svsrc/DcpCrossbarNxN.sv:52:9
							assign xbarConT[(i * N) + j].Vld = xbarCon[(j * N) + i].Vld;
							// Trace: src/src/rtl/design/svsrc/DcpCrossbarNxN.sv:53:9
							assign xbarConT[(i * N) + j].Pld = xbarCon[(j * N) + i].Pld;
							// Trace: src/src/rtl/design/svsrc/DcpCrossbarNxN.sv:54:9
							assign xbarConT[(i * N) + j].Dst = xbarCon[(j * N) + i].Dst;
							// Trace: src/src/rtl/design/svsrc/DcpCrossbarNxN.sv:55:9
							assign xbarCon[(j * N) + i].Rdy = xbarConT[(i * N) + j].Rdy;
						end
					end
					// Trace: src/src/rtl/design/svsrc/DcpCrossbarNxN.sv:60:3
					for (_gv_i_1 = 0; _gv_i_1 < N; _gv_i_1 = _gv_i_1 + 1) begin : GEN_CON
						localparam i = _gv_i_1;
						// Trace: src/src/rtl/design/svsrc/DcpCrossbarNxN.sv:62:7
						// expanded module instance: U_ROUTEUNIT
						localparam _bbase_08BCB_iDcpIn = _gv_i_1 + _mbase_iDcpIn;
						localparam _bbase_08BCB_oDcpOut = N * _gv_i_1;
						localparam _param_08BCB_DW = DW;
						localparam _param_08BCB_AW = AW;
						localparam _param_08BCB_RNUM = N;
						if (1) begin : U_ROUTEUNIT
							reg _sv2v_0;
							// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:3:13
							localparam DW = _param_08BCB_DW;
							// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:4:13
							localparam AW = _param_08BCB_AW;
							// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:5:13
							localparam RNUM = _param_08BCB_RNUM;
							// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:7:3
							wire iClk;
							// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:8:3
							wire iRst_n;
							// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:10:3
							localparam _mbase_iDcpIn = _bbase_08BCB_iDcpIn;
							// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:11:3
							localparam _mbase_oDcpOut = _bbase_08BCB_oDcpOut;
							// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:14:3
							reg swiInRdy;
							// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:15:3
							wire swiInVld;
							// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:16:3
							wire [32:0] swiInPld;
							// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:17:3
							wire [3:0] swiInDst;
							// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:19:3
							reg [15:0] swiOutVld;
							// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:20:3
							wire [15:0] swiOutRdy;
							// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:22:3
							localparam IDLE = 1'b0;
							// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:23:3
							localparam GRANT = 1'b1;
							// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:25:3
							gnrl_buf #(
								.DW(37),
								.CUT_RDY(1)
							) U_INBUF(
								.clk_i(iClk),
								.rst_n_i(iRst_n),
								.din_i({RdScheTopWrapper.U_RD_SCHE_TOP_SV.rddataCrsbarIn[_mbase_iDcpIn].Dst[3:0], RdScheTopWrapper.U_RD_SCHE_TOP_SV.rddataCrsbarIn[_mbase_iDcpIn].Pld}),
								.din_vld_i(RdScheTopWrapper.U_RD_SCHE_TOP_SV.rddataCrsbarIn[_mbase_iDcpIn].Vld),
								.din_rdy_o(RdScheTopWrapper.U_RD_SCHE_TOP_SV.rddataCrsbarIn[_mbase_iDcpIn].Rdy),
								.dout_o({swiInDst, swiInPld}),
								.dout_vld_o(swiInVld),
								.dout_rdy_i(swiInRdy)
							);
							// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:39:3
							genvar _gv_i_3;
							// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:40:3
							for (_gv_i_3 = 0; _gv_i_3 < RNUM; _gv_i_3 = _gv_i_3 + 1) begin : GEN_ROUTE
								localparam i = _gv_i_3;
								// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:42:7
								always @(*) begin
									if (_sv2v_0)
										;
									// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:44:9
									if (swiInVld && (swiInDst[3-:4] == i))
										// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:45:11
										swiOutVld[i] = swiInVld;
									else
										// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:47:11
										swiOutVld[i] = 1'b0;
								end
							end
							// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:53:3
							reg signed [31:0] j;
							// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:54:3
							always @(*) begin
								if (_sv2v_0)
									;
								// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:55:5
								if (swiInVld) begin
									begin
										// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:56:7
										for (j = 0; j < RNUM; j = j + 1)
											begin
												// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:58:9
												if (swiInDst[3-:4] == j)
													// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:59:11
													swiInRdy = swiOutRdy[j];
											end
									end
								end
								else
									// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:63:7
									swiInRdy = 1'b0;
							end
							// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:67:3
							for (_gv_i_3 = 0; _gv_i_3 < RNUM; _gv_i_3 = _gv_i_3 + 1) begin : GEN_OUTBUF
								localparam i = _gv_i_3;
								// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:69:7
								gnrl_buf #(
									.DW(37),
									.CUT_RDY(1)
								) U_OUTBUF(
									.clk_i(iClk),
									.rst_n_i(iRst_n),
									.din_i({swiInDst, swiInPld}),
									.din_vld_i(swiOutVld[i]),
									.din_rdy_o(swiOutRdy[i]),
									.dout_o({RdScheTopWrapper.U_RD_SCHE_TOP_SV.U_RDDATA_CRSBAR.U_CRSBAR.xbarCon[i + _mbase_oDcpOut].Dst[3:0], RdScheTopWrapper.U_RD_SCHE_TOP_SV.U_RDDATA_CRSBAR.U_CRSBAR.xbarCon[i + _mbase_oDcpOut].Pld}),
									.dout_vld_o(RdScheTopWrapper.U_RD_SCHE_TOP_SV.U_RDDATA_CRSBAR.U_CRSBAR.xbarCon[i + _mbase_oDcpOut].Vld),
									.dout_rdy_i(RdScheTopWrapper.U_RD_SCHE_TOP_SV.U_RDDATA_CRSBAR.U_CRSBAR.xbarCon[i + _mbase_oDcpOut].Rdy)
								);
							end
							initial _sv2v_0 = 0;
						end
						assign U_ROUTEUNIT.iClk = iClk;
						assign U_ROUTEUNIT.iRst_n = iRst_n;
						// Trace: src/src/rtl/design/svsrc/DcpCrossbarNxN.sv:72:7
						// expanded module instance: U_SWITCHUNIT
						localparam _bbase_C87B5_iDcpIn = N * _gv_i_1;
						localparam _bbase_C87B5_oDcpOut = _gv_i_1 + _mbase_oDcpOut;
						localparam _param_C87B5_DW = DW;
						localparam _param_C87B5_AW = AW;
						localparam _param_C87B5_SNUM = N;
						if (1) begin : U_SWITCHUNIT
							// Trace: src/src/rtl/design/svsrc/DcpSwitchUnit.sv:28:13
							localparam DW = _param_C87B5_DW;
							// Trace: src/src/rtl/design/svsrc/DcpSwitchUnit.sv:29:13
							localparam AW = _param_C87B5_AW;
							// Trace: src/src/rtl/design/svsrc/DcpSwitchUnit.sv:30:13
							localparam SNUM = _param_C87B5_SNUM;
							// Trace: src/src/rtl/design/svsrc/DcpSwitchUnit.sv:32:3
							wire iClk;
							// Trace: src/src/rtl/design/svsrc/DcpSwitchUnit.sv:33:3
							wire iRst_n;
							// Trace: src/src/rtl/design/svsrc/DcpSwitchUnit.sv:35:3
							localparam _mbase_iDcpIn = _bbase_C87B5_iDcpIn;
							// Trace: src/src/rtl/design/svsrc/DcpSwitchUnit.sv:36:3
							localparam _mbase_oDcpOut = _bbase_C87B5_oDcpOut;
							// Trace: src/src/rtl/design/svsrc/DcpSwitchUnit.sv:38:3
							wire [15:0] arbInReqArray;
							// Trace: src/src/rtl/design/svsrc/DcpSwitchUnit.sv:39:3
							wire [15:0] arbInGntArray;
							// Trace: src/src/rtl/design/svsrc/DcpSwitchUnit.sv:40:3
							wire [591:0] arbInPldArray;
							// Trace: src/src/rtl/design/svsrc/DcpSwitchUnit.sv:42:3
							wire arbOutReq;
							// Trace: src/src/rtl/design/svsrc/DcpSwitchUnit.sv:43:3
							wire arbOutGnt;
							// Trace: src/src/rtl/design/svsrc/DcpSwitchUnit.sv:44:3
							wire [36:0] arbOutPld;
							// Trace: src/src/rtl/design/svsrc/DcpSwitchUnit.sv:46:3
							genvar _gv_i_4;
							// Trace: src/src/rtl/design/svsrc/DcpSwitchUnit.sv:48:3
							for (_gv_i_4 = 0; _gv_i_4 < SNUM; _gv_i_4 = _gv_i_4 + 1) begin : GEN_INBUF
								localparam i = _gv_i_4;
								// Trace: src/src/rtl/design/svsrc/DcpSwitchUnit.sv:50:7
								gnrl_buf #(
									.DW(37),
									.CUT_RDY(1)
								) U_INBUF(
									.clk_i(iClk),
									.rst_n_i(iRst_n),
									.din_i({RdScheTopWrapper.U_RD_SCHE_TOP_SV.U_RDDATA_CRSBAR.U_CRSBAR.xbarConT[i + _mbase_iDcpIn].Dst, RdScheTopWrapper.U_RD_SCHE_TOP_SV.U_RDDATA_CRSBAR.U_CRSBAR.xbarConT[i + _mbase_iDcpIn].Pld}),
									.din_vld_i(RdScheTopWrapper.U_RD_SCHE_TOP_SV.U_RDDATA_CRSBAR.U_CRSBAR.xbarConT[i + _mbase_iDcpIn].Vld),
									.din_rdy_o(RdScheTopWrapper.U_RD_SCHE_TOP_SV.U_RDDATA_CRSBAR.U_CRSBAR.xbarConT[i + _mbase_iDcpIn].Rdy),
									.dout_o(arbInPldArray[i * 37+:37]),
									.dout_vld_o(arbInReqArray[i]),
									.dout_rdy_i(arbInGntArray[i])
								);
							end
							// Trace: src/src/rtl/design/svsrc/DcpSwitchUnit.sv:67:3
							rr_arb_tree #(
								.NumIn(SNUM),
								.DataWidth(37),
								.AxiVldRdy(1),
								.LockIn(0)
							) U_RR_ARB(
								.rst_ni(iRst_n),
								.clk_i(iClk),
								.req_i(arbInReqArray),
								.gnt_o(arbInGntArray),
								.data_i(arbInPldArray),
								.req_o(arbOutReq),
								.gnt_i(arbOutGnt),
								.data_o(arbOutPld)
							);
							// Trace: src/src/rtl/design/svsrc/DcpSwitchUnit.sv:86:3
							gnrl_buf #(
								.DW(37),
								.CUT_RDY(1)
							) U_INBUF(
								.clk_i(iClk),
								.rst_n_i(iRst_n),
								.din_i(arbOutPld),
								.din_vld_i(arbOutReq),
								.din_rdy_o(arbOutGnt),
								.dout_o({RdScheTopWrapper.U_RD_SCHE_TOP_SV.rddataCrsbarOut[_mbase_oDcpOut].Dst, RdScheTopWrapper.U_RD_SCHE_TOP_SV.rddataCrsbarOut[_mbase_oDcpOut].Pld}),
								.dout_vld_o(RdScheTopWrapper.U_RD_SCHE_TOP_SV.rddataCrsbarOut[_mbase_oDcpOut].Vld),
								.dout_rdy_i(RdScheTopWrapper.U_RD_SCHE_TOP_SV.rddataCrsbarOut[_mbase_oDcpOut].Rdy)
							);
						end
						assign U_SWITCHUNIT.iClk = iClk;
						assign U_SWITCHUNIT.iRst_n = iRst_n;
					end
				end
				assign U_CRSBAR.iClk = iClk;
				assign U_CRSBAR.iRst_n = iRst_n;
			end
			assign U_RDDATA_CRSBAR.iClk = iClk;
			assign U_RDDATA_CRSBAR.iRst_n = iRst_n;
			// Trace: src/src/rtl/design/svsrc/RdScheTop.sv:72:3
			// expanded module instance: U_RDCMD_CRSBAR
			localparam _bbase_FAFE3_iRdCmdIn = 0;
			localparam _bbase_FAFE3_oRdCmdOut = 0;
			if (1) begin : U_RDCMD_CRSBAR
				// Trace: src/src/rtl/design/svsrc/DcpRdCmd16x16.sv:27:3
				wire iClk;
				// Trace: src/src/rtl/design/svsrc/DcpRdCmd16x16.sv:28:3
				wire iRst_n;
				// Trace: src/src/rtl/design/svsrc/DcpRdCmd16x16.sv:30:3
				localparam _mbase_iRdCmdIn = 0;
				// Trace: src/src/rtl/design/svsrc/DcpRdCmd16x16.sv:31:3
				localparam _mbase_oRdCmdOut = 0;
				// Trace: src/src/rtl/design/svsrc/DcpRdCmd16x16.sv:33:3
				localparam CRSBAR_N = 4;
				// Trace: src/src/rtl/design/svsrc/DcpRdCmd16x16.sv:34:3
				localparam CRSBAR_WIDTH = 21;
				// Trace: src/src/rtl/design/svsrc/DcpRdCmd16x16.sv:36:3
				// expanded interface instance: switchOut
				localparam _param_CF9F8_DW = CRSBAR_WIDTH;
				localparam _param_CF9F8_AW = 4;
				genvar _arr_CF9F8;
				for (_arr_CF9F8 = 0; _arr_CF9F8 <= 3; _arr_CF9F8 = _arr_CF9F8 + 1) begin : switchOut
					// Trace: src/src/rtl/design/svsrc/interface_list.sv:64:33
					localparam DW = _param_CF9F8_DW;
					// Trace: src/src/rtl/design/svsrc/interface_list.sv:64:52
					localparam AW = _param_CF9F8_AW;
					// Trace: src/src/rtl/design/svsrc/interface_list.sv:65:3
					wire [20:0] Pld;
					// Trace: src/src/rtl/design/svsrc/interface_list.sv:66:3
					wire [3:0] Dst;
					// Trace: src/src/rtl/design/svsrc/interface_list.sv:67:3
					wire Vld;
					// Trace: src/src/rtl/design/svsrc/interface_list.sv:68:3
					wire Rdy;
					// Trace: src/src/rtl/design/svsrc/interface_list.sv:69:3
					// Trace: src/src/rtl/design/svsrc/interface_list.sv:75:3
				end
				// Trace: src/src/rtl/design/svsrc/DcpRdCmd16x16.sv:37:3
				// expanded interface instance: routeIn
				localparam _param_37094_DW = CRSBAR_WIDTH;
				localparam _param_37094_AW = 4;
				genvar _arr_37094;
				for (_arr_37094 = 0; _arr_37094 <= 3; _arr_37094 = _arr_37094 + 1) begin : routeIn
					// Trace: src/src/rtl/design/svsrc/interface_list.sv:64:33
					localparam DW = _param_37094_DW;
					// Trace: src/src/rtl/design/svsrc/interface_list.sv:64:52
					localparam AW = _param_37094_AW;
					// Trace: src/src/rtl/design/svsrc/interface_list.sv:65:3
					wire [20:0] Pld;
					// Trace: src/src/rtl/design/svsrc/interface_list.sv:66:3
					wire [3:0] Dst;
					// Trace: src/src/rtl/design/svsrc/interface_list.sv:67:3
					wire Vld;
					// Trace: src/src/rtl/design/svsrc/interface_list.sv:68:3
					wire Rdy;
					// Trace: src/src/rtl/design/svsrc/interface_list.sv:69:3
					// Trace: src/src/rtl/design/svsrc/interface_list.sv:75:3
				end
				// Trace: src/src/rtl/design/svsrc/DcpRdCmd16x16.sv:39:3
				// expanded interface instance: rdCmdIn
				localparam _param_93D41_DW = CRSBAR_WIDTH;
				localparam _param_93D41_AW = 4;
				genvar _arr_93D41;
				for (_arr_93D41 = 0; _arr_93D41 <= 15; _arr_93D41 = _arr_93D41 + 1) begin : rdCmdIn
					// Trace: src/src/rtl/design/svsrc/interface_list.sv:64:33
					localparam DW = _param_93D41_DW;
					// Trace: src/src/rtl/design/svsrc/interface_list.sv:64:52
					localparam AW = _param_93D41_AW;
					// Trace: src/src/rtl/design/svsrc/interface_list.sv:65:3
					wire [20:0] Pld;
					// Trace: src/src/rtl/design/svsrc/interface_list.sv:66:3
					wire [3:0] Dst;
					// Trace: src/src/rtl/design/svsrc/interface_list.sv:67:3
					wire Vld;
					// Trace: src/src/rtl/design/svsrc/interface_list.sv:68:3
					wire Rdy;
					// Trace: src/src/rtl/design/svsrc/interface_list.sv:69:3
					// Trace: src/src/rtl/design/svsrc/interface_list.sv:75:3
				end
				// Trace: src/src/rtl/design/svsrc/DcpRdCmd16x16.sv:40:3
				// expanded interface instance: rdCmdOut
				localparam _param_35D97_DW = CRSBAR_WIDTH;
				localparam _param_35D97_AW = 4;
				genvar _arr_35D97;
				for (_arr_35D97 = 0; _arr_35D97 <= 15; _arr_35D97 = _arr_35D97 + 1) begin : rdCmdOut
					// Trace: src/src/rtl/design/svsrc/interface_list.sv:64:33
					localparam DW = _param_35D97_DW;
					// Trace: src/src/rtl/design/svsrc/interface_list.sv:64:52
					localparam AW = _param_35D97_AW;
					// Trace: src/src/rtl/design/svsrc/interface_list.sv:65:3
					wire [20:0] Pld;
					// Trace: src/src/rtl/design/svsrc/interface_list.sv:66:3
					wire [3:0] Dst;
					// Trace: src/src/rtl/design/svsrc/interface_list.sv:67:3
					wire Vld;
					// Trace: src/src/rtl/design/svsrc/interface_list.sv:68:3
					wire Rdy;
					// Trace: src/src/rtl/design/svsrc/interface_list.sv:69:3
					// Trace: src/src/rtl/design/svsrc/interface_list.sv:75:3
				end
				// Trace: src/src/rtl/design/svsrc/DcpRdCmd16x16.sv:42:3
				genvar _gv_i_2;
				// Trace: src/src/rtl/design/svsrc/DcpRdCmd16x16.sv:44:3
				for (_gv_i_2 = 0; _gv_i_2 < 4; _gv_i_2 = _gv_i_2 + 1) begin : GEN_INPUT_SWITCH
					localparam i = _gv_i_2;
					// Trace: src/src/rtl/design/svsrc/DcpRdCmd16x16.sv:46:7
					// expanded module instance: U_INPUT_SWITCH
					localparam _bbase_66B98_iDcpIn = 4 * _gv_i_2;
					localparam _bbase_66B98_oDcpOut = _gv_i_2;
					localparam _param_66B98_DW = CRSBAR_WIDTH;
					localparam _param_66B98_AW = 4;
					localparam _param_66B98_SNUM = 4;
					if (1) begin : U_INPUT_SWITCH
						// Trace: src/src/rtl/design/svsrc/DcpSwitchUnit.sv:28:13
						localparam DW = _param_66B98_DW;
						// Trace: src/src/rtl/design/svsrc/DcpSwitchUnit.sv:29:13
						localparam AW = _param_66B98_AW;
						// Trace: src/src/rtl/design/svsrc/DcpSwitchUnit.sv:30:13
						localparam SNUM = _param_66B98_SNUM;
						// Trace: src/src/rtl/design/svsrc/DcpSwitchUnit.sv:32:3
						wire iClk;
						// Trace: src/src/rtl/design/svsrc/DcpSwitchUnit.sv:33:3
						wire iRst_n;
						// Trace: src/src/rtl/design/svsrc/DcpSwitchUnit.sv:35:3
						localparam _mbase_iDcpIn = _bbase_66B98_iDcpIn;
						// Trace: src/src/rtl/design/svsrc/DcpSwitchUnit.sv:36:3
						localparam _mbase_oDcpOut = _bbase_66B98_oDcpOut;
						// Trace: src/src/rtl/design/svsrc/DcpSwitchUnit.sv:38:3
						wire [3:0] arbInReqArray;
						// Trace: src/src/rtl/design/svsrc/DcpSwitchUnit.sv:39:3
						wire [3:0] arbInGntArray;
						// Trace: src/src/rtl/design/svsrc/DcpSwitchUnit.sv:40:3
						wire [99:0] arbInPldArray;
						// Trace: src/src/rtl/design/svsrc/DcpSwitchUnit.sv:42:3
						wire arbOutReq;
						// Trace: src/src/rtl/design/svsrc/DcpSwitchUnit.sv:43:3
						wire arbOutGnt;
						// Trace: src/src/rtl/design/svsrc/DcpSwitchUnit.sv:44:3
						wire [24:0] arbOutPld;
						// Trace: src/src/rtl/design/svsrc/DcpSwitchUnit.sv:46:3
						genvar _gv_i_4;
						// Trace: src/src/rtl/design/svsrc/DcpSwitchUnit.sv:48:3
						for (_gv_i_4 = 0; _gv_i_4 < SNUM; _gv_i_4 = _gv_i_4 + 1) begin : GEN_INBUF
							localparam i = _gv_i_4;
							// Trace: src/src/rtl/design/svsrc/DcpSwitchUnit.sv:50:7
							gnrl_buf #(
								.DW(25),
								.CUT_RDY(1)
							) U_INBUF(
								.clk_i(iClk),
								.rst_n_i(iRst_n),
								.din_i({RdScheTopWrapper.U_RD_SCHE_TOP_SV.U_RDCMD_CRSBAR.rdCmdIn[i + _mbase_iDcpIn].Dst, RdScheTopWrapper.U_RD_SCHE_TOP_SV.U_RDCMD_CRSBAR.rdCmdIn[i + _mbase_iDcpIn].Pld}),
								.din_vld_i(RdScheTopWrapper.U_RD_SCHE_TOP_SV.U_RDCMD_CRSBAR.rdCmdIn[i + _mbase_iDcpIn].Vld),
								.din_rdy_o(RdScheTopWrapper.U_RD_SCHE_TOP_SV.U_RDCMD_CRSBAR.rdCmdIn[i + _mbase_iDcpIn].Rdy),
								.dout_o(arbInPldArray[i * 25+:25]),
								.dout_vld_o(arbInReqArray[i]),
								.dout_rdy_i(arbInGntArray[i])
							);
						end
						// Trace: src/src/rtl/design/svsrc/DcpSwitchUnit.sv:67:3
						rr_arb_tree #(
							.NumIn(SNUM),
							.DataWidth(25),
							.AxiVldRdy(1),
							.LockIn(0)
						) U_RR_ARB(
							.rst_ni(iRst_n),
							.clk_i(iClk),
							.req_i(arbInReqArray),
							.gnt_o(arbInGntArray),
							.data_i(arbInPldArray),
							.req_o(arbOutReq),
							.gnt_i(arbOutGnt),
							.data_o(arbOutPld)
						);
						// Trace: src/src/rtl/design/svsrc/DcpSwitchUnit.sv:86:3
						gnrl_buf #(
							.DW(25),
							.CUT_RDY(1)
						) U_INBUF(
							.clk_i(iClk),
							.rst_n_i(iRst_n),
							.din_i(arbOutPld),
							.din_vld_i(arbOutReq),
							.din_rdy_o(arbOutGnt),
							.dout_o({RdScheTopWrapper.U_RD_SCHE_TOP_SV.U_RDCMD_CRSBAR.switchOut[_mbase_oDcpOut].Dst, RdScheTopWrapper.U_RD_SCHE_TOP_SV.U_RDCMD_CRSBAR.switchOut[_mbase_oDcpOut].Pld}),
							.dout_vld_o(RdScheTopWrapper.U_RD_SCHE_TOP_SV.U_RDCMD_CRSBAR.switchOut[_mbase_oDcpOut].Vld),
							.dout_rdy_i(RdScheTopWrapper.U_RD_SCHE_TOP_SV.U_RDCMD_CRSBAR.switchOut[_mbase_oDcpOut].Rdy)
						);
					end
					assign U_INPUT_SWITCH.iClk = iClk;
					assign U_INPUT_SWITCH.iRst_n = iRst_n;
				end
				// Trace: src/src/rtl/design/svsrc/DcpRdCmd16x16.sv:59:3
				// expanded module instance: U_CRSBAR
				localparam _bbase_509DC_iDcpIn = 0;
				localparam _bbase_509DC_oDcpOut = 0;
				localparam _param_509DC_DW = CRSBAR_WIDTH;
				localparam _param_509DC_AW = 4;
				localparam _param_509DC_N = 4;
				if (1) begin : U_CRSBAR
					// Trace: src/src/rtl/design/svsrc/DcpCrossbarNxN.sv:26:13
					localparam DW = _param_509DC_DW;
					// Trace: src/src/rtl/design/svsrc/DcpCrossbarNxN.sv:27:13
					localparam AW = _param_509DC_AW;
					// Trace: src/src/rtl/design/svsrc/DcpCrossbarNxN.sv:28:13
					localparam N = _param_509DC_N;
					// Trace: src/src/rtl/design/svsrc/DcpCrossbarNxN.sv:30:3
					wire iClk;
					// Trace: src/src/rtl/design/svsrc/DcpCrossbarNxN.sv:31:3
					wire iRst_n;
					// Trace: src/src/rtl/design/svsrc/DcpCrossbarNxN.sv:32:3
					localparam _mbase_iDcpIn = 0;
					// Trace: src/src/rtl/design/svsrc/DcpCrossbarNxN.sv:33:3
					localparam _mbase_oDcpOut = 0;
					// Trace: src/src/rtl/design/svsrc/DcpCrossbarNxN.sv:35:3
					// Trace: src/src/rtl/design/svsrc/DcpCrossbarNxN.sv:41:3
					// expanded interface instance: xbarCon
					localparam _param_7FFE1_DW = DW;
					localparam _param_7FFE1_AW = AW;
					genvar _arr_7FFE1;
					for (_arr_7FFE1 = 0; _arr_7FFE1 <= 15; _arr_7FFE1 = _arr_7FFE1 + 1) begin : xbarCon
						// Trace: src/src/rtl/design/svsrc/interface_list.sv:64:33
						localparam DW = _param_7FFE1_DW;
						// Trace: src/src/rtl/design/svsrc/interface_list.sv:64:52
						localparam AW = _param_7FFE1_AW;
						// Trace: src/src/rtl/design/svsrc/interface_list.sv:65:3
						wire [20:0] Pld;
						// Trace: src/src/rtl/design/svsrc/interface_list.sv:66:3
						wire [3:0] Dst;
						// Trace: src/src/rtl/design/svsrc/interface_list.sv:67:3
						wire Vld;
						// Trace: src/src/rtl/design/svsrc/interface_list.sv:68:3
						wire Rdy;
						// Trace: src/src/rtl/design/svsrc/interface_list.sv:69:3
						// Trace: src/src/rtl/design/svsrc/interface_list.sv:75:3
					end
					// Trace: src/src/rtl/design/svsrc/DcpCrossbarNxN.sv:42:3
					// expanded interface instance: xbarConT
					localparam _param_46BCA_DW = DW;
					localparam _param_46BCA_AW = AW;
					genvar _arr_46BCA;
					for (_arr_46BCA = 0; _arr_46BCA <= 15; _arr_46BCA = _arr_46BCA + 1) begin : xbarConT
						// Trace: src/src/rtl/design/svsrc/interface_list.sv:64:33
						localparam DW = _param_46BCA_DW;
						// Trace: src/src/rtl/design/svsrc/interface_list.sv:64:52
						localparam AW = _param_46BCA_AW;
						// Trace: src/src/rtl/design/svsrc/interface_list.sv:65:3
						wire [20:0] Pld;
						// Trace: src/src/rtl/design/svsrc/interface_list.sv:66:3
						wire [3:0] Dst;
						// Trace: src/src/rtl/design/svsrc/interface_list.sv:67:3
						wire Vld;
						// Trace: src/src/rtl/design/svsrc/interface_list.sv:68:3
						wire Rdy;
						// Trace: src/src/rtl/design/svsrc/interface_list.sv:69:3
						// Trace: src/src/rtl/design/svsrc/interface_list.sv:75:3
					end
					// Trace: src/src/rtl/design/svsrc/DcpCrossbarNxN.sv:44:3
					genvar _gv_i_1;
					// Trace: src/src/rtl/design/svsrc/DcpCrossbarNxN.sv:45:3
					genvar _gv_j_1;
					// Trace: src/src/rtl/design/svsrc/DcpCrossbarNxN.sv:46:3
					for (_gv_i_1 = 0; _gv_i_1 < N; _gv_i_1 = _gv_i_1 + 1) begin : GEN_XBAR_CON_TRANS_ROW
						localparam i = _gv_i_1;
						for (_gv_j_1 = 0; _gv_j_1 < N; _gv_j_1 = _gv_j_1 + 1) begin : GEN_XBAR_CON_TRANS_COL
							localparam j = _gv_j_1;
							// Trace: src/src/rtl/design/svsrc/DcpCrossbarNxN.sv:52:9
							assign xbarConT[(i * N) + j].Vld = xbarCon[(j * N) + i].Vld;
							// Trace: src/src/rtl/design/svsrc/DcpCrossbarNxN.sv:53:9
							assign xbarConT[(i * N) + j].Pld = xbarCon[(j * N) + i].Pld;
							// Trace: src/src/rtl/design/svsrc/DcpCrossbarNxN.sv:54:9
							assign xbarConT[(i * N) + j].Dst = xbarCon[(j * N) + i].Dst;
							// Trace: src/src/rtl/design/svsrc/DcpCrossbarNxN.sv:55:9
							assign xbarCon[(j * N) + i].Rdy = xbarConT[(i * N) + j].Rdy;
						end
					end
					// Trace: src/src/rtl/design/svsrc/DcpCrossbarNxN.sv:60:3
					for (_gv_i_1 = 0; _gv_i_1 < N; _gv_i_1 = _gv_i_1 + 1) begin : GEN_CON
						localparam i = _gv_i_1;
						// Trace: src/src/rtl/design/svsrc/DcpCrossbarNxN.sv:62:7
						// expanded module instance: U_ROUTEUNIT
						localparam _bbase_08BCB_iDcpIn = _gv_i_1 + _mbase_iDcpIn;
						localparam _bbase_08BCB_oDcpOut = N * _gv_i_1;
						localparam _param_08BCB_DW = DW;
						localparam _param_08BCB_AW = AW;
						localparam _param_08BCB_RNUM = N;
						if (1) begin : U_ROUTEUNIT
							reg _sv2v_0;
							// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:3:13
							localparam DW = _param_08BCB_DW;
							// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:4:13
							localparam AW = _param_08BCB_AW;
							// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:5:13
							localparam RNUM = _param_08BCB_RNUM;
							// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:7:3
							wire iClk;
							// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:8:3
							wire iRst_n;
							// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:10:3
							localparam _mbase_iDcpIn = _bbase_08BCB_iDcpIn;
							// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:11:3
							localparam _mbase_oDcpOut = _bbase_08BCB_oDcpOut;
							// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:14:3
							reg swiInRdy;
							// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:15:3
							wire swiInVld;
							// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:16:3
							wire [20:0] swiInPld;
							// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:17:3
							wire [3:0] swiInDst;
							// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:19:3
							reg [3:0] swiOutVld;
							// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:20:3
							wire [3:0] swiOutRdy;
							// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:22:3
							localparam IDLE = 1'b0;
							// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:23:3
							localparam GRANT = 1'b1;
							// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:25:3
							gnrl_buf #(
								.DW(25),
								.CUT_RDY(1)
							) U_INBUF(
								.clk_i(iClk),
								.rst_n_i(iRst_n),
								.din_i({RdScheTopWrapper.U_RD_SCHE_TOP_SV.U_RDCMD_CRSBAR.switchOut[_mbase_iDcpIn].Dst[3:0], RdScheTopWrapper.U_RD_SCHE_TOP_SV.U_RDCMD_CRSBAR.switchOut[_mbase_iDcpIn].Pld}),
								.din_vld_i(RdScheTopWrapper.U_RD_SCHE_TOP_SV.U_RDCMD_CRSBAR.switchOut[_mbase_iDcpIn].Vld),
								.din_rdy_o(RdScheTopWrapper.U_RD_SCHE_TOP_SV.U_RDCMD_CRSBAR.switchOut[_mbase_iDcpIn].Rdy),
								.dout_o({swiInDst, swiInPld}),
								.dout_vld_o(swiInVld),
								.dout_rdy_i(swiInRdy)
							);
							// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:39:3
							genvar _gv_i_3;
							// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:40:3
							for (_gv_i_3 = 0; _gv_i_3 < RNUM; _gv_i_3 = _gv_i_3 + 1) begin : GEN_ROUTE
								localparam i = _gv_i_3;
								// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:42:7
								always @(*) begin
									if (_sv2v_0)
										;
									// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:44:9
									if (swiInVld && (swiInDst[3-:2] == i))
										// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:45:11
										swiOutVld[i] = swiInVld;
									else
										// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:47:11
										swiOutVld[i] = 1'b0;
								end
							end
							// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:53:3
							reg signed [31:0] j;
							// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:54:3
							always @(*) begin
								if (_sv2v_0)
									;
								// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:55:5
								if (swiInVld) begin
									begin
										// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:56:7
										for (j = 0; j < RNUM; j = j + 1)
											begin
												// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:58:9
												if (swiInDst[3-:2] == j)
													// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:59:11
													swiInRdy = swiOutRdy[j];
											end
									end
								end
								else
									// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:63:7
									swiInRdy = 1'b0;
							end
							// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:67:3
							for (_gv_i_3 = 0; _gv_i_3 < RNUM; _gv_i_3 = _gv_i_3 + 1) begin : GEN_OUTBUF
								localparam i = _gv_i_3;
								// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:69:7
								gnrl_buf #(
									.DW(25),
									.CUT_RDY(1)
								) U_OUTBUF(
									.clk_i(iClk),
									.rst_n_i(iRst_n),
									.din_i({swiInDst, swiInPld}),
									.din_vld_i(swiOutVld[i]),
									.din_rdy_o(swiOutRdy[i]),
									.dout_o({RdScheTopWrapper.U_RD_SCHE_TOP_SV.U_RDCMD_CRSBAR.U_CRSBAR.xbarCon[i + _mbase_oDcpOut].Dst[3:0], RdScheTopWrapper.U_RD_SCHE_TOP_SV.U_RDCMD_CRSBAR.U_CRSBAR.xbarCon[i + _mbase_oDcpOut].Pld}),
									.dout_vld_o(RdScheTopWrapper.U_RD_SCHE_TOP_SV.U_RDCMD_CRSBAR.U_CRSBAR.xbarCon[i + _mbase_oDcpOut].Vld),
									.dout_rdy_i(RdScheTopWrapper.U_RD_SCHE_TOP_SV.U_RDCMD_CRSBAR.U_CRSBAR.xbarCon[i + _mbase_oDcpOut].Rdy)
								);
							end
							initial _sv2v_0 = 0;
						end
						assign U_ROUTEUNIT.iClk = iClk;
						assign U_ROUTEUNIT.iRst_n = iRst_n;
						// Trace: src/src/rtl/design/svsrc/DcpCrossbarNxN.sv:72:7
						// expanded module instance: U_SWITCHUNIT
						localparam _bbase_C87B5_iDcpIn = N * _gv_i_1;
						localparam _bbase_C87B5_oDcpOut = _gv_i_1 + _mbase_oDcpOut;
						localparam _param_C87B5_DW = DW;
						localparam _param_C87B5_AW = AW;
						localparam _param_C87B5_SNUM = N;
						if (1) begin : U_SWITCHUNIT
							// Trace: src/src/rtl/design/svsrc/DcpSwitchUnit.sv:28:13
							localparam DW = _param_C87B5_DW;
							// Trace: src/src/rtl/design/svsrc/DcpSwitchUnit.sv:29:13
							localparam AW = _param_C87B5_AW;
							// Trace: src/src/rtl/design/svsrc/DcpSwitchUnit.sv:30:13
							localparam SNUM = _param_C87B5_SNUM;
							// Trace: src/src/rtl/design/svsrc/DcpSwitchUnit.sv:32:3
							wire iClk;
							// Trace: src/src/rtl/design/svsrc/DcpSwitchUnit.sv:33:3
							wire iRst_n;
							// Trace: src/src/rtl/design/svsrc/DcpSwitchUnit.sv:35:3
							localparam _mbase_iDcpIn = _bbase_C87B5_iDcpIn;
							// Trace: src/src/rtl/design/svsrc/DcpSwitchUnit.sv:36:3
							localparam _mbase_oDcpOut = _bbase_C87B5_oDcpOut;
							// Trace: src/src/rtl/design/svsrc/DcpSwitchUnit.sv:38:3
							wire [3:0] arbInReqArray;
							// Trace: src/src/rtl/design/svsrc/DcpSwitchUnit.sv:39:3
							wire [3:0] arbInGntArray;
							// Trace: src/src/rtl/design/svsrc/DcpSwitchUnit.sv:40:3
							wire [99:0] arbInPldArray;
							// Trace: src/src/rtl/design/svsrc/DcpSwitchUnit.sv:42:3
							wire arbOutReq;
							// Trace: src/src/rtl/design/svsrc/DcpSwitchUnit.sv:43:3
							wire arbOutGnt;
							// Trace: src/src/rtl/design/svsrc/DcpSwitchUnit.sv:44:3
							wire [24:0] arbOutPld;
							// Trace: src/src/rtl/design/svsrc/DcpSwitchUnit.sv:46:3
							genvar _gv_i_4;
							// Trace: src/src/rtl/design/svsrc/DcpSwitchUnit.sv:48:3
							for (_gv_i_4 = 0; _gv_i_4 < SNUM; _gv_i_4 = _gv_i_4 + 1) begin : GEN_INBUF
								localparam i = _gv_i_4;
								// Trace: src/src/rtl/design/svsrc/DcpSwitchUnit.sv:50:7
								gnrl_buf #(
									.DW(25),
									.CUT_RDY(1)
								) U_INBUF(
									.clk_i(iClk),
									.rst_n_i(iRst_n),
									.din_i({RdScheTopWrapper.U_RD_SCHE_TOP_SV.U_RDCMD_CRSBAR.U_CRSBAR.xbarConT[i + _mbase_iDcpIn].Dst, RdScheTopWrapper.U_RD_SCHE_TOP_SV.U_RDCMD_CRSBAR.U_CRSBAR.xbarConT[i + _mbase_iDcpIn].Pld}),
									.din_vld_i(RdScheTopWrapper.U_RD_SCHE_TOP_SV.U_RDCMD_CRSBAR.U_CRSBAR.xbarConT[i + _mbase_iDcpIn].Vld),
									.din_rdy_o(RdScheTopWrapper.U_RD_SCHE_TOP_SV.U_RDCMD_CRSBAR.U_CRSBAR.xbarConT[i + _mbase_iDcpIn].Rdy),
									.dout_o(arbInPldArray[i * 25+:25]),
									.dout_vld_o(arbInReqArray[i]),
									.dout_rdy_i(arbInGntArray[i])
								);
							end
							// Trace: src/src/rtl/design/svsrc/DcpSwitchUnit.sv:67:3
							rr_arb_tree #(
								.NumIn(SNUM),
								.DataWidth(25),
								.AxiVldRdy(1),
								.LockIn(0)
							) U_RR_ARB(
								.rst_ni(iRst_n),
								.clk_i(iClk),
								.req_i(arbInReqArray),
								.gnt_o(arbInGntArray),
								.data_i(arbInPldArray),
								.req_o(arbOutReq),
								.gnt_i(arbOutGnt),
								.data_o(arbOutPld)
							);
							// Trace: src/src/rtl/design/svsrc/DcpSwitchUnit.sv:86:3
							gnrl_buf #(
								.DW(25),
								.CUT_RDY(1)
							) U_INBUF(
								.clk_i(iClk),
								.rst_n_i(iRst_n),
								.din_i(arbOutPld),
								.din_vld_i(arbOutReq),
								.din_rdy_o(arbOutGnt),
								.dout_o({RdScheTopWrapper.U_RD_SCHE_TOP_SV.U_RDCMD_CRSBAR.routeIn[_mbase_oDcpOut].Dst, RdScheTopWrapper.U_RD_SCHE_TOP_SV.U_RDCMD_CRSBAR.routeIn[_mbase_oDcpOut].Pld}),
								.dout_vld_o(RdScheTopWrapper.U_RD_SCHE_TOP_SV.U_RDCMD_CRSBAR.routeIn[_mbase_oDcpOut].Vld),
								.dout_rdy_i(RdScheTopWrapper.U_RD_SCHE_TOP_SV.U_RDCMD_CRSBAR.routeIn[_mbase_oDcpOut].Rdy)
							);
						end
						assign U_SWITCHUNIT.iClk = iClk;
						assign U_SWITCHUNIT.iRst_n = iRst_n;
					end
				end
				assign U_CRSBAR.iClk = iClk;
				assign U_CRSBAR.iRst_n = iRst_n;
				// Trace: src/src/rtl/design/svsrc/DcpRdCmd16x16.sv:70:3
				for (_gv_i_2 = 0; _gv_i_2 < 4; _gv_i_2 = _gv_i_2 + 1) begin : GEN_OUTPUT_ROUTE
					localparam i = _gv_i_2;
					// Trace: src/src/rtl/design/svsrc/DcpRdCmd16x16.sv:72:7
					// expanded module instance: U_OUTPUT_ROUTE
					localparam _bbase_37972_iDcpIn = _gv_i_2;
					localparam _bbase_37972_oDcpOut = _gv_i_2 * 4;
					localparam _param_37972_DW = CRSBAR_WIDTH;
					localparam _param_37972_AW = 2;
					localparam _param_37972_RNUM = 4;
					if (1) begin : U_OUTPUT_ROUTE
						reg _sv2v_0;
						// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:3:13
						localparam DW = _param_37972_DW;
						// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:4:13
						localparam AW = _param_37972_AW;
						// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:5:13
						localparam RNUM = _param_37972_RNUM;
						// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:7:3
						wire iClk;
						// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:8:3
						wire iRst_n;
						// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:10:3
						localparam _mbase_iDcpIn = _bbase_37972_iDcpIn;
						// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:11:3
						localparam _mbase_oDcpOut = _bbase_37972_oDcpOut;
						// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:14:3
						reg swiInRdy;
						// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:15:3
						wire swiInVld;
						// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:16:3
						wire [20:0] swiInPld;
						// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:17:3
						wire [1:0] swiInDst;
						// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:19:3
						reg [3:0] swiOutVld;
						// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:20:3
						wire [3:0] swiOutRdy;
						// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:22:3
						localparam IDLE = 1'b0;
						// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:23:3
						localparam GRANT = 1'b1;
						// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:25:3
						gnrl_buf #(
							.DW(23),
							.CUT_RDY(1)
						) U_INBUF(
							.clk_i(iClk),
							.rst_n_i(iRst_n),
							.din_i({RdScheTopWrapper.U_RD_SCHE_TOP_SV.U_RDCMD_CRSBAR.routeIn[_mbase_iDcpIn].Dst[1:0], RdScheTopWrapper.U_RD_SCHE_TOP_SV.U_RDCMD_CRSBAR.routeIn[_mbase_iDcpIn].Pld}),
							.din_vld_i(RdScheTopWrapper.U_RD_SCHE_TOP_SV.U_RDCMD_CRSBAR.routeIn[_mbase_iDcpIn].Vld),
							.din_rdy_o(RdScheTopWrapper.U_RD_SCHE_TOP_SV.U_RDCMD_CRSBAR.routeIn[_mbase_iDcpIn].Rdy),
							.dout_o({swiInDst, swiInPld}),
							.dout_vld_o(swiInVld),
							.dout_rdy_i(swiInRdy)
						);
						// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:39:3
						genvar _gv_i_3;
						// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:40:3
						for (_gv_i_3 = 0; _gv_i_3 < RNUM; _gv_i_3 = _gv_i_3 + 1) begin : GEN_ROUTE
							localparam i = _gv_i_3;
							// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:42:7
							always @(*) begin
								if (_sv2v_0)
									;
								// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:44:9
								if (swiInVld && (swiInDst[1-:2] == i))
									// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:45:11
									swiOutVld[i] = swiInVld;
								else
									// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:47:11
									swiOutVld[i] = 1'b0;
							end
						end
						// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:53:3
						reg signed [31:0] j;
						// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:54:3
						always @(*) begin
							if (_sv2v_0)
								;
							// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:55:5
							if (swiInVld) begin
								begin
									// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:56:7
									for (j = 0; j < RNUM; j = j + 1)
										begin
											// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:58:9
											if (swiInDst[1-:2] == j)
												// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:59:11
												swiInRdy = swiOutRdy[j];
										end
								end
							end
							else
								// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:63:7
								swiInRdy = 1'b0;
						end
						// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:67:3
						for (_gv_i_3 = 0; _gv_i_3 < RNUM; _gv_i_3 = _gv_i_3 + 1) begin : GEN_OUTBUF
							localparam i = _gv_i_3;
							// Trace: src/src/rtl/design/svsrc/DcpRouteUnit.sv:69:7
							gnrl_buf #(
								.DW(23),
								.CUT_RDY(1)
							) U_OUTBUF(
								.clk_i(iClk),
								.rst_n_i(iRst_n),
								.din_i({swiInDst, swiInPld}),
								.din_vld_i(swiOutVld[i]),
								.din_rdy_o(swiOutRdy[i]),
								.dout_o({RdScheTopWrapper.U_RD_SCHE_TOP_SV.U_RDCMD_CRSBAR.rdCmdOut[i + _mbase_oDcpOut].Dst[1:0], RdScheTopWrapper.U_RD_SCHE_TOP_SV.U_RDCMD_CRSBAR.rdCmdOut[i + _mbase_oDcpOut].Pld}),
								.dout_vld_o(RdScheTopWrapper.U_RD_SCHE_TOP_SV.U_RDCMD_CRSBAR.rdCmdOut[i + _mbase_oDcpOut].Vld),
								.dout_rdy_i(RdScheTopWrapper.U_RD_SCHE_TOP_SV.U_RDCMD_CRSBAR.rdCmdOut[i + _mbase_oDcpOut].Rdy)
							);
						end
						initial _sv2v_0 = 0;
					end
					assign U_OUTPUT_ROUTE.iClk = iClk;
					assign U_OUTPUT_ROUTE.iRst_n = iRst_n;
				end
				// Trace: src/src/rtl/design/svsrc/DcpRdCmd16x16.sv:86:3
				for (_gv_i_2 = 0; _gv_i_2 < 16; _gv_i_2 = _gv_i_2 + 1) begin : GENCON
					localparam i = _gv_i_2;
					// Trace: src/src/rtl/design/svsrc/DcpRdCmd16x16.sv:88:7
					assign rdCmdOut[i].Rdy = RdScheTopWrapper.U_RD_SCHE_TOP_SV.rdcmdCrsbarOut[i + _mbase_oRdCmdOut].Rdy;
					// Trace: src/src/rtl/design/svsrc/DcpRdCmd16x16.sv:89:7
					assign RdScheTopWrapper.U_RD_SCHE_TOP_SV.rdcmdCrsbarOut[i + _mbase_oRdCmdOut].Pld = rdCmdOut[i].Pld;
					// Trace: src/src/rtl/design/svsrc/DcpRdCmd16x16.sv:90:7
					assign RdScheTopWrapper.U_RD_SCHE_TOP_SV.rdcmdCrsbarOut[i + _mbase_oRdCmdOut].Vld = rdCmdOut[i].Vld;
					// Trace: src/src/rtl/design/svsrc/DcpRdCmd16x16.sv:91:7
					assign RdScheTopWrapper.U_RD_SCHE_TOP_SV.rdcmdCrsbarOut[i + _mbase_oRdCmdOut].Dst = rdCmdOut[i].Dst;
					// Trace: src/src/rtl/design/svsrc/DcpRdCmd16x16.sv:93:7
					assign RdScheTopWrapper.U_RD_SCHE_TOP_SV.rdcmdCrsbarIn[i + _mbase_iRdCmdIn].Rdy = rdCmdIn[i].Rdy;
					// Trace: src/src/rtl/design/svsrc/DcpRdCmd16x16.sv:94:7
					assign rdCmdIn[i].Pld = RdScheTopWrapper.U_RD_SCHE_TOP_SV.rdcmdCrsbarIn[i + _mbase_iRdCmdIn].Pld;
					// Trace: src/src/rtl/design/svsrc/DcpRdCmd16x16.sv:95:7
					assign rdCmdIn[i].Vld = RdScheTopWrapper.U_RD_SCHE_TOP_SV.rdcmdCrsbarIn[i + _mbase_iRdCmdIn].Vld;
					// Trace: src/src/rtl/design/svsrc/DcpRdCmd16x16.sv:96:7
					assign rdCmdIn[i].Dst = RdScheTopWrapper.U_RD_SCHE_TOP_SV.rdcmdCrsbarIn[i + _mbase_iRdCmdIn].Dst;
				end
			end
			assign U_RDCMD_CRSBAR.iClk = iClk;
			assign U_RDCMD_CRSBAR.iRst_n = iRst_n;
			// Trace: src/src/rtl/design/svsrc/RdScheTop.sv:80:3
			// expanded module instance: U_RDCTRLTOP16
			localparam _bbase_9AC28_iTagIn = 0;
			localparam _bbase_9AC28_oRdCmd = 0;
			localparam _bbase_9AC28_iRdData = 0;
			localparam _param_9AC28_PRI_DEPTH = PRI_DEPTH;
			localparam _param_9AC28_WRR_WEIGHT_NUM = WRR_WEIGHT_NUM;
			if (1) begin : U_RDCTRLTOP16
				// Trace: src/src/rtl/design/svsrc/RdCtrlTop16Ch.sv:26:13
				localparam PRI_DEPTH = _param_9AC28_PRI_DEPTH;
				// Trace: src/src/rtl/design/svsrc/RdCtrlTop16Ch.sv:28:13
				localparam PRI_NUM = 8;
				// Trace: src/src/rtl/design/svsrc/RdCtrlTop16Ch.sv:29:13
				localparam WRR_WEIGHT_NUM = _param_9AC28_WRR_WEIGHT_NUM;
				// Trace: src/src/rtl/design/svsrc/RdCtrlTop16Ch.sv:31:3
				wire iClk;
				// Trace: src/src/rtl/design/svsrc/RdCtrlTop16Ch.sv:32:3
				wire iRst_n;
				// Trace: src/src/rtl/design/svsrc/RdCtrlTop16Ch.sv:34:3
				localparam _mbase_iTagIn = 0;
				// Trace: src/src/rtl/design/svsrc/RdCtrlTop16Ch.sv:35:3
				localparam _mbase_oRdCmd = 0;
				// Trace: src/src/rtl/design/svsrc/RdCtrlTop16Ch.sv:37:3
				localparam _mbase_iRdData = 0;
				// Trace: src/src/rtl/design/svsrc/RdCtrlTop16Ch.sv:39:3
				wire [0:15] oRdSop;
				// Trace: src/src/rtl/design/svsrc/RdCtrlTop16Ch.sv:40:3
				wire [0:15] oRdEop;
				// Trace: src/src/rtl/design/svsrc/RdCtrlTop16Ch.sv:41:3
				wire [0:15] oRdVld;
				// Trace: src/src/rtl/design/svsrc/RdCtrlTop16Ch.sv:42:3
				wire [511:0] oRdData;
				// Trace: src/src/rtl/design/svsrc/RdCtrlTop16Ch.sv:43:3
				wire [0:15] iRdRdy;
				// Trace: src/src/rtl/design/svsrc/RdCtrlTop16Ch.sv:44:3
				wire [0:15] oRdLast;
				// Trace: src/src/rtl/design/svsrc/RdCtrlTop16Ch.sv:46:3
				wire [($clog2(WRR_WEIGHT_NUM) >= 0 ? (8 * ($clog2(WRR_WEIGHT_NUM) + 1)) - 1 : (8 * (1 - $clog2(WRR_WEIGHT_NUM))) + ($clog2(WRR_WEIGHT_NUM) - 1)):($clog2(WRR_WEIGHT_NUM) >= 0 ? 0 : $clog2(WRR_WEIGHT_NUM) + 0)] iWeightPld;
				// Trace: src/src/rtl/design/svsrc/RdCtrlTop16Ch.sv:47:3
				wire [3:0] iWeightIdx;
				// Trace: src/src/rtl/design/svsrc/RdCtrlTop16Ch.sv:48:3
				wire iWeightLoad;
				// Trace: src/src/rtl/design/svsrc/RdCtrlTop16Ch.sv:50:3
				genvar _gv_i_7;
				// Trace: src/src/rtl/design/svsrc/RdCtrlTop16Ch.sv:52:3
				wire [15:0] weightLoadArray;
				// Trace: src/src/rtl/design/svsrc/RdCtrlTop16Ch.sv:54:3
				for (_gv_i_7 = 0; _gv_i_7 < 16; _gv_i_7 = _gv_i_7 + 1) begin : genblk1
					localparam i = _gv_i_7;
					// Trace: src/src/rtl/design/svsrc/RdCtrlTop16Ch.sv:56:7
					assign weightLoadArray[i] = (iWeightIdx == i ? iWeightLoad : 1'b0);
					// Trace: src/src/rtl/design/svsrc/RdCtrlTop16Ch.sv:57:7
					// expanded module instance: U_RD_CHN
					localparam _bbase_177AB_iTagIn = _gv_i_7 + _mbase_iTagIn;
					localparam _bbase_177AB_oRdCmd = _gv_i_7 + _mbase_oRdCmd;
					localparam _bbase_177AB_iRdData = _gv_i_7 + _mbase_iRdData;
					localparam _param_177AB_PORT_ADDR = i;
					localparam _param_177AB_PRI_DEPTH = PRI_DEPTH;
					localparam _param_177AB_WRR_WEIGHT_NUM = WRR_WEIGHT_NUM;
					if (1) begin : U_RD_CHN
						// Trace: src/src/rtl/design/svsrc/RdCtrlTop1Ch.sv:26:13
						localparam PORT_ADDR = _param_177AB_PORT_ADDR;
						// Trace: src/src/rtl/design/svsrc/RdCtrlTop1Ch.sv:27:13
						localparam PRI_DEPTH = _param_177AB_PRI_DEPTH;
						// Trace: src/src/rtl/design/svsrc/RdCtrlTop1Ch.sv:29:13
						localparam PRI_NUM = 8;
						// Trace: src/src/rtl/design/svsrc/RdCtrlTop1Ch.sv:30:13
						localparam WRR_WEIGHT_NUM = _param_177AB_WRR_WEIGHT_NUM;
						// Trace: src/src/rtl/design/svsrc/RdCtrlTop1Ch.sv:33:3
						wire iClk;
						// Trace: src/src/rtl/design/svsrc/RdCtrlTop1Ch.sv:34:3
						wire iRst_n;
						// Trace: src/src/rtl/design/svsrc/RdCtrlTop1Ch.sv:36:3
						localparam _mbase_iTagIn = _bbase_177AB_iTagIn;
						// Trace: src/src/rtl/design/svsrc/RdCtrlTop1Ch.sv:37:3
						localparam _mbase_oRdCmd = _bbase_177AB_oRdCmd;
						// Trace: src/src/rtl/design/svsrc/RdCtrlTop1Ch.sv:39:3
						localparam _mbase_iRdData = _bbase_177AB_iRdData;
						// Trace: src/src/rtl/design/svsrc/RdCtrlTop1Ch.sv:41:3
						wire oRdSop;
						// Trace: src/src/rtl/design/svsrc/RdCtrlTop1Ch.sv:42:3
						wire oRdEop;
						// Trace: src/src/rtl/design/svsrc/RdCtrlTop1Ch.sv:43:3
						wire oRdVld;
						// Trace: src/src/rtl/design/svsrc/RdCtrlTop1Ch.sv:44:3
						wire [31:0] oRdData;
						// Trace: src/src/rtl/design/svsrc/RdCtrlTop1Ch.sv:45:3
						wire iRdRdy;
						// Trace: src/src/rtl/design/svsrc/RdCtrlTop1Ch.sv:46:3
						wire oRdLast;
						// Trace: src/src/rtl/design/svsrc/RdCtrlTop1Ch.sv:48:3
						wire [($clog2(WRR_WEIGHT_NUM) >= 0 ? (8 * ($clog2(WRR_WEIGHT_NUM) + 1)) - 1 : (8 * (1 - $clog2(WRR_WEIGHT_NUM))) + ($clog2(WRR_WEIGHT_NUM) - 1)):($clog2(WRR_WEIGHT_NUM) >= 0 ? 0 : $clog2(WRR_WEIGHT_NUM) + 0)] iWeight;
						// Trace: src/src/rtl/design/svsrc/RdCtrlTop1Ch.sv:49:3
						wire iWeightLoad;
						// Trace: src/src/rtl/design/svsrc/RdCtrlTop1Ch.sv:52:3
						localparam TAG_QUEUE_WIDTH = 20;
						// Trace: src/src/rtl/design/svsrc/RdCtrlTop1Ch.sv:54:3
						// expanded interface instance: tagQueueIn
						localparam _param_36243_DW = TAG_QUEUE_WIDTH;
						localparam _param_36243_AW = 1;
						genvar _arr_36243;
						for (_arr_36243 = 0; _arr_36243 <= 7; _arr_36243 = _arr_36243 + 1) begin : tagQueueIn
							// Trace: src/src/rtl/design/svsrc/interface_list.sv:64:33
							localparam DW = _param_36243_DW;
							// Trace: src/src/rtl/design/svsrc/interface_list.sv:64:52
							localparam AW = _param_36243_AW;
							// Trace: src/src/rtl/design/svsrc/interface_list.sv:65:3
							wire [19:0] Pld;
							// Trace: src/src/rtl/design/svsrc/interface_list.sv:66:3
							wire [0:0] Dst;
							// Trace: src/src/rtl/design/svsrc/interface_list.sv:67:3
							wire Vld;
							// Trace: src/src/rtl/design/svsrc/interface_list.sv:68:3
							wire Rdy;
							// Trace: src/src/rtl/design/svsrc/interface_list.sv:69:3
							// Trace: src/src/rtl/design/svsrc/interface_list.sv:75:3
						end
						// Trace: src/src/rtl/design/svsrc/RdCtrlTop1Ch.sv:55:3
						// expanded interface instance: tagQueueOut
						localparam _param_ACDEB_DW = TAG_QUEUE_WIDTH;
						localparam _param_ACDEB_AW = 1;
						genvar _arr_ACDEB;
						for (_arr_ACDEB = 0; _arr_ACDEB <= 7; _arr_ACDEB = _arr_ACDEB + 1) begin : tagQueueOut
							// Trace: src/src/rtl/design/svsrc/interface_list.sv:64:33
							localparam DW = _param_ACDEB_DW;
							// Trace: src/src/rtl/design/svsrc/interface_list.sv:64:52
							localparam AW = _param_ACDEB_AW;
							// Trace: src/src/rtl/design/svsrc/interface_list.sv:65:3
							wire [19:0] Pld;
							// Trace: src/src/rtl/design/svsrc/interface_list.sv:66:3
							wire [0:0] Dst;
							// Trace: src/src/rtl/design/svsrc/interface_list.sv:67:3
							wire Vld;
							// Trace: src/src/rtl/design/svsrc/interface_list.sv:68:3
							wire Rdy;
							// Trace: src/src/rtl/design/svsrc/interface_list.sv:69:3
							// Trace: src/src/rtl/design/svsrc/interface_list.sv:75:3
						end
						// Trace: src/src/rtl/design/svsrc/RdCtrlTop1Ch.sv:56:3
						// expanded interface instance: tagDrop
						localparam _param_642E1_DW = TAG_QUEUE_WIDTH;
						localparam _param_642E1_AW = 1;
						if (1) begin : tagDrop
							// Trace: src/src/rtl/design/svsrc/interface_list.sv:64:33
							localparam DW = _param_642E1_DW;
							// Trace: src/src/rtl/design/svsrc/interface_list.sv:64:52
							localparam AW = _param_642E1_AW;
							// Trace: src/src/rtl/design/svsrc/interface_list.sv:65:3
							wire [19:0] Pld;
							// Trace: src/src/rtl/design/svsrc/interface_list.sv:66:3
							wire [0:0] Dst;
							// Trace: src/src/rtl/design/svsrc/interface_list.sv:67:3
							wire Vld;
							// Trace: src/src/rtl/design/svsrc/interface_list.sv:68:3
							wire Rdy;
							// Trace: src/src/rtl/design/svsrc/interface_list.sv:69:3
							// Trace: src/src/rtl/design/svsrc/interface_list.sv:75:3
						end
						// Trace: src/src/rtl/design/svsrc/RdCtrlTop1Ch.sv:57:3
						// expanded interface instance: tagQueue
						localparam _param_0AAC6_DW = TAG_QUEUE_WIDTH;
						localparam _param_0AAC6_AW = 1;
						if (1) begin : tagQueue
							// Trace: src/src/rtl/design/svsrc/interface_list.sv:64:33
							localparam DW = _param_0AAC6_DW;
							// Trace: src/src/rtl/design/svsrc/interface_list.sv:64:52
							localparam AW = _param_0AAC6_AW;
							// Trace: src/src/rtl/design/svsrc/interface_list.sv:65:3
							wire [19:0] Pld;
							// Trace: src/src/rtl/design/svsrc/interface_list.sv:66:3
							wire [0:0] Dst;
							// Trace: src/src/rtl/design/svsrc/interface_list.sv:67:3
							wire Vld;
							// Trace: src/src/rtl/design/svsrc/interface_list.sv:68:3
							wire Rdy;
							// Trace: src/src/rtl/design/svsrc/interface_list.sv:69:3
							// Trace: src/src/rtl/design/svsrc/interface_list.sv:75:3
						end
						// Trace: src/src/rtl/design/svsrc/RdCtrlTop1Ch.sv:59:3
						// expanded module instance: U_TAGRX
						localparam _bbase_010B1_iTagIn = _gv_i_7 + 0;
						localparam _bbase_010B1_oTagQueueOut = 0;
						if (1) begin : U_TAGRX
							// Trace: src/src/rtl/design/svsrc/TagRx.sv:26:3
							wire iClk;
							// Trace: src/src/rtl/design/svsrc/TagRx.sv:27:3
							wire iRst_n;
							// Trace: src/src/rtl/design/svsrc/TagRx.sv:29:3
							localparam _mbase_iTagIn = _bbase_010B1_iTagIn;
							// Trace: src/src/rtl/design/svsrc/TagRx.sv:31:3
							localparam _mbase_oTagQueueOut = 0;
							// Trace: src/src/rtl/design/svsrc/TagRx.sv:32:3
							// removed modport instance oTagDropOut
							// Trace: src/src/rtl/design/svsrc/TagRx.sv:37:3
							wire [2:0] rxTagPri;
							// Trace: src/src/rtl/design/svsrc/TagRx.sv:38:3
							wire [3:0] rxTagSrcPort;
							// Trace: src/src/rtl/design/svsrc/TagRx.sv:39:3
							wire [15:0] rxTagMsg;
							// Trace: src/src/rtl/design/svsrc/TagRx.sv:42:3
							reg [2:0] tagPri;
							// Trace: src/src/rtl/design/svsrc/TagRx.sv:43:3
							reg [3:0] tagSrcPort;
							// Trace: src/src/rtl/design/svsrc/TagRx.sv:44:3
							reg [15:0] tagMsg;
							// Trace: src/src/rtl/design/svsrc/TagRx.sv:46:3
							wire [7:0] queueOutVld;
							// Trace: src/src/rtl/design/svsrc/TagRx.sv:47:3
							wire [7:0] queueOutRdy;
							// Trace: src/src/rtl/design/svsrc/TagRx.sv:49:3
							genvar _gv_i_11;
							// Trace: src/src/rtl/design/svsrc/TagRx.sv:51:3
							assign {rxTagPri, rxTagMsg, rxTagSrcPort} = RdScheTopWrapper.U_RD_SCHE_TOP_SV.tagCrsbarOut[_mbase_iTagIn].Pld;
							// Trace: src/src/rtl/design/svsrc/TagRx.sv:53:3
							assign RdScheTopWrapper.U_RD_SCHE_TOP_SV.U_RDCTRLTOP16.genblk1[_gv_i_7].U_RD_CHN.tagDrop.Pld = {tagMsg, tagSrcPort};
							// Trace: src/src/rtl/design/svsrc/TagRx.sv:54:3
							for (_gv_i_11 = 0; _gv_i_11 < 8; _gv_i_11 = _gv_i_11 + 1) begin : GEN_QUEUE_PLD
								localparam i = _gv_i_11;
								// Trace: src/src/rtl/design/svsrc/TagRx.sv:56:7
								assign RdScheTopWrapper.U_RD_SCHE_TOP_SV.U_RDCTRLTOP16.genblk1[_gv_i_7].U_RD_CHN.tagQueueIn[i + _mbase_oTagQueueOut].Pld = {tagMsg, tagSrcPort};
								// Trace: src/src/rtl/design/svsrc/TagRx.sv:57:7
								assign RdScheTopWrapper.U_RD_SCHE_TOP_SV.U_RDCTRLTOP16.genblk1[_gv_i_7].U_RD_CHN.tagQueueIn[i + _mbase_oTagQueueOut].Vld = queueOutVld[i];
								// Trace: src/src/rtl/design/svsrc/TagRx.sv:58:7
								assign queueOutRdy[i] = RdScheTopWrapper.U_RD_SCHE_TOP_SV.U_RDCTRLTOP16.genblk1[_gv_i_7].U_RD_CHN.tagQueueIn[i + _mbase_oTagQueueOut].Rdy;
							end
							// Trace: src/src/rtl/design/svsrc/TagRx.sv:63:3
							reg [1:0] fsmCstate;
							// Trace: src/src/rtl/design/svsrc/TagRx.sv:64:3
							reg [1:0] fsmNstate;
							// Trace: src/src/rtl/design/svsrc/TagRx.sv:66:3
							localparam FSM_IDLE = 2'b00;
							// Trace: src/src/rtl/design/svsrc/TagRx.sv:67:3
							localparam FSM_FETCH = 2'b01;
							// Trace: src/src/rtl/design/svsrc/TagRx.sv:68:3
							localparam FSM_DISPATCH = 2'b10;
							// Trace: src/src/rtl/design/svsrc/TagRx.sv:69:3
							localparam FSM_DROP = 2'b11;
							// Trace: src/src/rtl/design/svsrc/TagRx.sv:71:3
							wire signed [31:0] j;
							// Trace: src/src/rtl/design/svsrc/TagRx.sv:73:3
							always @(posedge iClk or negedge iRst_n)
								// Trace: src/src/rtl/design/svsrc/TagRx.sv:74:5
								if (!iRst_n)
									// Trace: src/src/rtl/design/svsrc/TagRx.sv:75:7
									fsmCstate <= FSM_IDLE;
								else
									// Trace: src/src/rtl/design/svsrc/TagRx.sv:77:7
									fsmCstate <= fsmNstate;
							// Trace: src/src/rtl/design/svsrc/TagRx.sv:81:3
							always @(*)
								// Trace: src/src/rtl/design/svsrc/TagRx.sv:82:5
								case (fsmCstate)
									FSM_IDLE:
										// Trace: src/src/rtl/design/svsrc/TagRx.sv:84:9
										if (RdScheTopWrapper.U_RD_SCHE_TOP_SV.tagCrsbarOut[_mbase_iTagIn].Vld && RdScheTopWrapper.U_RD_SCHE_TOP_SV.tagCrsbarOut[_mbase_iTagIn].Rdy)
											// Trace: src/src/rtl/design/svsrc/TagRx.sv:85:11
											fsmNstate = FSM_FETCH;
										else
											// Trace: src/src/rtl/design/svsrc/TagRx.sv:87:11
											fsmNstate = FSM_IDLE;
									FSM_FETCH:
										// Trace: src/src/rtl/design/svsrc/TagRx.sv:91:9
										if (queueOutRdy[tagPri])
											// Trace: src/src/rtl/design/svsrc/TagRx.sv:92:11
											fsmNstate = FSM_DISPATCH;
										else
											// Trace: src/src/rtl/design/svsrc/TagRx.sv:94:11
											fsmNstate = FSM_DROP;
									FSM_DISPATCH:
										// Trace: src/src/rtl/design/svsrc/TagRx.sv:98:9
										if (queueOutVld[tagPri] && queueOutRdy[tagPri])
											// Trace: src/src/rtl/design/svsrc/TagRx.sv:99:11
											fsmNstate = FSM_IDLE;
										else
											// Trace: src/src/rtl/design/svsrc/TagRx.sv:101:11
											fsmNstate = FSM_DISPATCH;
									FSM_DROP:
										// Trace: src/src/rtl/design/svsrc/TagRx.sv:105:9
										if (RdScheTopWrapper.U_RD_SCHE_TOP_SV.U_RDCTRLTOP16.genblk1[_gv_i_7].U_RD_CHN.tagDrop.Vld && RdScheTopWrapper.U_RD_SCHE_TOP_SV.U_RDCTRLTOP16.genblk1[_gv_i_7].U_RD_CHN.tagDrop.Rdy)
											// Trace: src/src/rtl/design/svsrc/TagRx.sv:106:11
											fsmNstate = FSM_IDLE;
										else
											// Trace: src/src/rtl/design/svsrc/TagRx.sv:108:11
											fsmNstate = FSM_DROP;
									default:
										// Trace: src/src/rtl/design/svsrc/TagRx.sv:111:17
										fsmNstate = FSM_IDLE;
								endcase
							// Trace: src/src/rtl/design/svsrc/TagRx.sv:115:3
							always @(posedge iClk or negedge iRst_n)
								// Trace: src/src/rtl/design/svsrc/TagRx.sv:116:5
								if (!iRst_n) begin
									// Trace: src/src/rtl/design/svsrc/TagRx.sv:117:7
									tagPri <= 0;
									// Trace: src/src/rtl/design/svsrc/TagRx.sv:118:7
									tagSrcPort <= 0;
									// Trace: src/src/rtl/design/svsrc/TagRx.sv:119:7
									tagMsg <= 0;
								end
								else if (RdScheTopWrapper.U_RD_SCHE_TOP_SV.tagCrsbarOut[_mbase_iTagIn].Vld && RdScheTopWrapper.U_RD_SCHE_TOP_SV.tagCrsbarOut[_mbase_iTagIn].Rdy) begin
									// Trace: src/src/rtl/design/svsrc/TagRx.sv:121:7
									tagPri <= rxTagPri;
									// Trace: src/src/rtl/design/svsrc/TagRx.sv:122:7
									tagSrcPort <= rxTagSrcPort;
									// Trace: src/src/rtl/design/svsrc/TagRx.sv:123:7
									tagMsg <= rxTagMsg;
								end
								else begin
									// Trace: src/src/rtl/design/svsrc/TagRx.sv:125:7
									tagPri <= tagPri;
									// Trace: src/src/rtl/design/svsrc/TagRx.sv:126:7
									tagSrcPort <= tagSrcPort;
									// Trace: src/src/rtl/design/svsrc/TagRx.sv:127:7
									tagMsg <= tagMsg;
								end
							// Trace: src/src/rtl/design/svsrc/TagRx.sv:131:3
							assign RdScheTopWrapper.U_RD_SCHE_TOP_SV.tagCrsbarOut[_mbase_iTagIn].Rdy = fsmCstate == FSM_IDLE;
							// Trace: src/src/rtl/design/svsrc/TagRx.sv:132:3
							assign RdScheTopWrapper.U_RD_SCHE_TOP_SV.U_RDCTRLTOP16.genblk1[_gv_i_7].U_RD_CHN.tagDrop.Vld = fsmCstate == FSM_DROP;
							// Trace: src/src/rtl/design/svsrc/TagRx.sv:134:3
							for (_gv_i_11 = 0; _gv_i_11 < 8; _gv_i_11 = _gv_i_11 + 1) begin : GEN_QUEUE_VLD
								localparam i = _gv_i_11;
								// Trace: src/src/rtl/design/svsrc/TagRx.sv:136:7
								assign queueOutVld[i] = (fsmCstate == FSM_DISPATCH) && (tagPri == i);
							end
						end
						assign U_TAGRX.iClk = iClk;
						assign U_TAGRX.iRst_n = iRst_n;
						// Trace: src/src/rtl/design/svsrc/RdCtrlTop1Ch.sv:67:3
						genvar _gv_i_8;
						// Trace: src/src/rtl/design/svsrc/RdCtrlTop1Ch.sv:68:3
						for (_gv_i_8 = 0; _gv_i_8 < PRI_NUM; _gv_i_8 = _gv_i_8 + 1) begin : GEN_PRI_FIFO
							localparam i = _gv_i_8;
							// Trace: src/src/rtl/design/svsrc/RdCtrlTop1Ch.sv:70:7
							// expanded module instance: U_PRIFIFO
							localparam _bbase_3FE19_iDcpIn = _gv_i_8;
							localparam _bbase_3FE19_oDcpOut = _gv_i_8;
							localparam _param_3FE19_DATA_WIDTH = TAG_QUEUE_WIDTH;
							localparam _param_3FE19_DEPTH = PRI_DEPTH;
							if (1) begin : U_PRIFIFO
								// Trace: src/src/rtl/design/svsrc/DcpFifo.sv:3:13
								localparam [0:0] FALL_THROUGH = 1'b0;
								// Trace: src/src/rtl/design/svsrc/DcpFifo.sv:5:13
								localparam [31:0] DATA_WIDTH = _param_3FE19_DATA_WIDTH;
								// Trace: src/src/rtl/design/svsrc/DcpFifo.sv:7:13
								localparam [31:0] DEPTH = _param_3FE19_DEPTH;
								// Trace: src/src/rtl/design/svsrc/DcpFifo.sv:9:13
								localparam [31:0] ADDR_DEPTH = (DEPTH > 1 ? $clog2(DEPTH) : 1);
								// Trace: src/src/rtl/design/svsrc/DcpFifo.sv:12:3
								wire iClk;
								// Trace: src/src/rtl/design/svsrc/DcpFifo.sv:13:3
								wire iRst_n;
								// Trace: src/src/rtl/design/svsrc/DcpFifo.sv:15:3
								localparam _mbase_iDcpIn = _bbase_3FE19_iDcpIn;
								// Trace: src/src/rtl/design/svsrc/DcpFifo.sv:16:3
								localparam _mbase_oDcpOut = _bbase_3FE19_oDcpOut;
								// Trace: src/src/rtl/design/svsrc/DcpFifo.sv:17:3
								wire [ADDR_DEPTH - 1:0] oUsage;
								// Trace: src/src/rtl/design/svsrc/DcpFifo.sv:18:3
								wire iTestmode;
								// Trace: src/src/rtl/design/svsrc/DcpFifo.sv:19:3
								wire iFlush;
								// Trace: src/src/rtl/design/svsrc/DcpFifo.sv:21:3
								// removed localparam type T
								// Trace: src/src/rtl/design/svsrc/DcpFifo.sv:23:3
								// expanded interface instance: fifoOut
								localparam _param_492B2_DW = DATA_WIDTH;
								localparam _param_492B2_AW = 1;
								if (1) begin : fifoOut
									// Trace: src/src/rtl/design/svsrc/interface_list.sv:64:33
									localparam DW = _param_492B2_DW;
									// Trace: src/src/rtl/design/svsrc/interface_list.sv:64:52
									localparam AW = _param_492B2_AW;
									// Trace: src/src/rtl/design/svsrc/interface_list.sv:65:3
									wire [19:0] Pld;
									// Trace: src/src/rtl/design/svsrc/interface_list.sv:66:3
									wire [0:0] Dst;
									// Trace: src/src/rtl/design/svsrc/interface_list.sv:67:3
									wire Vld;
									// Trace: src/src/rtl/design/svsrc/interface_list.sv:68:3
									wire Rdy;
									// Trace: src/src/rtl/design/svsrc/interface_list.sv:69:3
									// Trace: src/src/rtl/design/svsrc/interface_list.sv:75:3
								end
								// Trace: src/src/rtl/design/svsrc/DcpFifo.sv:25:5
								wire push;
								wire pop;
								// Trace: src/src/rtl/design/svsrc/DcpFifo.sv:26:5
								wire empty;
								wire full;
								// Trace: src/src/rtl/design/svsrc/DcpFifo.sv:28:5
								assign push = RdScheTopWrapper.U_RD_SCHE_TOP_SV.U_RDCTRLTOP16.genblk1[_gv_i_7].U_RD_CHN.tagQueueIn[_mbase_iDcpIn].Vld & ~full;
								// Trace: src/src/rtl/design/svsrc/DcpFifo.sv:29:5
								assign pop = fifoOut.Rdy & ~empty;
								// Trace: src/src/rtl/design/svsrc/DcpFifo.sv:30:5
								assign RdScheTopWrapper.U_RD_SCHE_TOP_SV.U_RDCTRLTOP16.genblk1[_gv_i_7].U_RD_CHN.tagQueueIn[_mbase_iDcpIn].Rdy = ~full;
								// Trace: src/src/rtl/design/svsrc/DcpFifo.sv:31:5
								assign fifoOut.Vld = ~empty;
								// Trace: src/src/rtl/design/svsrc/DcpFifo.sv:33:5
								fifo_v3_7703C #(
									.FALL_THROUGH(FALL_THROUGH),
									.DATA_WIDTH(DATA_WIDTH),
									.DEPTH(DEPTH)
								) U_FIFO(
									.clk_i(iClk),
									.rst_ni(iRst_n),
									.flush_i(iFlush),
									.testmode_i(iTestmode),
									.full_o(full),
									.empty_o(empty),
									.usage_o(oUsage),
									.data_i(RdScheTopWrapper.U_RD_SCHE_TOP_SV.U_RDCTRLTOP16.genblk1[_gv_i_7].U_RD_CHN.tagQueueIn[_mbase_iDcpIn].Pld),
									.push_i(push),
									.data_o(fifoOut.Pld),
									.pop_i(pop)
								);
								// Trace: src/src/rtl/design/svsrc/DcpFifo.sv:52:3
								gnrl_buf #(
									.DW(DATA_WIDTH),
									.CUT_RDY(1)
								) U_OUTBUF(
									.clk_i(iClk),
									.rst_n_i(iRst_n),
									.din_i(fifoOut.Pld),
									.din_vld_i(fifoOut.Vld),
									.din_rdy_o(fifoOut.Rdy),
									.dout_o(RdScheTopWrapper.U_RD_SCHE_TOP_SV.U_RDCTRLTOP16.genblk1[_gv_i_7].U_RD_CHN.tagQueueOut[_mbase_oDcpOut].Pld),
									.dout_vld_o(RdScheTopWrapper.U_RD_SCHE_TOP_SV.U_RDCTRLTOP16.genblk1[_gv_i_7].U_RD_CHN.tagQueueOut[_mbase_oDcpOut].Vld),
									.dout_rdy_i(RdScheTopWrapper.U_RD_SCHE_TOP_SV.U_RDCTRLTOP16.genblk1[_gv_i_7].U_RD_CHN.tagQueueOut[_mbase_oDcpOut].Rdy)
								);
							end
							assign U_PRIFIFO.iClk = iClk;
							assign U_PRIFIFO.iRst_n = iRst_n;
							assign U_PRIFIFO.iTestmode = 1'b0;
							assign U_PRIFIFO.iFlush = 1'b0;
						end
						// Trace: src/src/rtl/design/svsrc/RdCtrlTop1Ch.sv:85:3
						// expanded module instance: U_DCP_WRR_ARBITER
						localparam _bbase_ECC17_iDcpIn = 0;
						localparam _param_ECC17_DW = TAG_QUEUE_WIDTH;
						localparam _param_ECC17_WEIGHT_NUM = WRR_WEIGHT_NUM;
						localparam _param_ECC17_ARB_NUM = PRI_NUM;
						if (1) begin : U_DCP_WRR_ARBITER
							// Trace: src/src/rtl/design/svsrc/DcpWrrArbiter.sv:25:13
							localparam DW = _param_ECC17_DW;
							// Trace: src/src/rtl/design/svsrc/DcpWrrArbiter.sv:26:13
							localparam ARB_NUM = _param_ECC17_ARB_NUM;
							// Trace: src/src/rtl/design/svsrc/DcpWrrArbiter.sv:27:13
							localparam WEIGHT_NUM = _param_ECC17_WEIGHT_NUM;
							// Trace: src/src/rtl/design/svsrc/DcpWrrArbiter.sv:29:3
							wire iClk;
							// Trace: src/src/rtl/design/svsrc/DcpWrrArbiter.sv:30:3
							wire iRst_n;
							// Trace: src/src/rtl/design/svsrc/DcpWrrArbiter.sv:32:3
							localparam _mbase_iDcpIn = 0;
							// Trace: src/src/rtl/design/svsrc/DcpWrrArbiter.sv:33:3
							// removed modport instance oDcpOut
							// Trace: src/src/rtl/design/svsrc/DcpWrrArbiter.sv:35:3
							wire [($clog2(WEIGHT_NUM) >= 0 ? (8 * ($clog2(WEIGHT_NUM) + 1)) - 1 : (8 * (1 - $clog2(WEIGHT_NUM))) + ($clog2(WEIGHT_NUM) - 1)):($clog2(WEIGHT_NUM) >= 0 ? 0 : $clog2(WEIGHT_NUM) + 0)] iWeight;
							// Trace: src/src/rtl/design/svsrc/DcpWrrArbiter.sv:36:3
							wire iWeightLoad;
							// Trace: src/src/rtl/design/svsrc/DcpWrrArbiter.sv:38:3
							wire [7:0] iReq;
							// Trace: src/src/rtl/design/svsrc/DcpWrrArbiter.sv:39:3
							wire [7:0] oGnt;
							// Trace: src/src/rtl/design/svsrc/DcpWrrArbiter.sv:40:3
							wire [159:0] iData;
							// Trace: src/src/rtl/design/svsrc/DcpWrrArbiter.sv:42:3
							wire oReq;
							// Trace: src/src/rtl/design/svsrc/DcpWrrArbiter.sv:43:3
							wire iGnt;
							// Trace: src/src/rtl/design/svsrc/DcpWrrArbiter.sv:44:3
							wire [19:0] oData;
							// Trace: src/src/rtl/design/svsrc/DcpWrrArbiter.sv:46:3
							genvar _gv_i_6;
							// Trace: src/src/rtl/design/svsrc/DcpWrrArbiter.sv:47:3
							for (_gv_i_6 = 0; _gv_i_6 < ARB_NUM; _gv_i_6 = _gv_i_6 + 1) begin : genblk1
								localparam i = _gv_i_6;
								// Trace: src/src/rtl/design/svsrc/DcpWrrArbiter.sv:49:7
								assign iReq[i] = RdScheTopWrapper.U_RD_SCHE_TOP_SV.U_RDCTRLTOP16.genblk1[_gv_i_7].U_RD_CHN.tagQueueOut[i + _mbase_iDcpIn].Vld;
								// Trace: src/src/rtl/design/svsrc/DcpWrrArbiter.sv:50:7
								assign iData[i * 20+:20] = {RdScheTopWrapper.U_RD_SCHE_TOP_SV.U_RDCTRLTOP16.genblk1[_gv_i_7].U_RD_CHN.tagQueueOut[i + _mbase_iDcpIn].Pld};
								// Trace: src/src/rtl/design/svsrc/DcpWrrArbiter.sv:51:7
								assign RdScheTopWrapper.U_RD_SCHE_TOP_SV.U_RDCTRLTOP16.genblk1[_gv_i_7].U_RD_CHN.tagQueueOut[i + _mbase_iDcpIn].Rdy = oGnt[i];
							end
							// Trace: src/src/rtl/design/svsrc/DcpWrrArbiter.sv:55:3
							assign RdScheTopWrapper.U_RD_SCHE_TOP_SV.U_RDCTRLTOP16.genblk1[_gv_i_7].U_RD_CHN.tagQueue.Vld = oReq;
							// Trace: src/src/rtl/design/svsrc/DcpWrrArbiter.sv:56:3
							assign RdScheTopWrapper.U_RD_SCHE_TOP_SV.U_RDCTRLTOP16.genblk1[_gv_i_7].U_RD_CHN.tagQueue.Pld = oData;
							// Trace: src/src/rtl/design/svsrc/DcpWrrArbiter.sv:57:3
							assign iGnt = RdScheTopWrapper.U_RD_SCHE_TOP_SV.U_RDCTRLTOP16.genblk1[_gv_i_7].U_RD_CHN.tagQueue.Rdy;
							// Trace: src/src/rtl/design/svsrc/DcpWrrArbiter.sv:59:1
							WrrArbiter #(
								.DW(DW),
								.ARB_NUM(ARB_NUM),
								.WEIGHT_NUM(WEIGHT_NUM)
							) U_WRRARBITER(
								.iRst_n(iRst_n),
								.iClk(iClk),
								.iReq(iReq),
								.oGnt(oGnt),
								.iData(iData),
								.oReq(oReq),
								.iGnt(iGnt),
								.oData(oData),
								.iWeightLoad(iWeightLoad),
								.iWeight(iWeight)
							);
						end
						assign U_DCP_WRR_ARBITER.iClk = iClk;
						assign U_DCP_WRR_ARBITER.iRst_n = iRst_n;
						assign U_DCP_WRR_ARBITER.iWeightLoad = iWeightLoad;
						assign U_DCP_WRR_ARBITER.iWeight = iWeight;
						// Trace: src/src/rtl/design/svsrc/RdCtrlTop1Ch.sv:98:3
						// expanded module instance: U_PORT_CTRL
						localparam _bbase_0F4F7_oRdCmd = _gv_i_7 + 0;
						localparam _bbase_0F4F7_iRdData = _gv_i_7 + 0;
						localparam _param_0F4F7_PORT_ADDR = PORT_ADDR;
						if (1) begin : U_PORT_CTRL
							// Trace: src/src/rtl/design/svsrc/PortCtrl.sv:26:13
							localparam PORT_ADDR = _param_0F4F7_PORT_ADDR;
							// Trace: src/src/rtl/design/svsrc/PortCtrl.sv:28:3
							wire iClk;
							// Trace: src/src/rtl/design/svsrc/PortCtrl.sv:29:3
							wire iRst_n;
							// Trace: src/src/rtl/design/svsrc/PortCtrl.sv:31:3
							// removed modport instance iTagQueueIn
							// Trace: src/src/rtl/design/svsrc/PortCtrl.sv:32:3
							// removed modport instance iTagDropIn
							// Trace: src/src/rtl/design/svsrc/PortCtrl.sv:34:3
							localparam _mbase_oRdCmd = _bbase_0F4F7_oRdCmd;
							// Trace: src/src/rtl/design/svsrc/PortCtrl.sv:36:3
							localparam _mbase_iRdData = _bbase_0F4F7_iRdData;
							// Trace: src/src/rtl/design/svsrc/PortCtrl.sv:38:3
							reg oRdSop;
							// Trace: src/src/rtl/design/svsrc/PortCtrl.sv:39:3
							reg oRdEop;
							// Trace: src/src/rtl/design/svsrc/PortCtrl.sv:40:3
							wire oRdVld;
							// Trace: src/src/rtl/design/svsrc/PortCtrl.sv:41:3
							wire [31:0] oRdData;
							// Trace: src/src/rtl/design/svsrc/PortCtrl.sv:42:3
							wire iRdRdy;
							// Trace: src/src/rtl/design/svsrc/PortCtrl.sv:43:3
							wire oRdLast;
							// Trace: src/src/rtl/design/svsrc/PortCtrl.sv:46:3
							reg [3:0] queueSrcPort;
							// Trace: src/src/rtl/design/svsrc/PortCtrl.sv:47:3
							wire [3:0] queueDstPort;
							// Trace: src/src/rtl/design/svsrc/PortCtrl.sv:48:3
							reg [15:0] queueMsg;
							// Trace: src/src/rtl/design/svsrc/PortCtrl.sv:50:3
							reg [3:0] dropSrcPort;
							// Trace: src/src/rtl/design/svsrc/PortCtrl.sv:51:3
							reg [15:0] dropMsg;
							// Trace: src/src/rtl/design/svsrc/PortCtrl.sv:53:3
							wire rdCmdDrop;
							// Trace: src/src/rtl/design/svsrc/PortCtrl.sv:55:3
							wire rawRdLast;
							// Trace: src/src/rtl/design/svsrc/PortCtrl.sv:56:3
							wire [31:0] rawRdData;
							// Trace: src/src/rtl/design/svsrc/PortCtrl.sv:58:3
							wire tmpRdRdy;
							// Trace: src/src/rtl/design/svsrc/PortCtrl.sv:59:3
							wire tmpRdVld;
							// Trace: src/src/rtl/design/svsrc/PortCtrl.sv:60:3
							wire tmpRdLast;
							// Trace: src/src/rtl/design/svsrc/PortCtrl.sv:61:3
							reg [1:0] fsmCstate_d;
							// Trace: src/src/rtl/design/svsrc/PortCtrl.sv:63:3
							assign queueDstPort = PORT_ADDR;
							// Trace: src/src/rtl/design/svsrc/PortCtrl.sv:69:3
							always @(posedge iClk or negedge iRst_n)
								// Trace: src/src/rtl/design/svsrc/PortCtrl.sv:70:5
								if (!iRst_n) begin
									// Trace: src/src/rtl/design/svsrc/PortCtrl.sv:71:7
									queueMsg <= 'b0;
									// Trace: src/src/rtl/design/svsrc/PortCtrl.sv:72:7
									queueSrcPort <= 'b0;
								end
								else if (RdScheTopWrapper.U_RD_SCHE_TOP_SV.U_RDCTRLTOP16.genblk1[_gv_i_7].U_RD_CHN.tagQueue.Vld && RdScheTopWrapper.U_RD_SCHE_TOP_SV.U_RDCTRLTOP16.genblk1[_gv_i_7].U_RD_CHN.tagQueue.Rdy)
									// Trace: src/src/rtl/design/svsrc/PortCtrl.sv:74:7
									{queueMsg, queueSrcPort} <= RdScheTopWrapper.U_RD_SCHE_TOP_SV.U_RDCTRLTOP16.genblk1[_gv_i_7].U_RD_CHN.tagQueue.Pld;
								else
									// Trace: src/src/rtl/design/svsrc/PortCtrl.sv:76:7
									{queueMsg, queueSrcPort} <= {queueMsg, queueSrcPort};
							// Trace: src/src/rtl/design/svsrc/PortCtrl.sv:80:3
							always @(posedge iClk or negedge iRst_n)
								// Trace: src/src/rtl/design/svsrc/PortCtrl.sv:81:5
								if (!iRst_n) begin
									// Trace: src/src/rtl/design/svsrc/PortCtrl.sv:82:7
									dropMsg <= 'b0;
									// Trace: src/src/rtl/design/svsrc/PortCtrl.sv:83:7
									dropSrcPort <= 'b0;
								end
								else if (RdScheTopWrapper.U_RD_SCHE_TOP_SV.U_RDCTRLTOP16.genblk1[_gv_i_7].U_RD_CHN.tagDrop.Vld && RdScheTopWrapper.U_RD_SCHE_TOP_SV.U_RDCTRLTOP16.genblk1[_gv_i_7].U_RD_CHN.tagDrop.Rdy)
									// Trace: src/src/rtl/design/svsrc/PortCtrl.sv:85:7
									{dropMsg, dropSrcPort} <= RdScheTopWrapper.U_RD_SCHE_TOP_SV.U_RDCTRLTOP16.genblk1[_gv_i_7].U_RD_CHN.tagDrop.Pld;
								else
									// Trace: src/src/rtl/design/svsrc/PortCtrl.sv:87:7
									{dropMsg, dropSrcPort} <= {dropMsg, dropSrcPort};
							// Trace: src/src/rtl/design/svsrc/PortCtrl.sv:91:3
							assign {rawRdData, rawRdLast} = RdScheTopWrapper.U_RD_SCHE_TOP_SV.rddataCrsbarOut[_mbase_iRdData].Pld;
							// Trace: src/src/rtl/design/svsrc/PortCtrl.sv:94:3
							localparam FSM_IDLE = 2'b00;
							// Trace: src/src/rtl/design/svsrc/PortCtrl.sv:95:3
							localparam FSM_DROP = 2'b01;
							// Trace: src/src/rtl/design/svsrc/PortCtrl.sv:96:3
							localparam FSM_RDCMD = 2'b10;
							// Trace: src/src/rtl/design/svsrc/PortCtrl.sv:97:3
							localparam FSM_RDDATA = 2'b11;
							// Trace: src/src/rtl/design/svsrc/PortCtrl.sv:99:3
							reg [1:0] fsmCstate;
							reg [1:0] fsmNstate;
							// Trace: src/src/rtl/design/svsrc/PortCtrl.sv:103:3
							always @(posedge iClk or negedge iRst_n)
								// Trace: src/src/rtl/design/svsrc/PortCtrl.sv:104:5
								if (!iRst_n)
									// Trace: src/src/rtl/design/svsrc/PortCtrl.sv:105:7
									fsmCstate <= FSM_IDLE;
								else
									// Trace: src/src/rtl/design/svsrc/PortCtrl.sv:107:7
									fsmCstate <= fsmNstate;
							// Trace: src/src/rtl/design/svsrc/PortCtrl.sv:111:3
							always @(*)
								// Trace: src/src/rtl/design/svsrc/PortCtrl.sv:112:5
								case (fsmCstate)
									FSM_IDLE:
										// Trace: src/src/rtl/design/svsrc/PortCtrl.sv:114:7
										if (RdScheTopWrapper.U_RD_SCHE_TOP_SV.U_RDCTRLTOP16.genblk1[_gv_i_7].U_RD_CHN.tagDrop.Vld && RdScheTopWrapper.U_RD_SCHE_TOP_SV.U_RDCTRLTOP16.genblk1[_gv_i_7].U_RD_CHN.tagDrop.Rdy)
											// Trace: src/src/rtl/design/svsrc/PortCtrl.sv:115:9
											fsmNstate = FSM_DROP;
										else if (RdScheTopWrapper.U_RD_SCHE_TOP_SV.U_RDCTRLTOP16.genblk1[_gv_i_7].U_RD_CHN.tagQueue.Vld && RdScheTopWrapper.U_RD_SCHE_TOP_SV.U_RDCTRLTOP16.genblk1[_gv_i_7].U_RD_CHN.tagQueue.Rdy)
											// Trace: src/src/rtl/design/svsrc/PortCtrl.sv:117:9
											fsmNstate = FSM_RDCMD;
										else
											// Trace: src/src/rtl/design/svsrc/PortCtrl.sv:119:9
											fsmNstate = FSM_IDLE;
									FSM_DROP:
										// Trace: src/src/rtl/design/svsrc/PortCtrl.sv:123:7
										if (RdScheTopWrapper.U_RD_SCHE_TOP_SV.rdcmdCrsbarIn[_mbase_oRdCmd].Vld && RdScheTopWrapper.U_RD_SCHE_TOP_SV.rdcmdCrsbarIn[_mbase_oRdCmd].Rdy)
											// Trace: src/src/rtl/design/svsrc/PortCtrl.sv:124:9
											fsmNstate = FSM_IDLE;
										else
											// Trace: src/src/rtl/design/svsrc/PortCtrl.sv:126:9
											fsmNstate = FSM_DROP;
									FSM_RDCMD:
										// Trace: src/src/rtl/design/svsrc/PortCtrl.sv:130:7
										if (RdScheTopWrapper.U_RD_SCHE_TOP_SV.rdcmdCrsbarIn[_mbase_oRdCmd].Vld && RdScheTopWrapper.U_RD_SCHE_TOP_SV.rdcmdCrsbarIn[_mbase_oRdCmd].Rdy)
											// Trace: src/src/rtl/design/svsrc/PortCtrl.sv:131:9
											fsmNstate = FSM_RDDATA;
										else
											// Trace: src/src/rtl/design/svsrc/PortCtrl.sv:133:9
											fsmNstate = FSM_RDCMD;
									FSM_RDDATA:
										// Trace: src/src/rtl/design/svsrc/PortCtrl.sv:139:7
										if ((tmpRdLast && iRdRdy) && tmpRdVld)
											// Trace: src/src/rtl/design/svsrc/PortCtrl.sv:140:9
											fsmNstate = FSM_IDLE;
										else
											// Trace: src/src/rtl/design/svsrc/PortCtrl.sv:142:9
											fsmNstate = FSM_RDDATA;
									default:
										// Trace: src/src/rtl/design/svsrc/PortCtrl.sv:145:15
										fsmNstate = FSM_IDLE;
								endcase
							// Trace: src/src/rtl/design/svsrc/PortCtrl.sv:153:3
							rr_arb_tree #(
								.NumIn(2),
								.DataWidth(1),
								.AxiVldRdy(1),
								.LockIn(0)
							) U_RR_QUEUE_DROP(
								.rst_ni(iRst_n),
								.clk_i(iClk),
								.req_i({RdScheTopWrapper.U_RD_SCHE_TOP_SV.U_RDCTRLTOP16.genblk1[_gv_i_7].U_RD_CHN.tagDrop.Vld, RdScheTopWrapper.U_RD_SCHE_TOP_SV.U_RDCTRLTOP16.genblk1[_gv_i_7].U_RD_CHN.tagQueue.Vld}),
								.gnt_o({RdScheTopWrapper.U_RD_SCHE_TOP_SV.U_RDCTRLTOP16.genblk1[_gv_i_7].U_RD_CHN.tagDrop.Rdy, RdScheTopWrapper.U_RD_SCHE_TOP_SV.U_RDCTRLTOP16.genblk1[_gv_i_7].U_RD_CHN.tagQueue.Rdy}),
								.data_i(),
								.req_o(),
								.gnt_i(fsmCstate == FSM_IDLE),
								.data_o()
							);
							// Trace: src/src/rtl/design/svsrc/PortCtrl.sv:170:3
							assign rdCmdDrop = fsmCstate == FSM_DROP;
							// Trace: src/src/rtl/design/svsrc/PortCtrl.sv:172:3
							assign RdScheTopWrapper.U_RD_SCHE_TOP_SV.rdcmdCrsbarIn[_mbase_oRdCmd].Vld = ^fsmCstate;
							// Trace: src/src/rtl/design/svsrc/PortCtrl.sv:173:3
							assign RdScheTopWrapper.U_RD_SCHE_TOP_SV.rdcmdCrsbarIn[_mbase_oRdCmd].Pld = (fsmCstate[0] ? {dropMsg, queueDstPort, rdCmdDrop} : {queueMsg, queueDstPort, rdCmdDrop});
							// Trace: src/src/rtl/design/svsrc/PortCtrl.sv:174:3
							assign RdScheTopWrapper.U_RD_SCHE_TOP_SV.rdcmdCrsbarIn[_mbase_oRdCmd].Dst = (fsmCstate[0] ? dropSrcPort : queueSrcPort);
							// Trace: src/src/rtl/design/svsrc/PortCtrl.sv:181:3
							gnrl_buf #(
								.DW(33),
								.CUT_RDY(1)
							) U_INBUF(
								.clk_i(iClk),
								.rst_n_i(iRst_n),
								.din_i({rawRdData, rawRdLast}),
								.din_vld_i(RdScheTopWrapper.U_RD_SCHE_TOP_SV.rddataCrsbarOut[_mbase_iRdData].Vld),
								.din_rdy_o(RdScheTopWrapper.U_RD_SCHE_TOP_SV.rddataCrsbarOut[_mbase_iRdData].Rdy),
								.dout_o({oRdData, tmpRdLast}),
								.dout_vld_o(tmpRdVld),
								.dout_rdy_i(tmpRdRdy)
							);
							// Trace: src/src/rtl/design/svsrc/PortCtrl.sv:195:3
							always @(posedge iClk or negedge iRst_n)
								// Trace: src/src/rtl/design/svsrc/PortCtrl.sv:196:5
								if (!iRst_n)
									// Trace: src/src/rtl/design/svsrc/PortCtrl.sv:197:7
									fsmCstate_d <= FSM_IDLE;
								else
									// Trace: src/src/rtl/design/svsrc/PortCtrl.sv:199:7
									fsmCstate_d <= fsmCstate;
							// Trace: src/src/rtl/design/svsrc/PortCtrl.sv:203:3
							always @(posedge iClk or negedge iRst_n)
								// Trace: src/src/rtl/design/svsrc/PortCtrl.sv:204:5
								if (!iRst_n)
									// Trace: src/src/rtl/design/svsrc/PortCtrl.sv:205:7
									oRdSop <= 1'b0;
								else
									// Trace: src/src/rtl/design/svsrc/PortCtrl.sv:207:7
									oRdSop <= (fsmCstate == FSM_RDCMD) && (fsmCstate_d == FSM_IDLE);
							// Trace: src/src/rtl/design/svsrc/PortCtrl.sv:211:3
							always @(posedge iClk or negedge iRst_n)
								// Trace: src/src/rtl/design/svsrc/PortCtrl.sv:212:5
								if (!iRst_n)
									// Trace: src/src/rtl/design/svsrc/PortCtrl.sv:213:7
									oRdEop <= 1'b0;
								else
									// Trace: src/src/rtl/design/svsrc/PortCtrl.sv:215:7
									oRdEop <= (iRdRdy && oRdLast) && oRdVld;
							// Trace: src/src/rtl/design/svsrc/PortCtrl.sv:219:3
							assign tmpRdRdy = (fsmCstate_d == FSM_RDDATA ? iRdRdy : 1'b0);
							// Trace: src/src/rtl/design/svsrc/PortCtrl.sv:220:3
							assign oRdVld = ({fsmCstate_d == FSM_RDDATA} ? tmpRdVld : 1'b0);
							// Trace: src/src/rtl/design/svsrc/PortCtrl.sv:221:3
							assign oRdLast = tmpRdLast & tmpRdVld;
						end
						assign U_PORT_CTRL.iClk = iClk;
						assign U_PORT_CTRL.iRst_n = iRst_n;
						assign oRdSop = U_PORT_CTRL.oRdSop;
						assign oRdEop = U_PORT_CTRL.oRdEop;
						assign oRdVld = U_PORT_CTRL.oRdVld;
						assign oRdData = U_PORT_CTRL.oRdData;
						assign U_PORT_CTRL.iRdRdy = iRdRdy;
						assign oRdLast = U_PORT_CTRL.oRdLast;
					end
					assign U_RD_CHN.iClk = iClk;
					assign U_RD_CHN.iRst_n = iRst_n;
					assign oRdSop[i] = U_RD_CHN.oRdSop;
					assign oRdEop[i] = U_RD_CHN.oRdEop;
					assign oRdVld[i] = U_RD_CHN.oRdVld;
					assign oRdData[(15 - i) * 32+:32] = U_RD_CHN.oRdData;
					assign U_RD_CHN.iRdRdy = iRdRdy[i];
					assign oRdLast[i] = U_RD_CHN.oRdLast;
					assign U_RD_CHN.iWeight = iWeightPld;
					assign U_RD_CHN.iWeightLoad = weightLoadArray[i];
				end
			end
			assign U_RDCTRLTOP16.iClk = iClk;
			assign U_RDCTRLTOP16.iRst_n = iRst_n;
			assign oRdSop = U_RDCTRLTOP16.oRdSop;
			assign oRdEop = U_RDCTRLTOP16.oRdEop;
			assign oRdVld = U_RDCTRLTOP16.oRdVld;
			assign oRdData = U_RDCTRLTOP16.oRdData;
			assign U_RDCTRLTOP16.iRdRdy = iRdRdy;
			assign oRdLast = U_RDCTRLTOP16.oRdLast;
			assign U_RDCTRLTOP16.iWeightPld = iWeightPld;
			assign U_RDCTRLTOP16.iWeightIdx = iWeightIdx;
			assign U_RDCTRLTOP16.iWeightLoad = iWeightLoad;
		end
	endgenerate
	assign U_RD_SCHE_TOP_SV.iClk = iClk;
	assign U_RD_SCHE_TOP_SV.iRst_n = iRst_n;
	assign rdSop = U_RD_SCHE_TOP_SV.oRdSop;
	assign rdEop = U_RD_SCHE_TOP_SV.oRdEop;
	assign rdVld = U_RD_SCHE_TOP_SV.oRdVld;
	assign rdData = U_RD_SCHE_TOP_SV.oRdData;
	assign U_RD_SCHE_TOP_SV.iRdRdy = rdRdy;
	assign rdLast = U_RD_SCHE_TOP_SV.oRdLast;
	assign U_RD_SCHE_TOP_SV.iWeightPld = weightPld;
	assign U_RD_SCHE_TOP_SV.iWeightIdx = iWrrWeightIdx;
	assign U_RD_SCHE_TOP_SV.iWeightLoad = iWrrWeightLoad;
endmodule
