// removed module with interface ports: DcpCrossbarNxN
