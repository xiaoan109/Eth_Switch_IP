************************************************************************
* Cdl Netlist:
*
* Top Cell Name: dpram16x4096
* Configuration: 4096X16CM8
* View Name:     schematic
* Netlist on:    2024-3-29 10:27:320
************************************************************************


************************************************************************
* Library Name: XMC55_DPS
* Created by buildSchLib.pl  at Fri Oct 25 16:34:57 CST 2019
************************************************************************
************************************************************************




************************************************************************
* Library Name: XMC55_DPS
* Cell Name:    xmc55_dps_collar_edge
************************************************************************
.SUBCKT xmc55_dps_collar_edge tie_low vdd vss
** N=75 EP=3 IP=0 FDC=4
M0 tie_low 1 vss vss hvtnfet l=6e-08 w=9e-07 $X=1025 $Y=1120 $D=616
M1 vss 1 tie_low vss hvtnfet l=6e-08 w=9e-07 $X=1285 $Y=1120 $D=616
M2 1 1 vdd vdd hvtpfet l=6e-08 w=9e-07 $X=1025 $Y=2340 $D=636
M3 vdd 1 1 vdd hvtpfet l=6e-08 w=9e-07 $X=1285 $Y=2340 $D=636
.ends

************************************************************************
* Library Name: XMC55_DPS
* Cell Name:    xmc55_dps_collar_corner
************************************************************************
.SUBCKT xmc55_dps_collar_corner aa<12> aa<11> aa<10> aa<9> aa<8> aa<7> aa<6> 
+ aa<5> aa<4> aa<3> aa<2> aa<1> aa<0> aa_int<12> aa_int<11> aa_int<10> 
+ aa_int<9> aa_int<8> aa_int<7> aa_int<6> aa_int<5> aa_int<4> aa_int<3> 
+ aa_int<2> aa_int<1> aa_int<0> ab<12> ab<11> ab<10> ab<9> ab<8> ab<7> ab<6> 
+ ab<5> ab<4> ab<3> ab<2> ab<1> ab<0> ab_int<12> ab_int<11> ab_int<10> 
+ ab_int<9> ab_int<8> ab_int<7> ab_int<6> ab_int<5> ab_int<4> ab_int<3> 
+ ab_int<2> ab_int<1> ab_int<0> cena cena_int cenb cenb_int clka clka_int clkb 
+ clkb_int tie_vdd tie_vss tm<9> tm<8> tm<7> tm<6> tm<5> tm<4> tm<3> tm<2> 
+ tm<1> tm<0> tm_int<9> tm_int<8> tm_int<7> tm_int<6> tm_int<5> tm_int<4> 
+ tm_int<3> tm_int<2> tm_int<1> tm_int<0> vdd vss wena wena_int wenb wenb_int
** N=1833 EP=88 IP=0 FDC=299
D0 vss ab<0> diodenx AREA=7.04e-14 $X=290 $Y=130 $D=2
D1 vss ab<2> diodenx AREA=7.04e-14 $X=2500 $Y=130 $D=2
D2 vss ab<1> diodenx AREA=7.04e-14 $X=2850 $Y=130 $D=2
D3 vss ab<3> diodenx AREA=7.04e-14 $X=3990 $Y=130 $D=2
D4 vss ab<4> diodenx AREA=7.04e-14 $X=4900 $Y=130 $D=2
D5 vss ab<5> diodenx AREA=7.04e-14 $X=6065 $Y=130 $D=2
D6 vss ab<6> diodenx AREA=7.04e-14 $X=6415 $Y=130 $D=2
D7 vss ab<7> diodenx AREA=7.04e-14 $X=7580 $Y=130 $D=2
D8 vss ab<8> diodenx AREA=7.04e-14 $X=8530 $Y=130 $D=2
D9 vss ab<9> diodenx AREA=7.04e-14 $X=9980 $Y=130 $D=2
D10 vss ab<10> diodenx AREA=7.04e-14 $X=10900 $Y=130 $D=2
D11 vss ab<11> diodenx AREA=7.04e-14 $X=11339 $Y=130 $D=2
D12 vss ab<12> diodenx AREA=7.04e-14 $X=11780 $Y=130 $D=2
D13 vss wenb diodenx AREA=7.04e-14 $X=14180 $Y=130 $D=2
D14 vss cenb diodenx AREA=7.04e-14 $X=15100 $Y=130 $D=2
D15 vss clkb diodenx AREA=7.04e-14 $X=16700 $Y=130 $D=2
D16 vss tm<0> diodenx AREA=7.04e-14 $X=17180 $Y=130 $D=2
D17 vss tm<2> diodenx AREA=7.04e-14 $X=18065 $Y=130 $D=2
D18 vss tm<6> diodenx AREA=7.04e-14 $X=18415 $Y=130 $D=2
D19 vss tm<3> diodenx AREA=7.04e-14 $X=19265 $Y=130 $D=2
D20 vss tm<4> diodenx AREA=7.04e-14 $X=19615 $Y=130 $D=2
D21 vss tm<9> diodenx AREA=7.04e-14 $X=23725 $Y=130 $D=2
D22 vss tm<8> diodenx AREA=7.04e-14 $X=24075 $Y=130 $D=2
D23 vss tm<7> diodenx AREA=7.04e-14 $X=24925 $Y=130 $D=2
D24 vss tm<5> diodenx AREA=7.04e-14 $X=25275 $Y=130 $D=2
D25 vss tm<1> diodenx AREA=7.04e-14 $X=26160 $Y=130 $D=2
D26 vss clka diodenx AREA=7.04e-14 $X=26640 $Y=130 $D=2
D27 vss cena diodenx AREA=7.04e-14 $X=28240 $Y=130 $D=2
D28 vss wena diodenx AREA=7.04e-14 $X=29160 $Y=130 $D=2
D29 vss aa<12> diodenx AREA=7.04e-14 $X=31560 $Y=130 $D=2
D30 vss aa<11> diodenx AREA=7.04e-14 $X=32001 $Y=130 $D=2
D31 vss aa<10> diodenx AREA=7.04e-14 $X=32440 $Y=130 $D=2
D32 vss aa<9> diodenx AREA=7.04e-14 $X=33360 $Y=130 $D=2
D33 vss aa<8> diodenx AREA=7.04e-14 $X=34810 $Y=130 $D=2
D34 vss aa<7> diodenx AREA=7.04e-14 $X=35760 $Y=130 $D=2
D35 vss aa<6> diodenx AREA=7.04e-14 $X=36925 $Y=130 $D=2
D36 vss aa<5> diodenx AREA=7.04e-14 $X=37275 $Y=130 $D=2
D37 vss aa<4> diodenx AREA=7.04e-14 $X=38440 $Y=130 $D=2
D38 vss aa<3> diodenx AREA=7.04e-14 $X=39350 $Y=130 $D=2
D39 vss aa<1> diodenx AREA=7.04e-14 $X=40490 $Y=130 $D=2
D40 vss aa<2> diodenx AREA=7.04e-14 $X=40840 $Y=130 $D=2
D41 vss aa<0> diodenx AREA=7.04e-14 $X=43050 $Y=130 $D=2
M42 vss ab<0> 2 vss hvtnfet l=6e-08 w=5e-07 $X=290 $Y=1620 $D=616
M43 ab_int<0> 2 vss vss hvtnfet l=6e-08 w=1e-06 $X=560 $Y=1120 $D=616
M44 vss 2 ab_int<0> vss hvtnfet l=6e-08 w=1e-06 $X=820 $Y=1120 $D=616
M45 ab_int<1> 3 vss vss hvtnfet l=6e-08 w=1e-06 $X=1080 $Y=1120 $D=616
M46 vss 3 ab_int<1> vss hvtnfet l=6e-08 w=1e-06 $X=1340 $Y=1120 $D=616
M47 vss ab<1> 3 vss hvtnfet l=6e-08 w=5e-07 $X=1850 $Y=1620 $D=616
M48 6 ab<2> vss vss hvtnfet l=6e-08 w=5e-07 $X=2110 $Y=1620 $D=616
M49 ab_int<2> 6 vss vss hvtnfet l=6e-08 w=1e-06 $X=2620 $Y=1120 $D=616
M50 vss 6 ab_int<2> vss hvtnfet l=6e-08 w=1e-06 $X=2880 $Y=1120 $D=616
M51 ab_int<3> 7 vss vss hvtnfet l=6e-08 w=1e-06 $X=3140 $Y=1120 $D=616
M52 vss 7 ab_int<3> vss hvtnfet l=6e-08 w=1e-06 $X=3400 $Y=1120 $D=616
M53 vss ab<3> 7 vss hvtnfet l=6e-08 w=5e-07 $X=3910 $Y=1620 $D=616
M54 10 ab<4> vss vss hvtnfet l=6e-08 w=5e-07 $X=4170 $Y=1620 $D=616
M55 ab_int<4> 10 vss vss hvtnfet l=6e-08 w=1e-06 $X=4680 $Y=1120 $D=616
M56 vss 10 ab_int<4> vss hvtnfet l=6e-08 w=1e-06 $X=4940 $Y=1120 $D=616
M57 ab_int<5> 11 vss vss hvtnfet l=6e-08 w=1e-06 $X=5200 $Y=1120 $D=616
M58 vss 11 ab_int<5> vss hvtnfet l=6e-08 w=1e-06 $X=5460 $Y=1120 $D=616
M59 vss ab<5> 11 vss hvtnfet l=6e-08 w=5e-07 $X=5970 $Y=1620 $D=616
M60 14 ab<6> vss vss hvtnfet l=6e-08 w=5e-07 $X=6230 $Y=1620 $D=616
M61 ab_int<6> 14 vss vss hvtnfet l=6e-08 w=1e-06 $X=6740 $Y=1120 $D=616
M62 vss 14 ab_int<6> vss hvtnfet l=6e-08 w=1e-06 $X=7000 $Y=1120 $D=616
M63 ab_int<7> 15 vss vss hvtnfet l=6e-08 w=1e-06 $X=7260 $Y=1120 $D=616
M64 vss 15 ab_int<7> vss hvtnfet l=6e-08 w=1e-06 $X=7520 $Y=1120 $D=616
M65 vss ab<7> 15 vss hvtnfet l=6e-08 w=5e-07 $X=8030 $Y=1620 $D=616
M66 18 ab<8> vss vss hvtnfet l=6e-08 w=5e-07 $X=8290 $Y=1620 $D=616
M67 ab_int<8> 18 vss vss hvtnfet l=6e-08 w=1e-06 $X=8800 $Y=1120 $D=616
M68 vss 18 ab_int<8> vss hvtnfet l=6e-08 w=1e-06 $X=9060 $Y=1120 $D=616
M69 ab_int<9> 19 vss vss hvtnfet l=6e-08 w=1e-06 $X=9320 $Y=1120 $D=616
M70 vss 19 ab_int<9> vss hvtnfet l=6e-08 w=1e-06 $X=9580 $Y=1120 $D=616
M71 vss ab<9> 19 vss hvtnfet l=6e-08 w=5e-07 $X=10090 $Y=1620 $D=616
M72 22 ab<10> vss vss hvtnfet l=6e-08 w=5e-07 $X=10350 $Y=1620 $D=616
M73 ab_int<10> 22 vss vss hvtnfet l=6e-08 w=1e-06 $X=10860 $Y=1120 $D=616
M74 vss 22 ab_int<10> vss hvtnfet l=6e-08 w=1e-06 $X=11120 $Y=1120 $D=616
M75 ab_int<11> 23 vss vss hvtnfet l=6e-08 w=1e-06 $X=11380 $Y=1120 $D=616
M76 vss 23 ab_int<11> vss hvtnfet l=6e-08 w=1e-06 $X=11640 $Y=1120 $D=616
M77 vss ab<11> 23 vss hvtnfet l=6e-08 w=5e-07 $X=12150 $Y=1620 $D=616
M78 26 ab<12> vss vss hvtnfet l=6e-08 w=5e-07 $X=12410 $Y=1620 $D=616
M79 ab_int<12> 26 vss vss hvtnfet l=6e-08 w=1e-06 $X=12920 $Y=1120 $D=616
M80 vss 26 ab_int<12> vss hvtnfet l=6e-08 w=1e-06 $X=13180 $Y=1120 $D=616
M81 wenb_int 27 vss vss hvtnfet l=6e-08 w=1e-06 $X=13440 $Y=1120 $D=616
M82 vss 27 wenb_int vss hvtnfet l=6e-08 w=1e-06 $X=13700 $Y=1120 $D=616
M83 27 wenb vss vss hvtnfet l=6e-08 w=5e-07 $X=13970 $Y=1620 $D=616
M84 105 cenb vss vss hvtnfet l=6e-08 w=3.2e-07 $X=14670 $Y=2067 $D=616
M85 33 31 105 vss hvtnfet l=6e-08 w=3.2e-07 $X=14930 $Y=2067 $D=616
M86 106 32 33 vss hvtnfet l=6e-08 w=2.1e-07 $X=15190 $Y=2177 $D=616
M87 vss clkb 31 vss hvtnfet l=6e-08 w=3.2e-07 $X=15276 $Y=1147 $D=616
M88 vss clkb 106 vss hvtnfet l=6e-08 w=2.1e-07 $X=15450 $Y=2177 $D=616
M89 32 33 vss vss hvtnfet l=6e-08 w=2.1e-07 $X=15710 $Y=2177 $D=616
M90 148 33 vss vss hvtnfet l=6e-08 w=1.5e-06 $X=16220 $Y=1125 $D=616
M91 34 clkb 148 vss hvtnfet l=6e-08 w=1.5e-06 $X=16480 $Y=1125 $D=616
M92 vss 34 clkb_int vss hvtnfet l=6e-08 w=1.15e-06 $X=17250 $Y=1120 $D=616
M93 clkb_int 34 vss vss hvtnfet l=6e-08 w=1.15e-06 $X=17510 $Y=1120 $D=616
M94 vss 34 clkb_int vss hvtnfet l=6e-08 w=1.15e-06 $X=17770 $Y=1120 $D=616
M95 tm_int<0> 35 vss vss hvtnfet l=6e-08 w=1e-06 $X=18030 $Y=1270 $D=616
M96 vss tm<0> 35 vss hvtnfet l=6e-08 w=5e-07 $X=18540 $Y=1620 $D=616
M97 38 tm<2> vss vss hvtnfet l=6e-08 w=5e-07 $X=18800 $Y=1620 $D=616
M98 vss 38 tm_int<2> vss hvtnfet l=6e-08 w=1e-06 $X=19310 $Y=1120 $D=616
M99 tm_int<6> 39 vss vss hvtnfet l=6e-08 w=1e-06 $X=19570 $Y=1120 $D=616
M100 vss tm<6> 39 vss hvtnfet l=6e-08 w=5e-07 $X=20080 $Y=1620 $D=616
M101 42 tm<3> vss vss hvtnfet l=6e-08 w=5e-07 $X=20340 $Y=1620 $D=616
M102 vss 42 tm_int<3> vss hvtnfet l=6e-08 w=1e-06 $X=20850 $Y=1120 $D=616
M103 tm_int<4> 43 vss vss hvtnfet l=6e-08 w=1e-06 $X=21110 $Y=1120 $D=616
M104 vss tm<4> 43 vss hvtnfet l=6e-08 w=5e-07 $X=21620 $Y=1620 $D=616
M105 46 tm<9> vss vss hvtnfet l=6e-08 w=5e-07 $X=21880 $Y=1620 $D=616
M106 vss 46 tm_int<9> vss hvtnfet l=6e-08 w=1e-06 $X=22390 $Y=1120 $D=616
M107 tm_int<8> 47 vss vss hvtnfet l=6e-08 w=1e-06 $X=22650 $Y=1120 $D=616
M108 vss tm<8> 47 vss hvtnfet l=6e-08 w=5e-07 $X=23160 $Y=1620 $D=616
M109 50 tm<7> vss vss hvtnfet l=6e-08 w=5e-07 $X=23420 $Y=1620 $D=616
M110 vss 50 tm_int<7> vss hvtnfet l=6e-08 w=1e-06 $X=23930 $Y=1120 $D=616
M111 tm_int<5> 51 vss vss hvtnfet l=6e-08 w=1e-06 $X=24190 $Y=1120 $D=616
M112 vss tm<5> 51 vss hvtnfet l=6e-08 w=5e-07 $X=24700 $Y=1620 $D=616
M113 54 tm<1> vss vss hvtnfet l=6e-08 w=5e-07 $X=24960 $Y=1620 $D=616
M114 vss 54 tm_int<1> vss hvtnfet l=6e-08 w=1e-06 $X=25470 $Y=1270 $D=616
M115 clka_int 55 vss vss hvtnfet l=6e-08 w=1.15e-06 $X=25730 $Y=1120 $D=616
M116 vss 55 clka_int vss hvtnfet l=6e-08 w=1.15e-06 $X=25990 $Y=1120 $D=616
M117 clka_int 55 vss vss hvtnfet l=6e-08 w=1.15e-06 $X=26250 $Y=1120 $D=616
M118 149 clka 55 vss hvtnfet l=6e-08 w=1.5e-06 $X=27020 $Y=1125 $D=616
M119 vss 57 149 vss hvtnfet l=6e-08 w=1.5e-06 $X=27280 $Y=1125 $D=616
M120 vss 57 58 vss hvtnfet l=6e-08 w=2.1e-07 $X=27790 $Y=2177 $D=616
M121 120 clka vss vss hvtnfet l=6e-08 w=2.1e-07 $X=28050 $Y=2177 $D=616
M122 59 clka vss vss hvtnfet l=6e-08 w=3.2e-07 $X=28224 $Y=1147 $D=616
M123 57 58 120 vss hvtnfet l=6e-08 w=2.1e-07 $X=28310 $Y=2177 $D=616
M124 122 59 57 vss hvtnfet l=6e-08 w=3.2e-07 $X=28570 $Y=2067 $D=616
M125 vss cena 122 vss hvtnfet l=6e-08 w=3.2e-07 $X=28830 $Y=2067 $D=616
M126 vss wena 62 vss hvtnfet l=6e-08 w=5e-07 $X=29530 $Y=1620 $D=616
M127 wena_int 62 vss vss hvtnfet l=6e-08 w=1e-06 $X=29800 $Y=1120 $D=616
M128 vss 62 wena_int vss hvtnfet l=6e-08 w=1e-06 $X=30060 $Y=1120 $D=616
M129 aa_int<12> 63 vss vss hvtnfet l=6e-08 w=1e-06 $X=30320 $Y=1120 $D=616
M130 vss 63 aa_int<12> vss hvtnfet l=6e-08 w=1e-06 $X=30580 $Y=1120 $D=616
M131 vss aa<12> 63 vss hvtnfet l=6e-08 w=5e-07 $X=31090 $Y=1620 $D=616
M132 66 aa<11> vss vss hvtnfet l=6e-08 w=5e-07 $X=31350 $Y=1620 $D=616
M133 aa_int<11> 66 vss vss hvtnfet l=6e-08 w=1e-06 $X=31860 $Y=1120 $D=616
M134 vss 66 aa_int<11> vss hvtnfet l=6e-08 w=1e-06 $X=32120 $Y=1120 $D=616
M135 aa_int<10> 67 vss vss hvtnfet l=6e-08 w=1e-06 $X=32380 $Y=1120 $D=616
M136 vss 67 aa_int<10> vss hvtnfet l=6e-08 w=1e-06 $X=32640 $Y=1120 $D=616
M137 vss aa<10> 67 vss hvtnfet l=6e-08 w=5e-07 $X=33150 $Y=1620 $D=616
M138 70 aa<9> vss vss hvtnfet l=6e-08 w=5e-07 $X=33410 $Y=1620 $D=616
M139 aa_int<9> 70 vss vss hvtnfet l=6e-08 w=1e-06 $X=33920 $Y=1120 $D=616
M140 vss 70 aa_int<9> vss hvtnfet l=6e-08 w=1e-06 $X=34180 $Y=1120 $D=616
M141 aa_int<8> 71 vss vss hvtnfet l=6e-08 w=1e-06 $X=34440 $Y=1120 $D=616
M142 vss 71 aa_int<8> vss hvtnfet l=6e-08 w=1e-06 $X=34700 $Y=1120 $D=616
M143 vss aa<8> 71 vss hvtnfet l=6e-08 w=5e-07 $X=35210 $Y=1620 $D=616
M144 74 aa<7> vss vss hvtnfet l=6e-08 w=5e-07 $X=35470 $Y=1620 $D=616
M145 aa_int<7> 74 vss vss hvtnfet l=6e-08 w=1e-06 $X=35980 $Y=1120 $D=616
M146 vss 74 aa_int<7> vss hvtnfet l=6e-08 w=1e-06 $X=36240 $Y=1120 $D=616
M147 aa_int<6> 75 vss vss hvtnfet l=6e-08 w=1e-06 $X=36500 $Y=1120 $D=616
M148 vss 75 aa_int<6> vss hvtnfet l=6e-08 w=1e-06 $X=36760 $Y=1120 $D=616
M149 vss aa<6> 75 vss hvtnfet l=6e-08 w=5e-07 $X=37270 $Y=1620 $D=616
M150 78 aa<5> vss vss hvtnfet l=6e-08 w=5e-07 $X=37530 $Y=1620 $D=616
M151 aa_int<5> 78 vss vss hvtnfet l=6e-08 w=1e-06 $X=38040 $Y=1120 $D=616
M152 vss 78 aa_int<5> vss hvtnfet l=6e-08 w=1e-06 $X=38300 $Y=1120 $D=616
M153 aa_int<4> 79 vss vss hvtnfet l=6e-08 w=1e-06 $X=38560 $Y=1120 $D=616
M154 vss 79 aa_int<4> vss hvtnfet l=6e-08 w=1e-06 $X=38820 $Y=1120 $D=616
M155 vss aa<4> 79 vss hvtnfet l=6e-08 w=5e-07 $X=39330 $Y=1620 $D=616
M156 82 aa<3> vss vss hvtnfet l=6e-08 w=5e-07 $X=39590 $Y=1620 $D=616
M157 aa_int<3> 82 vss vss hvtnfet l=6e-08 w=1e-06 $X=40100 $Y=1120 $D=616
M158 vss 82 aa_int<3> vss hvtnfet l=6e-08 w=1e-06 $X=40360 $Y=1120 $D=616
M159 aa_int<2> 83 vss vss hvtnfet l=6e-08 w=1e-06 $X=40620 $Y=1120 $D=616
M160 vss 83 aa_int<2> vss hvtnfet l=6e-08 w=1e-06 $X=40880 $Y=1120 $D=616
M161 vss aa<2> 83 vss hvtnfet l=6e-08 w=5e-07 $X=41390 $Y=1620 $D=616
M162 86 aa<1> vss vss hvtnfet l=6e-08 w=5e-07 $X=41650 $Y=1620 $D=616
M163 aa_int<1> 86 vss vss hvtnfet l=6e-08 w=1e-06 $X=42160 $Y=1120 $D=616
M164 vss 86 aa_int<1> vss hvtnfet l=6e-08 w=1e-06 $X=42420 $Y=1120 $D=616
M165 aa_int<0> 87 vss vss hvtnfet l=6e-08 w=1e-06 $X=42680 $Y=1120 $D=616
M166 vss 87 aa_int<0> vss hvtnfet l=6e-08 w=1e-06 $X=42940 $Y=1120 $D=616
M167 87 aa<0> vss vss hvtnfet l=6e-08 w=5e-07 $X=43210 $Y=1620 $D=616
M168 tie_vss tie_vss vss vss hvtnfet l=6e-08 w=2e-07 $X=43750 $Y=1650 $D=616
M169 vss tie_vdd tie_vss vss hvtnfet l=6e-08 w=2e-07 $X=44010 $Y=1650 $D=616
M170 tie_vss tie_vdd cena_int vss hvtnfet l=6e-08 w=2e-07 $X=44520 $Y=1341 $D=616
M171 cenb_int tie_vdd tie_vss vss hvtnfet l=6e-08 w=2e-07 $X=44780 $Y=1341 $D=616
M172 vdd ab<0> 2 vdd hvtpfet l=6e-08 w=1e-06 $X=290 $Y=2440 $D=636
M173 ab_int<0> 2 vdd vdd hvtpfet l=6e-08 w=2e-06 $X=560 $Y=2440 $D=636
M174 vdd 2 ab_int<0> vdd hvtpfet l=6e-08 w=2e-06 $X=820 $Y=2440 $D=636
M175 ab_int<1> 3 vdd vdd hvtpfet l=6e-08 w=2e-06 $X=1080 $Y=2440 $D=636
M176 vdd 3 ab_int<1> vdd hvtpfet l=6e-08 w=2e-06 $X=1340 $Y=2440 $D=636
M177 vdd ab<1> 3 vdd hvtpfet l=6e-08 w=1e-06 $X=1850 $Y=2440 $D=636
M178 6 ab<2> vdd vdd hvtpfet l=6e-08 w=1e-06 $X=2110 $Y=2440 $D=636
M179 ab_int<2> 6 vdd vdd hvtpfet l=6e-08 w=2e-06 $X=2620 $Y=2440 $D=636
M180 vdd 6 ab_int<2> vdd hvtpfet l=6e-08 w=2e-06 $X=2880 $Y=2440 $D=636
M181 ab_int<3> 7 vdd vdd hvtpfet l=6e-08 w=2e-06 $X=3140 $Y=2440 $D=636
M182 vdd 7 ab_int<3> vdd hvtpfet l=6e-08 w=2e-06 $X=3400 $Y=2440 $D=636
M183 vdd ab<3> 7 vdd hvtpfet l=6e-08 w=1e-06 $X=3910 $Y=2440 $D=636
M184 10 ab<4> vdd vdd hvtpfet l=6e-08 w=1e-06 $X=4170 $Y=2440 $D=636
M185 ab_int<4> 10 vdd vdd hvtpfet l=6e-08 w=2e-06 $X=4680 $Y=2440 $D=636
M186 vdd 10 ab_int<4> vdd hvtpfet l=6e-08 w=2e-06 $X=4940 $Y=2440 $D=636
M187 ab_int<5> 11 vdd vdd hvtpfet l=6e-08 w=2e-06 $X=5200 $Y=2440 $D=636
M188 vdd 11 ab_int<5> vdd hvtpfet l=6e-08 w=2e-06 $X=5460 $Y=2440 $D=636
M189 vdd ab<5> 11 vdd hvtpfet l=6e-08 w=1e-06 $X=5970 $Y=2440 $D=636
M190 14 ab<6> vdd vdd hvtpfet l=6e-08 w=1e-06 $X=6230 $Y=2440 $D=636
M191 ab_int<6> 14 vdd vdd hvtpfet l=6e-08 w=2e-06 $X=6740 $Y=2440 $D=636
M192 vdd 14 ab_int<6> vdd hvtpfet l=6e-08 w=2e-06 $X=7000 $Y=2440 $D=636
M193 ab_int<7> 15 vdd vdd hvtpfet l=6e-08 w=2e-06 $X=7260 $Y=2440 $D=636
M194 vdd 15 ab_int<7> vdd hvtpfet l=6e-08 w=2e-06 $X=7520 $Y=2440 $D=636
M195 vdd ab<7> 15 vdd hvtpfet l=6e-08 w=1e-06 $X=8030 $Y=2440 $D=636
M196 18 ab<8> vdd vdd hvtpfet l=6e-08 w=1e-06 $X=8290 $Y=2440 $D=636
M197 ab_int<8> 18 vdd vdd hvtpfet l=6e-08 w=2e-06 $X=8800 $Y=2440 $D=636
M198 vdd 18 ab_int<8> vdd hvtpfet l=6e-08 w=2e-06 $X=9060 $Y=2440 $D=636
M199 ab_int<9> 19 vdd vdd hvtpfet l=6e-08 w=2e-06 $X=9320 $Y=2440 $D=636
M200 vdd 19 ab_int<9> vdd hvtpfet l=6e-08 w=2e-06 $X=9580 $Y=2440 $D=636
M201 vdd ab<9> 19 vdd hvtpfet l=6e-08 w=1e-06 $X=10090 $Y=2440 $D=636
M202 22 ab<10> vdd vdd hvtpfet l=6e-08 w=1e-06 $X=10350 $Y=2440 $D=636
M203 ab_int<10> 22 vdd vdd hvtpfet l=6e-08 w=2e-06 $X=10860 $Y=2440 $D=636
M204 vdd 22 ab_int<10> vdd hvtpfet l=6e-08 w=2e-06 $X=11120 $Y=2440 $D=636
M205 ab_int<11> 23 vdd vdd hvtpfet l=6e-08 w=2e-06 $X=11380 $Y=2440 $D=636
M206 vdd 23 ab_int<11> vdd hvtpfet l=6e-08 w=2e-06 $X=11640 $Y=2440 $D=636
M207 vdd ab<11> 23 vdd hvtpfet l=6e-08 w=1e-06 $X=12150 $Y=2440 $D=636
M208 26 ab<12> vdd vdd hvtpfet l=6e-08 w=1e-06 $X=12410 $Y=2440 $D=636
M209 ab_int<12> 26 vdd vdd hvtpfet l=6e-08 w=2e-06 $X=12920 $Y=2440 $D=636
M210 vdd 26 ab_int<12> vdd hvtpfet l=6e-08 w=2e-06 $X=13180 $Y=2440 $D=636
M211 wenb_int 27 vdd vdd hvtpfet l=6e-08 w=2e-06 $X=13440 $Y=2440 $D=636
M212 vdd 27 wenb_int vdd hvtpfet l=6e-08 w=2e-06 $X=13700 $Y=2440 $D=636
M213 27 wenb vdd vdd hvtpfet l=6e-08 w=1e-06 $X=13970 $Y=2440 $D=636
M214 150 cenb vdd vdd hvtpfet l=6e-08 w=4.8e-07 $X=14670 $Y=3431 $D=636
M215 33 clkb 150 vdd hvtpfet l=6e-08 w=4.8e-07 $X=14930 $Y=3431 $D=636
M216 107 32 33 vdd hvtpfet l=6e-08 w=3.2e-07 $X=15190 $Y=3431 $D=636
M217 vdd clkb 31 vdd hvtpfet l=6e-08 w=4.8e-07 $X=15276 $Y=4410 $D=636
M218 vdd 31 107 vdd hvtpfet l=6e-08 w=3.2e-07 $X=15450 $Y=3431 $D=636
M219 32 33 vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=15710 $Y=3431 $D=636
M220 vdd 33 34 vdd hvtpfet l=6e-08 w=1.5e-06 $X=16220 $Y=3390 $D=636
M221 34 clkb vdd vdd hvtpfet l=6e-08 w=1.5e-06 $X=16480 $Y=3390 $D=636
M222 vdd 34 clkb_int vdd hvtpfet l=6e-08 w=2.3e-06 $X=17250 $Y=2590 $D=636
M223 clkb_int 34 vdd vdd hvtpfet l=6e-08 w=2.3e-06 $X=17510 $Y=2590 $D=636
M224 vdd 34 clkb_int vdd hvtpfet l=6e-08 w=2.3e-06 $X=17770 $Y=2590 $D=636
M225 tm_int<0> 35 vdd vdd hvtpfet l=6e-08 w=2e-06 $X=18030 $Y=2590 $D=636
M226 vdd tm<0> 35 vdd hvtpfet l=6e-08 w=1e-06 $X=18540 $Y=2590 $D=636
M227 38 tm<2> vdd vdd hvtpfet l=6e-08 w=1e-06 $X=18800 $Y=2590 $D=636
M228 vdd 38 tm_int<2> vdd hvtpfet l=6e-08 w=2e-06 $X=19310 $Y=2590 $D=636
M229 tm_int<6> 39 vdd vdd hvtpfet l=6e-08 w=2e-06 $X=19570 $Y=2590 $D=636
M230 vdd tm<6> 39 vdd hvtpfet l=6e-08 w=1e-06 $X=20080 $Y=2590 $D=636
M231 42 tm<3> vdd vdd hvtpfet l=6e-08 w=1e-06 $X=20340 $Y=2590 $D=636
M232 vdd 42 tm_int<3> vdd hvtpfet l=6e-08 w=2e-06 $X=20850 $Y=2590 $D=636
M233 tm_int<4> 43 vdd vdd hvtpfet l=6e-08 w=2e-06 $X=21110 $Y=2590 $D=636
M234 vdd tm<4> 43 vdd hvtpfet l=6e-08 w=1e-06 $X=21620 $Y=2590 $D=636
M235 46 tm<9> vdd vdd hvtpfet l=6e-08 w=1e-06 $X=21880 $Y=2590 $D=636
M236 vdd 46 tm_int<9> vdd hvtpfet l=6e-08 w=2e-06 $X=22390 $Y=2590 $D=636
M237 tm_int<8> 47 vdd vdd hvtpfet l=6e-08 w=2e-06 $X=22650 $Y=2590 $D=636
M238 vdd tm<8> 47 vdd hvtpfet l=6e-08 w=1e-06 $X=23160 $Y=2590 $D=636
M239 50 tm<7> vdd vdd hvtpfet l=6e-08 w=1e-06 $X=23420 $Y=2590 $D=636
M240 vdd 50 tm_int<7> vdd hvtpfet l=6e-08 w=2e-06 $X=23930 $Y=2590 $D=636
M241 tm_int<5> 51 vdd vdd hvtpfet l=6e-08 w=2e-06 $X=24190 $Y=2590 $D=636
M242 vdd tm<5> 51 vdd hvtpfet l=6e-08 w=1e-06 $X=24700 $Y=2590 $D=636
M243 54 tm<1> vdd vdd hvtpfet l=6e-08 w=1e-06 $X=24960 $Y=2590 $D=636
M244 vdd 54 tm_int<1> vdd hvtpfet l=6e-08 w=2e-06 $X=25470 $Y=2590 $D=636
M245 clka_int 55 vdd vdd hvtpfet l=6e-08 w=2.3e-06 $X=25730 $Y=2590 $D=636
M246 vdd 55 clka_int vdd hvtpfet l=6e-08 w=2.3e-06 $X=25990 $Y=2590 $D=636
M247 clka_int 55 vdd vdd hvtpfet l=6e-08 w=2.3e-06 $X=26250 $Y=2590 $D=636
M248 vdd clka 55 vdd hvtpfet l=6e-08 w=1.5e-06 $X=27020 $Y=3390 $D=636
M249 55 57 vdd vdd hvtpfet l=6e-08 w=1.5e-06 $X=27280 $Y=3390 $D=636
M250 vdd 57 58 vdd hvtpfet l=6e-08 w=3.2e-07 $X=27790 $Y=3431 $D=636
M251 121 59 vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=28050 $Y=3431 $D=636
M252 59 clka vdd vdd hvtpfet l=6e-08 w=4.8e-07 $X=28224 $Y=4410 $D=636
M253 57 58 121 vdd hvtpfet l=6e-08 w=3.2e-07 $X=28310 $Y=3431 $D=636
M254 151 clka 57 vdd hvtpfet l=6e-08 w=4.8e-07 $X=28570 $Y=3431 $D=636
M255 vdd cena 151 vdd hvtpfet l=6e-08 w=4.8e-07 $X=28830 $Y=3431 $D=636
M256 vdd wena 62 vdd hvtpfet l=6e-08 w=1e-06 $X=29530 $Y=2440 $D=636
M257 wena_int 62 vdd vdd hvtpfet l=6e-08 w=2e-06 $X=29800 $Y=2440 $D=636
M258 vdd 62 wena_int vdd hvtpfet l=6e-08 w=2e-06 $X=30060 $Y=2440 $D=636
M259 aa_int<12> 63 vdd vdd hvtpfet l=6e-08 w=2e-06 $X=30320 $Y=2440 $D=636
M260 vdd 63 aa_int<12> vdd hvtpfet l=6e-08 w=2e-06 $X=30580 $Y=2440 $D=636
M261 vdd aa<12> 63 vdd hvtpfet l=6e-08 w=1e-06 $X=31090 $Y=2440 $D=636
M262 66 aa<11> vdd vdd hvtpfet l=6e-08 w=1e-06 $X=31350 $Y=2440 $D=636
M263 aa_int<11> 66 vdd vdd hvtpfet l=6e-08 w=2e-06 $X=31860 $Y=2440 $D=636
M264 vdd 66 aa_int<11> vdd hvtpfet l=6e-08 w=2e-06 $X=32120 $Y=2440 $D=636
M265 aa_int<10> 67 vdd vdd hvtpfet l=6e-08 w=2e-06 $X=32380 $Y=2440 $D=636
M266 vdd 67 aa_int<10> vdd hvtpfet l=6e-08 w=2e-06 $X=32640 $Y=2440 $D=636
M267 vdd aa<10> 67 vdd hvtpfet l=6e-08 w=1e-06 $X=33150 $Y=2440 $D=636
M268 70 aa<9> vdd vdd hvtpfet l=6e-08 w=1e-06 $X=33410 $Y=2440 $D=636
M269 aa_int<9> 70 vdd vdd hvtpfet l=6e-08 w=2e-06 $X=33920 $Y=2440 $D=636
M270 vdd 70 aa_int<9> vdd hvtpfet l=6e-08 w=2e-06 $X=34180 $Y=2440 $D=636
M271 aa_int<8> 71 vdd vdd hvtpfet l=6e-08 w=2e-06 $X=34440 $Y=2440 $D=636
M272 vdd 71 aa_int<8> vdd hvtpfet l=6e-08 w=2e-06 $X=34700 $Y=2440 $D=636
M273 vdd aa<8> 71 vdd hvtpfet l=6e-08 w=1e-06 $X=35210 $Y=2440 $D=636
M274 74 aa<7> vdd vdd hvtpfet l=6e-08 w=1e-06 $X=35470 $Y=2440 $D=636
M275 aa_int<7> 74 vdd vdd hvtpfet l=6e-08 w=2e-06 $X=35980 $Y=2440 $D=636
M276 vdd 74 aa_int<7> vdd hvtpfet l=6e-08 w=2e-06 $X=36240 $Y=2440 $D=636
M277 aa_int<6> 75 vdd vdd hvtpfet l=6e-08 w=2e-06 $X=36500 $Y=2440 $D=636
M278 vdd 75 aa_int<6> vdd hvtpfet l=6e-08 w=2e-06 $X=36760 $Y=2440 $D=636
M279 vdd aa<6> 75 vdd hvtpfet l=6e-08 w=1e-06 $X=37270 $Y=2440 $D=636
M280 78 aa<5> vdd vdd hvtpfet l=6e-08 w=1e-06 $X=37530 $Y=2440 $D=636
M281 aa_int<5> 78 vdd vdd hvtpfet l=6e-08 w=2e-06 $X=38040 $Y=2440 $D=636
M282 vdd 78 aa_int<5> vdd hvtpfet l=6e-08 w=2e-06 $X=38300 $Y=2440 $D=636
M283 aa_int<4> 79 vdd vdd hvtpfet l=6e-08 w=2e-06 $X=38560 $Y=2440 $D=636
M284 vdd 79 aa_int<4> vdd hvtpfet l=6e-08 w=2e-06 $X=38820 $Y=2440 $D=636
M285 vdd aa<4> 79 vdd hvtpfet l=6e-08 w=1e-06 $X=39330 $Y=2440 $D=636
M286 82 aa<3> vdd vdd hvtpfet l=6e-08 w=1e-06 $X=39590 $Y=2440 $D=636
M287 aa_int<3> 82 vdd vdd hvtpfet l=6e-08 w=2e-06 $X=40100 $Y=2440 $D=636
M288 vdd 82 aa_int<3> vdd hvtpfet l=6e-08 w=2e-06 $X=40360 $Y=2440 $D=636
M289 aa_int<2> 83 vdd vdd hvtpfet l=6e-08 w=2e-06 $X=40620 $Y=2440 $D=636
M290 vdd 83 aa_int<2> vdd hvtpfet l=6e-08 w=2e-06 $X=40880 $Y=2440 $D=636
M291 vdd aa<2> 83 vdd hvtpfet l=6e-08 w=1e-06 $X=41390 $Y=2440 $D=636
M292 86 aa<1> vdd vdd hvtpfet l=6e-08 w=1e-06 $X=41650 $Y=2440 $D=636
M293 aa_int<1> 86 vdd vdd hvtpfet l=6e-08 w=2e-06 $X=42160 $Y=2440 $D=636
M294 vdd 86 aa_int<1> vdd hvtpfet l=6e-08 w=2e-06 $X=42420 $Y=2440 $D=636
M295 aa_int<0> 87 vdd vdd hvtpfet l=6e-08 w=2e-06 $X=42680 $Y=2440 $D=636
M296 vdd 87 aa_int<0> vdd hvtpfet l=6e-08 w=2e-06 $X=42940 $Y=2440 $D=636
M297 87 aa<0> vdd vdd hvtpfet l=6e-08 w=1e-06 $X=43210 $Y=2440 $D=636
M298 tie_vdd tie_vss vdd vdd hvtpfet l=6e-08 w=2e-07 $X=43750 $Y=2440 $D=636
.ends

************************************************************************
* Library Name: XMC55_DPS
* Cell Name:    xmc55_dps_local_ctrl16
************************************************************************
.SUBCKT xmc55_dps_local_ctrl16 aa<12> aa<11> aa<10> aa<9> aa<8> aa<7> aa<6> 
+ aa<5> aa<4> aa<3> aa<2> aa<1> aa<0> ab<12> ab<11> ab<10> ab<9> ab<8> ab<7> 
+ ab<6> ab<5> ab<4> ab<3> ab<2> ab<1> ab<0> b_pxaa<3> b_pxaa<2> b_pxaa<1> 
+ b_pxaa<0> b_pxab<3> b_pxab<2> b_pxab<1> b_pxab<0> b_pxba_n<7> b_pxba_n<6> 
+ b_pxba_n<5> b_pxba_n<4> b_pxba_n<3> b_pxba_n<2> b_pxba_n<1> b_pxba_n<0> 
+ b_pxbb_n<7> b_pxbb_n<6> b_pxbb_n<5> b_pxbb_n<4> b_pxbb_n<3> b_pxbb_n<2> 
+ b_pxbb_n<1> b_pxbb_n<0> b_pxca_n<7> b_pxca_n<6> b_pxca_n<5> b_pxca_n<4> 
+ b_pxca_n<3> b_pxca_n<2> b_pxca_n<1> b_pxca_n<0> b_pxcb_n<7> b_pxcb_n<6> 
+ b_pxcb_n<5> b_pxcb_n<4> b_pxcb_n<3> b_pxcb_n<2> b_pxcb_n<1> b_pxcb_n<0> cena 
+ cenb clka clkb dbl_pd_n<3> dbl_pd_n<2> dbl_pd_n<1> dbl_pd_n<0> ddqa ddqa_n 
+ ddqb ddqb_n dwla<1> dwla<0> dwlb<1> dwlb<0> l_clk_dqa l_clk_dqa_n l_clk_dqb 
+ l_clk_dqb_n l_lwea l_lweb l_sa_prea_n l_sa_preb_n l_saea_n l_saeb_n lb_ca<3> 
+ lb_ca<2> lb_ca<1> lb_ca<0> lb_cb<3> lb_cb<2> lb_cb<1> lb_cb<0> lb_ma<3> 
+ lb_ma<2> lb_ma<1> lb_ma<0> lb_mb<3> lb_mb<2> lb_mb<1> lb_mb<0> lb_tm_prea_n 
+ lb_tm_preb_n lt_ca<3> lt_ca<2> lt_ca<1> lt_ca<0> lt_cb<3> lt_cb<2> lt_cb<1> 
+ lt_cb<0> lt_ma<3> lt_ma<2> lt_ma<1> lt_ma<0> lt_mb<3> lt_mb<2> lt_mb<1> 
+ lt_mb<0> lt_tm_prea_n lt_tm_preb_n r_clk_dqa r_clk_dqa_n r_clk_dqb 
+ r_clk_dqb_n r_lwea r_lweb r_sa_prea_n r_sa_preb_n r_saea_n r_saeb_n rb_ca<3> 
+ rb_ca<2> rb_ca<1> rb_ca<0> rb_cb<3> rb_cb<2> rb_cb<1> rb_cb<0> rb_ma<3> 
+ rb_ma<2> rb_ma<1> rb_ma<0> rb_mb<3> rb_mb<2> rb_mb<1> rb_mb<0> rb_tm_prea_n 
+ rb_tm_preb_n rt_ca<3> rt_ca<2> rt_ca<1> rt_ca<0> rt_cb<3> rt_cb<2> rt_cb<1> 
+ rt_cb<0> rt_ma<3> rt_ma<2> rt_ma<1> rt_ma<0> rt_mb<3> rt_mb<2> rt_mb<1> 
+ rt_mb<0> rt_tm_prea_n rt_tm_preb_n stclka stclkb t_pxaa<3> t_pxaa<2> 
+ t_pxaa<1> t_pxaa<0> t_pxab<3> t_pxab<2> t_pxab<1> t_pxab<0> t_pxba_n<7> 
+ t_pxba_n<6> t_pxba_n<5> t_pxba_n<4> t_pxba_n<3> t_pxba_n<2> t_pxba_n<1> 
+ t_pxba_n<0> t_pxbb_n<7> t_pxbb_n<6> t_pxbb_n<5> t_pxbb_n<4> t_pxbb_n<3> 
+ t_pxbb_n<2> t_pxbb_n<1> t_pxbb_n<0> t_pxca_n<7> t_pxca_n<6> t_pxca_n<5> 
+ t_pxca_n<4> t_pxca_n<3> t_pxca_n<2> t_pxca_n<1> t_pxca_n<0> t_pxcb_n<7> 
+ t_pxcb_n<6> t_pxcb_n<5> t_pxcb_n<4> t_pxcb_n<3> t_pxcb_n<2> t_pxcb_n<1> 
+ t_pxcb_n<0> tm<9> tm<8> tm<7> tm<6> tm<5> tm<4> tm<3> tm<2> tm<1> tm<0> vdd 
+ vss wena wenb
** N=19585 EP=230 IP=0 FDC=3266
M0 vss 5 15 vss hvtnfet l=6e-08 w=6e-07 $X=965 $Y=37277 $D=616
M1 11 1 vss vss hvtnfet l=6e-08 w=6e-07 $X=1225 $Y=336 $D=616
M2 12 2 vss vss hvtnfet l=6e-08 w=6e-07 $X=1225 $Y=5566 $D=616
M3 13 3 vss vss hvtnfet l=6e-08 w=6e-07 $X=1225 $Y=6796 $D=616
M4 14 4 vss vss hvtnfet l=6e-08 w=6e-07 $X=1225 $Y=12026 $D=616
M5 lb_tm_preb_n 20 vss vss hvtnfet l=6e-08 w=1.287e-06 $X=1225 $Y=13280 $D=616
M6 lt_tm_preb_n 21 vss vss hvtnfet l=6e-08 w=1.287e-06 $X=1225 $Y=20124 $D=616
M7 vss 8 l_clk_dqb vss hvtnfet l=6e-08 w=1.26e-06 $X=1225 $Y=22041 $D=616
M8 vss 9 l_clk_dqb_n vss hvtnfet l=6e-08 w=1.26e-06 $X=1225 $Y=29007 $D=616
M9 l_lweb 10 vss vss hvtnfet l=6e-08 w=1.287e-06 $X=1225 $Y=30897 $D=616
M10 15 5 vss vss hvtnfet l=6e-08 w=6e-07 $X=1225 $Y=37277 $D=616
M11 16 4 vss vss hvtnfet l=6e-08 w=6e-07 $X=1225 $Y=38507 $D=616
M12 17 3 vss vss hvtnfet l=6e-08 w=6e-07 $X=1225 $Y=43737 $D=616
M13 18 6 vss vss hvtnfet l=6e-08 w=6e-07 $X=1225 $Y=44967 $D=616
M14 19 7 vss vss hvtnfet l=6e-08 w=6e-07 $X=1225 $Y=50197 $D=616
M15 vss 20 lb_tm_preb_n vss hvtnfet l=6e-08 w=1.287e-06 $X=1485 $Y=13280 $D=616
M16 vss 21 lt_tm_preb_n vss hvtnfet l=6e-08 w=1.287e-06 $X=1485 $Y=20124 $D=616
M17 l_clk_dqb 8 vss vss hvtnfet l=6e-08 w=1.26e-06 $X=1485 $Y=22041 $D=616
M18 l_clk_dqb_n 9 vss vss hvtnfet l=6e-08 w=1.26e-06 $X=1485 $Y=29007 $D=616
M19 vss 10 l_lweb vss hvtnfet l=6e-08 w=1.287e-06 $X=1485 $Y=30897 $D=616
M20 lb_cb<0> 11 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=1735 $Y=328 $D=616
M21 lb_cb<2> 12 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=1735 $Y=5316 $D=616
M22 lb_mb<0> 13 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=1735 $Y=6788 $D=616
M23 lb_mb<2> 14 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=1735 $Y=11776 $D=616
M24 l_saeb_n 15 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=1735 $Y=37027 $D=616
M25 lt_mb<2> 16 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=1735 $Y=38499 $D=616
M26 lt_mb<0> 17 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=1735 $Y=43487 $D=616
M27 lt_cb<2> 18 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=1735 $Y=44959 $D=616
M28 lt_cb<0> 19 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=1735 $Y=49947 $D=616
M29 vss 8 l_clk_dqb vss hvtnfet l=6e-08 w=1.26e-06 $X=1745 $Y=22041 $D=616
M30 vss 9 l_clk_dqb_n vss hvtnfet l=6e-08 w=1.26e-06 $X=1745 $Y=29007 $D=616
M31 vss 11 lb_cb<0> vss hvtnfet l=6e-08 w=8.58e-07 $X=1995 $Y=328 $D=616
M32 vss 12 lb_cb<2> vss hvtnfet l=6e-08 w=8.58e-07 $X=1995 $Y=5316 $D=616
M33 vss 13 lb_mb<0> vss hvtnfet l=6e-08 w=8.58e-07 $X=1995 $Y=6788 $D=616
M34 vss 14 lb_mb<2> vss hvtnfet l=6e-08 w=8.58e-07 $X=1995 $Y=11776 $D=616
M35 vss 24 20 vss hvtnfet l=6e-08 w=6e-07 $X=1995 $Y=13282 $D=616
M36 vss 25 21 vss hvtnfet l=6e-08 w=6e-07 $X=1995 $Y=20809 $D=616
M37 vss 15 l_saeb_n vss hvtnfet l=6e-08 w=8.58e-07 $X=1995 $Y=37027 $D=616
M38 vss 16 lt_mb<2> vss hvtnfet l=6e-08 w=8.58e-07 $X=1995 $Y=38499 $D=616
M39 vss 17 lt_mb<0> vss hvtnfet l=6e-08 w=8.58e-07 $X=1995 $Y=43487 $D=616
M40 vss 18 lt_cb<2> vss hvtnfet l=6e-08 w=8.58e-07 $X=1995 $Y=44959 $D=616
M41 vss 19 lt_cb<0> vss hvtnfet l=6e-08 w=8.58e-07 $X=1995 $Y=49947 $D=616
M42 8 clkb vss vss hvtnfet l=6e-08 w=1.05e-06 $X=2005 $Y=22251 $D=616
M43 9 23 vss vss hvtnfet l=6e-08 w=1.05e-06 $X=2005 $Y=29007 $D=616
M44 lb_cb<0> 11 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=2255 $Y=328 $D=616
M45 lb_cb<2> 12 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=2255 $Y=5316 $D=616
M46 lb_mb<0> 13 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=2255 $Y=6788 $D=616
M47 lb_mb<2> 14 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=2255 $Y=11776 $D=616
M48 l_saeb_n 15 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=2255 $Y=37027 $D=616
M49 lt_mb<2> 16 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=2255 $Y=38499 $D=616
M50 lt_mb<0> 17 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=2255 $Y=43487 $D=616
M51 lt_cb<2> 18 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=2255 $Y=44959 $D=616
M52 lt_cb<0> 19 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=2255 $Y=49947 $D=616
M53 vss 15 l_saeb_n vss hvtnfet l=6e-08 w=8.58e-07 $X=2515 $Y=37027 $D=616
M54 vss 34 lb_cb<1> vss hvtnfet l=6e-08 w=8.58e-07 $X=2765 $Y=328 $D=616
M55 vss 35 lb_cb<3> vss hvtnfet l=6e-08 w=8.58e-07 $X=2765 $Y=5316 $D=616
M56 vss 36 lb_mb<1> vss hvtnfet l=6e-08 w=8.58e-07 $X=2765 $Y=6788 $D=616
M57 vss 37 lb_mb<3> vss hvtnfet l=6e-08 w=8.58e-07 $X=2765 $Y=11776 $D=616
M58 vss 39 lt_mb<3> vss hvtnfet l=6e-08 w=8.58e-07 $X=2765 $Y=38499 $D=616
M59 vss 40 lt_mb<1> vss hvtnfet l=6e-08 w=8.58e-07 $X=2765 $Y=43487 $D=616
M60 vss 41 lt_cb<3> vss hvtnfet l=6e-08 w=8.58e-07 $X=2765 $Y=44959 $D=616
M61 vss 42 lt_cb<1> vss hvtnfet l=6e-08 w=8.58e-07 $X=2765 $Y=49947 $D=616
M62 l_saeb_n 15 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=2775 $Y=37027 $D=616
M63 909 26 vss vss hvtnfet l=6e-08 w=1.8e-07 $X=2821 $Y=17143 $D=616
M64 26 28 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=2821 $Y=17812 $D=616
M65 4 29 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=2821 $Y=18983 $D=616
M66 910 4 vss vss hvtnfet l=6e-08 w=1.8e-07 $X=2821 $Y=19609 $D=616
M67 911 27 vss vss hvtnfet l=6e-08 w=1.8e-07 $X=2821 $Y=24063 $D=616
M68 27 30 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=2821 $Y=24732 $D=616
M69 3 31 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=2821 $Y=25903 $D=616
M70 912 3 vss vss hvtnfet l=6e-08 w=1.8e-07 $X=2821 $Y=26529 $D=616
M71 lb_cb<1> 34 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=3025 $Y=328 $D=616
M72 lb_cb<3> 35 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=3025 $Y=5316 $D=616
M73 lb_mb<1> 36 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=3025 $Y=6788 $D=616
M74 lb_mb<3> 37 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=3025 $Y=11776 $D=616
M75 lt_mb<3> 39 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=3025 $Y=38499 $D=616
M76 lt_mb<1> 40 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=3025 $Y=43487 $D=616
M77 lt_cb<3> 41 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=3025 $Y=44959 $D=616
M78 lt_cb<1> 42 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=3025 $Y=49947 $D=616
M79 28 33 909 vss hvtnfet l=6e-08 w=1.8e-07 $X=3081 $Y=17143 $D=616
M80 vss 28 26 vss hvtnfet l=6e-08 w=1.37e-07 $X=3081 $Y=17812 $D=616
M81 vss 29 4 vss hvtnfet l=6e-08 w=1.37e-07 $X=3081 $Y=18983 $D=616
M82 29 33 910 vss hvtnfet l=6e-08 w=1.8e-07 $X=3081 $Y=19609 $D=616
M83 30 33 911 vss hvtnfet l=6e-08 w=1.8e-07 $X=3081 $Y=24063 $D=616
M84 vss 30 27 vss hvtnfet l=6e-08 w=1.37e-07 $X=3081 $Y=24732 $D=616
M85 vss 31 3 vss hvtnfet l=6e-08 w=1.37e-07 $X=3081 $Y=25903 $D=616
M86 31 33 912 vss hvtnfet l=6e-08 w=1.8e-07 $X=3081 $Y=26529 $D=616
M87 vss 34 lb_cb<1> vss hvtnfet l=6e-08 w=8.58e-07 $X=3285 $Y=328 $D=616
M88 vss 35 lb_cb<3> vss hvtnfet l=6e-08 w=8.58e-07 $X=3285 $Y=5316 $D=616
M89 vss 36 lb_mb<1> vss hvtnfet l=6e-08 w=8.58e-07 $X=3285 $Y=6788 $D=616
M90 vss 37 lb_mb<3> vss hvtnfet l=6e-08 w=8.58e-07 $X=3285 $Y=11776 $D=616
M91 vss 51 l_sa_preb_n vss hvtnfet l=6e-08 w=8.58e-07 $X=3285 $Y=37027 $D=616
M92 vss 39 lt_mb<3> vss hvtnfet l=6e-08 w=8.58e-07 $X=3285 $Y=38499 $D=616
M93 vss 40 lt_mb<1> vss hvtnfet l=6e-08 w=8.58e-07 $X=3285 $Y=43487 $D=616
M94 vss 41 lt_cb<3> vss hvtnfet l=6e-08 w=8.58e-07 $X=3285 $Y=44959 $D=616
M95 vss 42 lt_cb<1> vss hvtnfet l=6e-08 w=8.58e-07 $X=3285 $Y=49947 $D=616
M96 vss ab<2> 44 vss hvtnfet l=6e-08 w=2.74e-07 $X=3396 $Y=13476 $D=616
M97 l_sa_preb_n 51 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=3545 $Y=37027 $D=616
M98 913 43 vss vss hvtnfet l=6e-08 w=8.23e-07 $X=3591 $Y=17143 $D=616
M99 914 43 vss vss hvtnfet l=6e-08 w=8.23e-07 $X=3591 $Y=18966 $D=616
M100 915 43 vss vss hvtnfet l=6e-08 w=8.23e-07 $X=3591 $Y=24063 $D=616
M101 916 43 vss vss hvtnfet l=6e-08 w=8.23e-07 $X=3591 $Y=25886 $D=616
M102 52 stclkb vss vss hvtnfet l=6e-08 w=2.74e-07 $X=3705 $Y=30668 $D=616
M103 vss 47 34 vss hvtnfet l=6e-08 w=6e-07 $X=3795 $Y=336 $D=616
M104 vss 48 35 vss hvtnfet l=6e-08 w=6e-07 $X=3795 $Y=5566 $D=616
M105 vss 27 36 vss hvtnfet l=6e-08 w=6e-07 $X=3795 $Y=6796 $D=616
M106 vss 26 37 vss hvtnfet l=6e-08 w=6e-07 $X=3795 $Y=12026 $D=616
M107 vss 26 39 vss hvtnfet l=6e-08 w=6e-07 $X=3795 $Y=38507 $D=616
M108 vss 27 40 vss hvtnfet l=6e-08 w=6e-07 $X=3795 $Y=43737 $D=616
M109 vss 49 41 vss hvtnfet l=6e-08 w=6e-07 $X=3795 $Y=44967 $D=616
M110 vss 50 42 vss hvtnfet l=6e-08 w=6e-07 $X=3795 $Y=50197 $D=616
M111 vss 51 l_sa_preb_n vss hvtnfet l=6e-08 w=8.58e-07 $X=3805 $Y=37027 $D=616
M112 917 45 913 vss hvtnfet l=6e-08 w=5.49e-07 $X=3861 $Y=17143 $D=616
M113 918 45 914 vss hvtnfet l=6e-08 w=5.49e-07 $X=3861 $Y=19240 $D=616
M114 919 46 915 vss hvtnfet l=6e-08 w=5.49e-07 $X=3861 $Y=24063 $D=616
M115 920 46 916 vss hvtnfet l=6e-08 w=5.49e-07 $X=3861 $Y=26160 $D=616
M116 53 44 vss vss hvtnfet l=6e-08 w=2.74e-07 $X=3906 $Y=13476 $D=616
M117 vss clkb 43 vss hvtnfet l=6e-08 w=6e-07 $X=4066 $Y=32403 $D=616
M118 28 53 917 vss hvtnfet l=6e-08 w=5.49e-07 $X=4121 $Y=17143 $D=616
M119 29 44 918 vss hvtnfet l=6e-08 w=5.49e-07 $X=4121 $Y=19240 $D=616
M120 30 53 919 vss hvtnfet l=6e-08 w=5.49e-07 $X=4121 $Y=24063 $D=616
M121 31 44 920 vss hvtnfet l=6e-08 w=5.49e-07 $X=4121 $Y=26160 $D=616
M122 vss 52 59 vss hvtnfet l=6e-08 w=5.49e-07 $X=4215 $Y=30668 $D=616
M123 vss 55 51 vss hvtnfet l=6e-08 w=6e-07 $X=4315 $Y=37277 $D=616
M124 43 clkb vss vss hvtnfet l=6e-08 w=6e-07 $X=4326 $Y=32403 $D=616
M125 vss ab<3> 46 vss hvtnfet l=6e-08 w=2.74e-07 $X=4416 $Y=13476 $D=616
M126 59 56 vss vss hvtnfet l=6e-08 w=5.49e-07 $X=4475 $Y=30668 $D=616
M127 b_pxab<0> 60 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=4550 $Y=336 $D=616
M128 60 61 vss vss hvtnfet l=6e-08 w=5e-07 $X=4550 $Y=6701 $D=616
M129 61 62 vss vss hvtnfet l=6e-08 w=3e-07 $X=4550 $Y=7831 $D=616
M130 921 57 vss vss hvtnfet l=6e-08 w=4.11e-07 $X=4550 $Y=11276 $D=616
M131 922 57 vss vss hvtnfet l=6e-08 w=4.11e-07 $X=4550 $Y=39446 $D=616
M132 64 63 vss vss hvtnfet l=6e-08 w=3e-07 $X=4550 $Y=43002 $D=616
M133 65 64 vss vss hvtnfet l=6e-08 w=5e-07 $X=4550 $Y=43932 $D=616
M134 t_pxab<0> 65 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=4550 $Y=49512 $D=616
M135 vss 60 b_pxab<0> vss hvtnfet l=6e-08 w=1.285e-06 $X=4810 $Y=336 $D=616
M136 vss 61 60 vss hvtnfet l=6e-08 w=5e-07 $X=4810 $Y=6701 $D=616
M137 vss 62 61 vss hvtnfet l=6e-08 w=3e-07 $X=4810 $Y=7831 $D=616
M138 62 24 921 vss hvtnfet l=6e-08 w=4.11e-07 $X=4810 $Y=11276 $D=616
M139 63 25 922 vss hvtnfet l=6e-08 w=4.11e-07 $X=4810 $Y=39446 $D=616
M140 vss 63 64 vss hvtnfet l=6e-08 w=3e-07 $X=4810 $Y=43002 $D=616
M141 vss 64 65 vss hvtnfet l=6e-08 w=5e-07 $X=4810 $Y=43932 $D=616
M142 vss 65 t_pxab<0> vss hvtnfet l=6e-08 w=1.285e-06 $X=4810 $Y=49512 $D=616
M143 45 46 vss vss hvtnfet l=6e-08 w=2.74e-07 $X=4926 $Y=13476 $D=616
M144 vss 66 586 vss hvtnfet l=1.4e-07 w=3.2e-07 $X=4939 $Y=37127 $D=616
M145 vss 59 56 vss hvtnfet l=6e-08 w=5.49e-07 $X=4985 $Y=30668 $D=616
M146 vss 58 587 vss hvtnfet l=6e-08 w=3.2e-07 $X=5069 $Y=32828 $D=616
M147 923 67 vss vss hvtnfet l=6e-08 w=1.8e-07 $X=5141 $Y=17143 $D=616
M148 67 73 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=5141 $Y=17812 $D=616
M149 68 74 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=5141 $Y=18983 $D=616
M150 924 68 vss vss hvtnfet l=6e-08 w=1.8e-07 $X=5141 $Y=19609 $D=616
M151 925 69 vss vss hvtnfet l=6e-08 w=1.8e-07 $X=5141 $Y=24063 $D=616
M152 69 75 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=5141 $Y=24732 $D=616
M153 57 76 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=5141 $Y=25903 $D=616
M154 926 57 vss vss hvtnfet l=6e-08 w=1.8e-07 $X=5141 $Y=26529 $D=616
M155 56 70 vss vss hvtnfet l=6e-08 w=5.49e-07 $X=5245 $Y=30668 $D=616
M156 66 71 vss vss hvtnfet l=1.4e-07 w=3.2e-07 $X=5279 $Y=37127 $D=616
M157 b_pxab<1> 78 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=5320 $Y=336 $D=616
M158 78 79 vss vss hvtnfet l=6e-08 w=5e-07 $X=5320 $Y=6701 $D=616
M159 79 80 vss vss hvtnfet l=6e-08 w=3e-07 $X=5320 $Y=7831 $D=616
M160 927 24 80 vss hvtnfet l=6e-08 w=4.11e-07 $X=5320 $Y=11276 $D=616
M161 928 25 81 vss hvtnfet l=6e-08 w=4.11e-07 $X=5320 $Y=39446 $D=616
M162 82 81 vss vss hvtnfet l=6e-08 w=3e-07 $X=5320 $Y=43002 $D=616
M163 83 82 vss vss hvtnfet l=6e-08 w=5e-07 $X=5320 $Y=43932 $D=616
M164 t_pxab<1> 83 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=5320 $Y=49512 $D=616
M165 73 33 923 vss hvtnfet l=6e-08 w=1.8e-07 $X=5401 $Y=17143 $D=616
M166 vss 73 67 vss hvtnfet l=6e-08 w=1.37e-07 $X=5401 $Y=17812 $D=616
M167 vss 74 68 vss hvtnfet l=6e-08 w=1.37e-07 $X=5401 $Y=18983 $D=616
M168 74 33 924 vss hvtnfet l=6e-08 w=1.8e-07 $X=5401 $Y=19609 $D=616
M169 75 33 925 vss hvtnfet l=6e-08 w=1.8e-07 $X=5401 $Y=24063 $D=616
M170 vss 75 69 vss hvtnfet l=6e-08 w=1.37e-07 $X=5401 $Y=24732 $D=616
M171 vss 76 57 vss hvtnfet l=6e-08 w=1.37e-07 $X=5401 $Y=25903 $D=616
M172 76 33 926 vss hvtnfet l=6e-08 w=1.8e-07 $X=5401 $Y=26529 $D=616
M173 929 72 vss vss hvtnfet l=6e-08 w=6.4e-07 $X=5579 $Y=32508 $D=616
M174 vss 78 b_pxab<1> vss hvtnfet l=6e-08 w=1.285e-06 $X=5580 $Y=336 $D=616
M175 vss 79 78 vss hvtnfet l=6e-08 w=5e-07 $X=5580 $Y=6701 $D=616
M176 vss 80 79 vss hvtnfet l=6e-08 w=3e-07 $X=5580 $Y=7831 $D=616
M177 vss 69 927 vss hvtnfet l=6e-08 w=4.11e-07 $X=5580 $Y=11276 $D=616
M178 vss 69 928 vss hvtnfet l=6e-08 w=4.11e-07 $X=5580 $Y=39446 $D=616
M179 vss 81 82 vss hvtnfet l=6e-08 w=3e-07 $X=5580 $Y=43002 $D=616
M180 vss 82 83 vss hvtnfet l=6e-08 w=5e-07 $X=5580 $Y=43932 $D=616
M181 vss 83 t_pxab<1> vss hvtnfet l=6e-08 w=1.285e-06 $X=5580 $Y=49512 $D=616
M182 vss ab<5> 86 vss hvtnfet l=6e-08 w=2.74e-07 $X=5716 $Y=13476 $D=616
M183 5 85 929 vss hvtnfet l=6e-08 w=6.4e-07 $X=5839 $Y=32508 $D=616
M184 930 43 vss vss hvtnfet l=6e-08 w=8.23e-07 $X=5911 $Y=17143 $D=616
M185 931 43 vss vss hvtnfet l=6e-08 w=8.23e-07 $X=5911 $Y=18966 $D=616
M186 932 43 vss vss hvtnfet l=6e-08 w=8.23e-07 $X=5911 $Y=24063 $D=616
M187 933 43 vss vss hvtnfet l=6e-08 w=8.23e-07 $X=5911 $Y=25886 $D=616
M188 70 clkb vss vss hvtnfet l=6e-08 w=6e-07 $X=6015 $Y=30668 $D=616
M189 vss ddqb 71 vss hvtnfet l=6e-08 w=2.4e-07 $X=6079 $Y=37292 $D=616
M190 b_pxab<2> 90 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=6090 $Y=336 $D=616
M191 90 91 vss vss hvtnfet l=6e-08 w=5e-07 $X=6090 $Y=6701 $D=616
M192 91 92 vss vss hvtnfet l=6e-08 w=3e-07 $X=6090 $Y=7831 $D=616
M193 934 68 vss vss hvtnfet l=6e-08 w=4.11e-07 $X=6090 $Y=11276 $D=616
M194 935 68 vss vss hvtnfet l=6e-08 w=4.11e-07 $X=6090 $Y=39446 $D=616
M195 94 93 vss vss hvtnfet l=6e-08 w=3e-07 $X=6090 $Y=43002 $D=616
M196 95 94 vss vss hvtnfet l=6e-08 w=5e-07 $X=6090 $Y=43932 $D=616
M197 t_pxab<2> 95 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=6090 $Y=49512 $D=616
M198 936 87 930 vss hvtnfet l=6e-08 w=5.49e-07 $X=6181 $Y=17143 $D=616
M199 937 87 931 vss hvtnfet l=6e-08 w=5.49e-07 $X=6181 $Y=19240 $D=616
M200 938 88 932 vss hvtnfet l=6e-08 w=5.49e-07 $X=6181 $Y=24063 $D=616
M201 939 88 933 vss hvtnfet l=6e-08 w=5.49e-07 $X=6181 $Y=26160 $D=616
M202 97 86 vss vss hvtnfet l=6e-08 w=2.74e-07 $X=6226 $Y=13476 $D=616
M203 71 ddqb_n vss vss hvtnfet l=6e-08 w=2.4e-07 $X=6339 $Y=37292 $D=616
M204 vss 90 b_pxab<2> vss hvtnfet l=6e-08 w=1.285e-06 $X=6350 $Y=336 $D=616
M205 vss 91 90 vss hvtnfet l=6e-08 w=5e-07 $X=6350 $Y=6701 $D=616
M206 vss 92 91 vss hvtnfet l=6e-08 w=3e-07 $X=6350 $Y=7831 $D=616
M207 92 24 934 vss hvtnfet l=6e-08 w=4.11e-07 $X=6350 $Y=11276 $D=616
M208 93 25 935 vss hvtnfet l=6e-08 w=4.11e-07 $X=6350 $Y=39446 $D=616
M209 vss 93 94 vss hvtnfet l=6e-08 w=3e-07 $X=6350 $Y=43002 $D=616
M210 vss 94 95 vss hvtnfet l=6e-08 w=5e-07 $X=6350 $Y=43932 $D=616
M211 vss 95 t_pxab<2> vss hvtnfet l=6e-08 w=1.285e-06 $X=6350 $Y=49512 $D=616
M212 73 97 936 vss hvtnfet l=6e-08 w=5.49e-07 $X=6441 $Y=17143 $D=616
M213 74 86 937 vss hvtnfet l=6e-08 w=5.49e-07 $X=6441 $Y=19240 $D=616
M214 75 97 938 vss hvtnfet l=6e-08 w=5.49e-07 $X=6441 $Y=24063 $D=616
M215 76 86 939 vss hvtnfet l=6e-08 w=5.49e-07 $X=6441 $Y=26160 $D=616
M216 85 89 vss vss hvtnfet l=6e-08 w=3.2e-07 $X=6524 $Y=32828 $D=616
M217 142 clkb 595 vss hvtnfet l=6e-08 w=8e-07 $X=6525 $Y=30668 $D=616
M218 vss ab<6> 88 vss hvtnfet l=6e-08 w=2.74e-07 $X=6736 $Y=13476 $D=616
M219 595 clkb 142 vss hvtnfet l=6e-08 w=8e-07 $X=6785 $Y=30668 $D=616
M220 b_pxab<3> 99 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=6860 $Y=336 $D=616
M221 99 100 vss vss hvtnfet l=6e-08 w=5e-07 $X=6860 $Y=6701 $D=616
M222 100 101 vss vss hvtnfet l=6e-08 w=3e-07 $X=6860 $Y=7831 $D=616
M223 940 24 101 vss hvtnfet l=6e-08 w=4.11e-07 $X=6860 $Y=11276 $D=616
M224 941 25 102 vss hvtnfet l=6e-08 w=4.11e-07 $X=6860 $Y=39446 $D=616
M225 103 102 vss vss hvtnfet l=6e-08 w=3e-07 $X=6860 $Y=43002 $D=616
M226 104 103 vss vss hvtnfet l=6e-08 w=5e-07 $X=6860 $Y=43932 $D=616
M227 t_pxab<3> 104 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=6860 $Y=49512 $D=616
M228 109 85 vss vss hvtnfet l=6e-08 w=3.2e-07 $X=7034 $Y=32828 $D=616
M229 89 58 vss vss hvtnfet l=6e-08 w=3.2e-07 $X=7069 $Y=37292 $D=616
M230 vss 99 b_pxab<3> vss hvtnfet l=6e-08 w=1.285e-06 $X=7120 $Y=336 $D=616
M231 vss 100 99 vss hvtnfet l=6e-08 w=5e-07 $X=7120 $Y=6701 $D=616
M232 vss 101 100 vss hvtnfet l=6e-08 w=3e-07 $X=7120 $Y=7831 $D=616
M233 vss 67 940 vss hvtnfet l=6e-08 w=4.11e-07 $X=7120 $Y=11276 $D=616
M234 vss 67 941 vss hvtnfet l=6e-08 w=4.11e-07 $X=7120 $Y=39446 $D=616
M235 vss 102 103 vss hvtnfet l=6e-08 w=3e-07 $X=7120 $Y=43002 $D=616
M236 vss 103 104 vss hvtnfet l=6e-08 w=5e-07 $X=7120 $Y=43932 $D=616
M237 vss 104 t_pxab<3> vss hvtnfet l=6e-08 w=1.285e-06 $X=7120 $Y=49512 $D=616
M238 87 88 vss vss hvtnfet l=6e-08 w=2.74e-07 $X=7246 $Y=13476 $D=616
M239 595 59 vss vss hvtnfet l=6e-08 w=8e-07 $X=7295 $Y=30668 $D=616
M240 942 105 vss vss hvtnfet l=6e-08 w=1.8e-07 $X=7461 $Y=17143 $D=616
M241 943 106 vss vss hvtnfet l=6e-08 w=1.8e-07 $X=7461 $Y=19609 $D=616
M242 944 107 vss vss hvtnfet l=6e-08 w=1.8e-07 $X=7461 $Y=24063 $D=616
M243 945 108 vss vss hvtnfet l=6e-08 w=1.8e-07 $X=7461 $Y=26529 $D=616
M244 105 111 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=7476 $Y=17812 $D=616
M245 106 112 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=7476 $Y=18983 $D=616
M246 107 113 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=7476 $Y=24732 $D=616
M247 108 114 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=7476 $Y=25903 $D=616
M248 vss 59 595 vss hvtnfet l=6e-08 w=8e-07 $X=7555 $Y=30668 $D=616
M249 vss 110 89 vss hvtnfet l=1.2e-07 w=1.5e-07 $X=7579 $Y=37297 $D=616
M250 vss 109 119 vss hvtnfet l=2.5e-07 w=3.5e-07 $X=7604 $Y=32613 $D=616
M251 b_pxbb_n<0> 115 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=7630 $Y=336 $D=616
M252 115 116 vss vss hvtnfet l=6e-08 w=5e-07 $X=7630 $Y=6701 $D=616
M253 116 107 vss vss hvtnfet l=6e-08 w=3e-07 $X=7630 $Y=7831 $D=616
M254 117 107 vss vss hvtnfet l=6e-08 w=3e-07 $X=7630 $Y=43002 $D=616
M255 118 117 vss vss hvtnfet l=6e-08 w=5e-07 $X=7630 $Y=43932 $D=616
M256 t_pxbb_n<0> 118 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=7630 $Y=49512 $D=616
M257 111 33 942 vss hvtnfet l=6e-08 w=1.8e-07 $X=7721 $Y=17143 $D=616
M258 112 33 943 vss hvtnfet l=6e-08 w=1.8e-07 $X=7721 $Y=19609 $D=616
M259 113 33 944 vss hvtnfet l=6e-08 w=1.8e-07 $X=7721 $Y=24063 $D=616
M260 114 33 945 vss hvtnfet l=6e-08 w=1.8e-07 $X=7721 $Y=26529 $D=616
M261 vss 111 105 vss hvtnfet l=6e-08 w=1.37e-07 $X=7736 $Y=17812 $D=616
M262 vss 112 106 vss hvtnfet l=6e-08 w=1.37e-07 $X=7736 $Y=18983 $D=616
M263 vss 113 107 vss hvtnfet l=6e-08 w=1.37e-07 $X=7736 $Y=24732 $D=616
M264 vss 114 108 vss hvtnfet l=6e-08 w=1.37e-07 $X=7736 $Y=25903 $D=616
M265 vss 115 b_pxbb_n<0> vss hvtnfet l=6e-08 w=1.285e-06 $X=7890 $Y=336 $D=616
M266 vss 116 115 vss hvtnfet l=6e-08 w=5e-07 $X=7890 $Y=6701 $D=616
M267 vss 107 116 vss hvtnfet l=6e-08 w=3e-07 $X=7890 $Y=7831 $D=616
M268 vss 107 117 vss hvtnfet l=6e-08 w=3e-07 $X=7890 $Y=43002 $D=616
M269 vss 117 118 vss hvtnfet l=6e-08 w=5e-07 $X=7890 $Y=43932 $D=616
M270 vss 118 t_pxbb_n<0> vss hvtnfet l=6e-08 w=1.285e-06 $X=7890 $Y=49512 $D=616
M271 120 119 vss vss hvtnfet l=6e-08 w=3.5e-07 $X=8054 $Y=32613 $D=616
M272 110 89 vss vss hvtnfet l=6e-08 w=3e-07 $X=8149 $Y=37257 $D=616
M273 946 43 vss vss hvtnfet l=6e-08 w=8.23e-07 $X=8231 $Y=17143 $D=616
M274 947 43 vss vss hvtnfet l=6e-08 w=8.23e-07 $X=8231 $Y=18966 $D=616
M275 948 43 vss vss hvtnfet l=6e-08 w=8.23e-07 $X=8231 $Y=24063 $D=616
M276 949 43 vss vss hvtnfet l=6e-08 w=8.23e-07 $X=8231 $Y=25886 $D=616
M277 b_pxbb_n<1> 125 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=8400 $Y=336 $D=616
M278 125 126 vss vss hvtnfet l=6e-08 w=5e-07 $X=8400 $Y=6701 $D=616
M279 126 108 vss vss hvtnfet l=6e-08 w=3e-07 $X=8400 $Y=7831 $D=616
M280 127 108 vss vss hvtnfet l=6e-08 w=3e-07 $X=8400 $Y=43002 $D=616
M281 128 127 vss vss hvtnfet l=6e-08 w=5e-07 $X=8400 $Y=43932 $D=616
M282 t_pxbb_n<1> 128 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=8400 $Y=49512 $D=616
M283 vss 122 121 vss hvtnfet l=6e-08 w=2.74e-07 $X=8466 $Y=13476 $D=616
M284 950 121 946 vss hvtnfet l=6e-08 w=5.49e-07 $X=8501 $Y=17417 $D=616
M285 951 121 947 vss hvtnfet l=6e-08 w=5.49e-07 $X=8501 $Y=18966 $D=616
M286 952 122 948 vss hvtnfet l=6e-08 w=5.49e-07 $X=8501 $Y=24337 $D=616
M287 953 122 949 vss hvtnfet l=6e-08 w=5.49e-07 $X=8501 $Y=25886 $D=616
M288 123 123 vss vss hvtnfet l=6e-08 w=2e-07 $X=8594 $Y=11546 $D=616
M289 954 120 55 vss hvtnfet l=6e-08 w=6.4e-07 $X=8619 $Y=32508 $D=616
M290 dwlb<0> 124 vss vss hvtnfet l=6e-08 w=3e-07 $X=8659 $Y=31098 $D=616
M291 25 124 vss vss hvtnfet l=6e-08 w=3e-07 $X=8659 $Y=37457 $D=616
M292 vss 125 b_pxbb_n<1> vss hvtnfet l=6e-08 w=1.285e-06 $X=8660 $Y=336 $D=616
M293 vss 126 125 vss hvtnfet l=6e-08 w=5e-07 $X=8660 $Y=6701 $D=616
M294 vss 108 126 vss hvtnfet l=6e-08 w=3e-07 $X=8660 $Y=7831 $D=616
M295 vss 108 127 vss hvtnfet l=6e-08 w=3e-07 $X=8660 $Y=43002 $D=616
M296 vss 127 128 vss hvtnfet l=6e-08 w=5e-07 $X=8660 $Y=43932 $D=616
M297 vss 128 t_pxbb_n<1> vss hvtnfet l=6e-08 w=1.285e-06 $X=8660 $Y=49512 $D=616
M298 955 129 950 vss hvtnfet l=6e-08 w=5.49e-07 $X=8761 $Y=17417 $D=616
M299 956 129 951 vss hvtnfet l=6e-08 w=5.49e-07 $X=8761 $Y=18966 $D=616
M300 957 129 952 vss hvtnfet l=6e-08 w=5.49e-07 $X=8761 $Y=24337 $D=616
M301 958 129 953 vss hvtnfet l=6e-08 w=5.49e-07 $X=8761 $Y=25886 $D=616
M302 vss 131 123 vss hvtnfet l=6e-08 w=2e-07 $X=8854 $Y=11546 $D=616
M303 vss vdd 954 vss hvtnfet l=6e-08 w=6.4e-07 $X=8879 $Y=32508 $D=616
M304 vss 124 dwlb<0> vss hvtnfet l=6e-08 w=3e-07 $X=8919 $Y=31098 $D=616
M305 vss 124 25 vss hvtnfet l=6e-08 w=3e-07 $X=8919 $Y=37457 $D=616
M306 122 ab<9> vss vss hvtnfet l=6e-08 w=2.74e-07 $X=8976 $Y=13476 $D=616
M307 111 132 955 vss hvtnfet l=6e-08 w=5.49e-07 $X=9021 $Y=17417 $D=616
M308 112 133 956 vss hvtnfet l=6e-08 w=5.49e-07 $X=9021 $Y=18966 $D=616
M309 113 132 957 vss hvtnfet l=6e-08 w=5.49e-07 $X=9021 $Y=24337 $D=616
M310 114 133 958 vss hvtnfet l=6e-08 w=5.49e-07 $X=9021 $Y=25886 $D=616
M311 b_pxbb_n<2> 135 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=9170 $Y=336 $D=616
M312 135 136 vss vss hvtnfet l=6e-08 w=5e-07 $X=9170 $Y=6701 $D=616
M313 136 137 vss vss hvtnfet l=6e-08 w=3e-07 $X=9170 $Y=7831 $D=616
M314 138 137 vss vss hvtnfet l=6e-08 w=3e-07 $X=9170 $Y=43002 $D=616
M315 139 138 vss vss hvtnfet l=6e-08 w=5e-07 $X=9170 $Y=43932 $D=616
M316 t_pxbb_n<2> 139 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=9170 $Y=49512 $D=616
M317 dwlb<0> 142 vss vss hvtnfet l=6e-08 w=3e-07 $X=9429 $Y=31098 $D=616
M318 25 143 vss vss hvtnfet l=6e-08 w=3e-07 $X=9429 $Y=37457 $D=616
M319 vss 135 b_pxbb_n<2> vss hvtnfet l=6e-08 w=1.285e-06 $X=9430 $Y=336 $D=616
M320 vss 136 135 vss hvtnfet l=6e-08 w=5e-07 $X=9430 $Y=6701 $D=616
M321 vss 137 136 vss hvtnfet l=6e-08 w=3e-07 $X=9430 $Y=7831 $D=616
M322 vss 137 138 vss hvtnfet l=6e-08 w=3e-07 $X=9430 $Y=43002 $D=616
M323 vss 138 139 vss hvtnfet l=6e-08 w=5e-07 $X=9430 $Y=43932 $D=616
M324 vss 139 t_pxbb_n<2> vss hvtnfet l=6e-08 w=1.285e-06 $X=9430 $Y=49512 $D=616
M325 vss 140 1 vss hvtnfet l=6e-08 w=2e-07 $X=9586 $Y=11276 $D=616
M326 vss 141 7 vss hvtnfet l=6e-08 w=2e-07 $X=9586 $Y=39657 $D=616
M327 vss 142 dwlb<0> vss hvtnfet l=6e-08 w=3e-07 $X=9689 $Y=31098 $D=616
M328 vss 143 25 vss hvtnfet l=6e-08 w=3e-07 $X=9689 $Y=37457 $D=616
M329 b_pxbb_n<3> 146 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=9940 $Y=336 $D=616
M330 146 147 vss vss hvtnfet l=6e-08 w=5e-07 $X=9940 $Y=6701 $D=616
M331 147 148 vss vss hvtnfet l=6e-08 w=3e-07 $X=9940 $Y=7831 $D=616
M332 149 148 vss vss hvtnfet l=6e-08 w=3e-07 $X=9940 $Y=43002 $D=616
M333 150 149 vss vss hvtnfet l=6e-08 w=5e-07 $X=9940 $Y=43932 $D=616
M334 t_pxbb_n<3> 150 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=9940 $Y=49512 $D=616
M335 vss ab<8> 129 vss hvtnfet l=6e-08 w=2.74e-07 $X=9986 $Y=13476 $D=616
M336 959 145 vss vss hvtnfet l=6e-08 w=4.11e-07 $X=10096 $Y=11276 $D=616
M337 960 145 vss vss hvtnfet l=6e-08 w=4.11e-07 $X=10096 $Y=39446 $D=616
M338 dwlb<1> 142 vss vss hvtnfet l=6e-08 w=3e-07 $X=10199 $Y=31098 $D=616
M339 24 143 vss vss hvtnfet l=6e-08 w=3e-07 $X=10199 $Y=37457 $D=616
M340 vss 146 b_pxbb_n<3> vss hvtnfet l=6e-08 w=1.285e-06 $X=10200 $Y=336 $D=616
M341 vss 147 146 vss hvtnfet l=6e-08 w=5e-07 $X=10200 $Y=6701 $D=616
M342 vss 148 147 vss hvtnfet l=6e-08 w=3e-07 $X=10200 $Y=7831 $D=616
M343 vss 148 149 vss hvtnfet l=6e-08 w=3e-07 $X=10200 $Y=43002 $D=616
M344 vss 149 150 vss hvtnfet l=6e-08 w=5e-07 $X=10200 $Y=43932 $D=616
M345 vss 150 t_pxbb_n<3> vss hvtnfet l=6e-08 w=1.285e-06 $X=10200 $Y=49512 $D=616
M346 160 129 vss vss hvtnfet l=6e-08 w=2.74e-07 $X=10246 $Y=13476 $D=616
M347 140 dwlb<1> 959 vss hvtnfet l=6e-08 w=4.11e-07 $X=10356 $Y=11276 $D=616
M348 141 dwlb<0> 960 vss hvtnfet l=6e-08 w=4.11e-07 $X=10356 $Y=39446 $D=616
M349 vss 153 124 vss hvtnfet l=6e-08 w=4e-07 $X=10406 $Y=32543 $D=616
M350 vss 142 dwlb<1> vss hvtnfet l=6e-08 w=3e-07 $X=10459 $Y=31098 $D=616
M351 vss 143 24 vss hvtnfet l=6e-08 w=3e-07 $X=10459 $Y=37457 $D=616
M352 b_pxbb_n<4> 156 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=10710 $Y=336 $D=616
M353 156 157 vss vss hvtnfet l=6e-08 w=5e-07 $X=10710 $Y=6701 $D=616
M354 157 105 vss vss hvtnfet l=6e-08 w=3e-07 $X=10710 $Y=7831 $D=616
M355 158 105 vss vss hvtnfet l=6e-08 w=3e-07 $X=10710 $Y=43002 $D=616
M356 159 158 vss vss hvtnfet l=6e-08 w=5e-07 $X=10710 $Y=43932 $D=616
M357 t_pxbb_n<4> 159 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=10710 $Y=49512 $D=616
M358 vss 132 133 vss hvtnfet l=6e-08 w=2.74e-07 $X=10846 $Y=13476 $D=616
M359 961 132 168 vss hvtnfet l=6e-08 w=5.49e-07 $X=10861 $Y=17417 $D=616
M360 962 133 169 vss hvtnfet l=6e-08 w=5.49e-07 $X=10861 $Y=18966 $D=616
M361 963 132 170 vss hvtnfet l=6e-08 w=5.49e-07 $X=10861 $Y=24337 $D=616
M362 964 133 171 vss hvtnfet l=6e-08 w=5.49e-07 $X=10861 $Y=25886 $D=616
M363 965 dwlb<1> 162 vss hvtnfet l=6e-08 w=4.11e-07 $X=10866 $Y=11276 $D=616
M364 966 dwlb<0> 163 vss hvtnfet l=6e-08 w=4.11e-07 $X=10866 $Y=39446 $D=616
M365 dwlb<1> 153 vss vss hvtnfet l=6e-08 w=3e-07 $X=10969 $Y=31098 $D=616
M366 24 153 vss vss hvtnfet l=6e-08 w=3e-07 $X=10969 $Y=37457 $D=616
M367 vss 156 b_pxbb_n<4> vss hvtnfet l=6e-08 w=1.285e-06 $X=10970 $Y=336 $D=616
M368 vss 157 156 vss hvtnfet l=6e-08 w=5e-07 $X=10970 $Y=6701 $D=616
M369 vss 105 157 vss hvtnfet l=6e-08 w=3e-07 $X=10970 $Y=7831 $D=616
M370 vss 105 158 vss hvtnfet l=6e-08 w=3e-07 $X=10970 $Y=43002 $D=616
M371 vss 158 159 vss hvtnfet l=6e-08 w=5e-07 $X=10970 $Y=43932 $D=616
M372 vss 159 t_pxbb_n<4> vss hvtnfet l=6e-08 w=1.285e-06 $X=10970 $Y=49512 $D=616
M373 132 ab<7> vss vss hvtnfet l=6e-08 w=2.74e-07 $X=11106 $Y=13476 $D=616
M374 153 154 vss vss hvtnfet l=6e-08 w=5e-07 $X=11106 $Y=32443 $D=616
M375 967 160 961 vss hvtnfet l=6e-08 w=5.49e-07 $X=11121 $Y=17417 $D=616
M376 968 160 962 vss hvtnfet l=6e-08 w=5.49e-07 $X=11121 $Y=18966 $D=616
M377 969 160 963 vss hvtnfet l=6e-08 w=5.49e-07 $X=11121 $Y=24337 $D=616
M378 970 160 964 vss hvtnfet l=6e-08 w=5.49e-07 $X=11121 $Y=25886 $D=616
M379 vss 155 965 vss hvtnfet l=6e-08 w=4.11e-07 $X=11126 $Y=11276 $D=616
M380 vss 155 966 vss hvtnfet l=6e-08 w=4.11e-07 $X=11126 $Y=39446 $D=616
M381 vss 153 dwlb<1> vss hvtnfet l=6e-08 w=3e-07 $X=11229 $Y=31098 $D=616
M382 vss 153 24 vss hvtnfet l=6e-08 w=3e-07 $X=11229 $Y=37457 $D=616
M383 971 121 967 vss hvtnfet l=6e-08 w=5.49e-07 $X=11381 $Y=17417 $D=616
M384 972 121 968 vss hvtnfet l=6e-08 w=5.49e-07 $X=11381 $Y=18966 $D=616
M385 973 122 969 vss hvtnfet l=6e-08 w=5.49e-07 $X=11381 $Y=24337 $D=616
M386 974 122 970 vss hvtnfet l=6e-08 w=5.49e-07 $X=11381 $Y=25886 $D=616
M387 b_pxbb_n<5> 164 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=11480 $Y=336 $D=616
M388 164 165 vss vss hvtnfet l=6e-08 w=5e-07 $X=11480 $Y=6701 $D=616
M389 165 106 vss vss hvtnfet l=6e-08 w=3e-07 $X=11480 $Y=7831 $D=616
M390 166 106 vss vss hvtnfet l=6e-08 w=3e-07 $X=11480 $Y=43002 $D=616
M391 167 166 vss vss hvtnfet l=6e-08 w=5e-07 $X=11480 $Y=43932 $D=616
M392 t_pxbb_n<5> 167 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=11480 $Y=49512 $D=616
M393 47 162 vss vss hvtnfet l=6e-08 w=2e-07 $X=11636 $Y=11276 $D=616
M394 50 163 vss vss hvtnfet l=6e-08 w=2e-07 $X=11636 $Y=39657 $D=616
M395 vss 43 971 vss hvtnfet l=6e-08 w=8.23e-07 $X=11651 $Y=17143 $D=616
M396 vss 43 972 vss hvtnfet l=6e-08 w=8.23e-07 $X=11651 $Y=18966 $D=616
M397 vss 43 973 vss hvtnfet l=6e-08 w=8.23e-07 $X=11651 $Y=24063 $D=616
M398 vss 43 974 vss hvtnfet l=6e-08 w=8.23e-07 $X=11651 $Y=25886 $D=616
M399 172 142 vss vss hvtnfet l=6e-08 w=2e-07 $X=11739 $Y=31098 $D=616
M400 vss 164 b_pxbb_n<5> vss hvtnfet l=6e-08 w=1.285e-06 $X=11740 $Y=336 $D=616
M401 vss 165 164 vss hvtnfet l=6e-08 w=5e-07 $X=11740 $Y=6701 $D=616
M402 vss 106 165 vss hvtnfet l=6e-08 w=3e-07 $X=11740 $Y=7831 $D=616
M403 vss 106 166 vss hvtnfet l=6e-08 w=3e-07 $X=11740 $Y=43002 $D=616
M404 vss 166 167 vss hvtnfet l=6e-08 w=5e-07 $X=11740 $Y=43932 $D=616
M405 vss 167 t_pxbb_n<5> vss hvtnfet l=6e-08 w=1.285e-06 $X=11740 $Y=49512 $D=616
M406 vss tm<0> dbl_pd_n<0> vss hvtnfet l=6e-08 w=2.14e-07 $X=11746 $Y=13361 $D=616
M407 dbl_pd_n<0> tm<0> vss vss hvtnfet l=6e-08 w=2.14e-07 $X=12006 $Y=13361 $D=616
M408 179 173 vss vss hvtnfet l=6e-08 w=2e-07 $X=12086 $Y=32533 $D=616
M409 vss 174 2 vss hvtnfet l=6e-08 w=2e-07 $X=12146 $Y=11276 $D=616
M410 177 168 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=12146 $Y=17812 $D=616
M411 178 169 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=12146 $Y=18983 $D=616
M412 137 170 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=12146 $Y=24732 $D=616
M413 148 171 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=12146 $Y=25903 $D=616
M414 vss 175 6 vss hvtnfet l=6e-08 w=2e-07 $X=12146 $Y=39657 $D=616
M415 975 33 168 vss hvtnfet l=6e-08 w=1.8e-07 $X=12161 $Y=17143 $D=616
M416 976 33 169 vss hvtnfet l=6e-08 w=1.8e-07 $X=12161 $Y=19609 $D=616
M417 977 33 170 vss hvtnfet l=6e-08 w=1.8e-07 $X=12161 $Y=24063 $D=616
M418 978 33 171 vss hvtnfet l=6e-08 w=1.8e-07 $X=12161 $Y=26529 $D=616
M419 vss 172 143 vss hvtnfet l=6e-08 w=6e-07 $X=12193 $Y=37037 $D=616
M420 b_pxbb_n<6> 180 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=12250 $Y=336 $D=616
M421 180 181 vss vss hvtnfet l=6e-08 w=5e-07 $X=12250 $Y=6701 $D=616
M422 181 177 vss vss hvtnfet l=6e-08 w=3e-07 $X=12250 $Y=7831 $D=616
M423 182 177 vss vss hvtnfet l=6e-08 w=3e-07 $X=12250 $Y=43002 $D=616
M424 183 182 vss vss hvtnfet l=6e-08 w=5e-07 $X=12250 $Y=43932 $D=616
M425 t_pxbb_n<6> 183 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=12250 $Y=49512 $D=616
M426 vss tm<0> dbl_pd_n<0> vss hvtnfet l=6e-08 w=2.14e-07 $X=12266 $Y=13361 $D=616
M427 vss 142 184 vss hvtnfet l=2.5e-07 w=3.5e-07 $X=12309 $Y=30853 $D=616
M428 vss 168 177 vss hvtnfet l=6e-08 w=1.37e-07 $X=12406 $Y=17812 $D=616
M429 vss 169 178 vss hvtnfet l=6e-08 w=1.37e-07 $X=12406 $Y=18983 $D=616
M430 vss 170 137 vss hvtnfet l=6e-08 w=1.37e-07 $X=12406 $Y=24732 $D=616
M431 vss 171 148 vss hvtnfet l=6e-08 w=1.37e-07 $X=12406 $Y=25903 $D=616
M432 vss 177 975 vss hvtnfet l=6e-08 w=1.8e-07 $X=12421 $Y=17143 $D=616
M433 vss 178 976 vss hvtnfet l=6e-08 w=1.8e-07 $X=12421 $Y=19609 $D=616
M434 vss 137 977 vss hvtnfet l=6e-08 w=1.8e-07 $X=12421 $Y=24063 $D=616
M435 vss 148 978 vss hvtnfet l=6e-08 w=1.8e-07 $X=12421 $Y=26529 $D=616
M436 vss 180 b_pxbb_n<6> vss hvtnfet l=6e-08 w=1.285e-06 $X=12510 $Y=336 $D=616
M437 vss 181 180 vss hvtnfet l=6e-08 w=5e-07 $X=12510 $Y=6701 $D=616
M438 vss 177 181 vss hvtnfet l=6e-08 w=3e-07 $X=12510 $Y=7831 $D=616
M439 vss 177 182 vss hvtnfet l=6e-08 w=3e-07 $X=12510 $Y=43002 $D=616
M440 vss 182 183 vss hvtnfet l=6e-08 w=5e-07 $X=12510 $Y=43932 $D=616
M441 vss 183 t_pxbb_n<6> vss hvtnfet l=6e-08 w=1.285e-06 $X=12510 $Y=49512 $D=616
M442 vss 179 186 vss hvtnfet l=6e-08 w=2e-07 $X=12596 $Y=32533 $D=616
M443 979 185 vss vss hvtnfet l=6e-08 w=4.11e-07 $X=12656 $Y=11276 $D=616
M444 980 185 vss vss hvtnfet l=6e-08 w=4.11e-07 $X=12656 $Y=39446 $D=616
M445 191 184 vss vss hvtnfet l=6e-08 w=3.5e-07 $X=12759 $Y=30853 $D=616
M446 vss 131 dbl_pd_n<2> vss hvtnfet l=6e-08 w=2.14e-07 $X=12776 $Y=13361 $D=616
M447 186 191 vss vss hvtnfet l=6e-08 w=2e-07 $X=12856 $Y=32533 $D=616
M448 174 dwlb<1> 979 vss hvtnfet l=6e-08 w=4.11e-07 $X=12916 $Y=11276 $D=616
M449 175 dwlb<0> 980 vss hvtnfet l=6e-08 w=4.11e-07 $X=12916 $Y=39446 $D=616
M450 981 187 vss vss hvtnfet l=6e-08 w=1.8e-07 $X=12931 $Y=17143 $D=616
M451 982 188 vss vss hvtnfet l=6e-08 w=1.8e-07 $X=12931 $Y=19609 $D=616
M452 983 189 vss vss hvtnfet l=6e-08 w=1.8e-07 $X=12931 $Y=24063 $D=616
M453 984 190 vss vss hvtnfet l=6e-08 w=1.8e-07 $X=12931 $Y=26529 $D=616
M454 187 192 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=12946 $Y=17812 $D=616
M455 188 193 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=12946 $Y=18983 $D=616
M456 189 194 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=12946 $Y=24732 $D=616
M457 190 195 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=12946 $Y=25903 $D=616
M458 vss 186 143 vss hvtnfet l=6e-08 w=6e-07 $X=12973 $Y=37037 $D=616
M459 b_pxbb_n<7> 196 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=13020 $Y=336 $D=616
M460 196 197 vss vss hvtnfet l=6e-08 w=5e-07 $X=13020 $Y=6701 $D=616
M461 197 178 vss vss hvtnfet l=6e-08 w=3e-07 $X=13020 $Y=7831 $D=616
M462 198 178 vss vss hvtnfet l=6e-08 w=3e-07 $X=13020 $Y=43002 $D=616
M463 199 198 vss vss hvtnfet l=6e-08 w=5e-07 $X=13020 $Y=43932 $D=616
M464 t_pxbb_n<7> 199 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=13020 $Y=49512 $D=616
M465 dbl_pd_n<2> 131 vss vss hvtnfet l=6e-08 w=2.14e-07 $X=13036 $Y=13361 $D=616
M466 192 33 981 vss hvtnfet l=6e-08 w=1.8e-07 $X=13191 $Y=17143 $D=616
M467 193 33 982 vss hvtnfet l=6e-08 w=1.8e-07 $X=13191 $Y=19609 $D=616
M468 194 33 983 vss hvtnfet l=6e-08 w=1.8e-07 $X=13191 $Y=24063 $D=616
M469 195 33 984 vss hvtnfet l=6e-08 w=1.8e-07 $X=13191 $Y=26529 $D=616
M470 vss 192 187 vss hvtnfet l=6e-08 w=1.37e-07 $X=13206 $Y=17812 $D=616
M471 vss 193 188 vss hvtnfet l=6e-08 w=1.37e-07 $X=13206 $Y=18983 $D=616
M472 vss 194 189 vss hvtnfet l=6e-08 w=1.37e-07 $X=13206 $Y=24732 $D=616
M473 vss 195 190 vss hvtnfet l=6e-08 w=1.37e-07 $X=13206 $Y=25903 $D=616
M474 vss 196 b_pxbb_n<7> vss hvtnfet l=6e-08 w=1.285e-06 $X=13280 $Y=336 $D=616
M475 vss 197 196 vss hvtnfet l=6e-08 w=5e-07 $X=13280 $Y=6701 $D=616
M476 vss 178 197 vss hvtnfet l=6e-08 w=3e-07 $X=13280 $Y=7831 $D=616
M477 vss 178 198 vss hvtnfet l=6e-08 w=3e-07 $X=13280 $Y=43002 $D=616
M478 vss 198 199 vss hvtnfet l=6e-08 w=5e-07 $X=13280 $Y=43932 $D=616
M479 vss 199 t_pxbb_n<7> vss hvtnfet l=6e-08 w=1.285e-06 $X=13280 $Y=49512 $D=616
M480 vss 131 dbl_pd_n<2> vss hvtnfet l=6e-08 w=2.14e-07 $X=13296 $Y=13361 $D=616
M481 vss 191 202 vss hvtnfet l=2.5e-07 w=3.5e-07 $X=13429 $Y=30853 $D=616
M482 vss tm<7> 203 vss hvtnfet l=6e-08 w=2e-07 $X=13432 $Y=32533 $D=616
M483 985 43 vss vss hvtnfet l=6e-08 w=8.23e-07 $X=13701 $Y=17143 $D=616
M484 986 43 vss vss hvtnfet l=6e-08 w=8.23e-07 $X=13701 $Y=18966 $D=616
M485 987 43 vss vss hvtnfet l=6e-08 w=8.23e-07 $X=13701 $Y=24063 $D=616
M486 988 43 vss vss hvtnfet l=6e-08 w=8.23e-07 $X=13701 $Y=25886 $D=616
M487 vss 200 143 vss hvtnfet l=6e-08 w=6e-07 $X=13753 $Y=37037 $D=616
M488 b_pxcb_n<0> 206 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=13790 $Y=336 $D=616
M489 206 207 vss vss hvtnfet l=6e-08 w=5e-07 $X=13790 $Y=6701 $D=616
M490 207 189 vss vss hvtnfet l=6e-08 w=3e-07 $X=13790 $Y=7831 $D=616
M491 208 189 vss vss hvtnfet l=6e-08 w=3e-07 $X=13790 $Y=43002 $D=616
M492 209 208 vss vss hvtnfet l=6e-08 w=5e-07 $X=13790 $Y=43932 $D=616
M493 t_pxcb_n<0> 209 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=13790 $Y=49512 $D=616
M494 211 202 vss vss hvtnfet l=6e-08 w=3.5e-07 $X=13879 $Y=30853 $D=616
M495 vss 205 204 vss hvtnfet l=6e-08 w=2.74e-07 $X=13936 $Y=13476 $D=616
M496 vss 203 200 vss hvtnfet l=6e-08 w=2e-07 $X=13942 $Y=32533 $D=616
M497 989 204 985 vss hvtnfet l=6e-08 w=5.49e-07 $X=13971 $Y=17417 $D=616
M498 990 204 986 vss hvtnfet l=6e-08 w=5.49e-07 $X=13971 $Y=18966 $D=616
M499 991 205 987 vss hvtnfet l=6e-08 w=5.49e-07 $X=13971 $Y=24337 $D=616
M500 992 205 988 vss hvtnfet l=6e-08 w=5.49e-07 $X=13971 $Y=25886 $D=616
M501 vss 206 b_pxcb_n<0> vss hvtnfet l=6e-08 w=1.285e-06 $X=14050 $Y=336 $D=616
M502 vss 207 206 vss hvtnfet l=6e-08 w=5e-07 $X=14050 $Y=6701 $D=616
M503 vss 189 207 vss hvtnfet l=6e-08 w=3e-07 $X=14050 $Y=7831 $D=616
M504 vss 189 208 vss hvtnfet l=6e-08 w=3e-07 $X=14050 $Y=43002 $D=616
M505 vss 208 209 vss hvtnfet l=6e-08 w=5e-07 $X=14050 $Y=43932 $D=616
M506 vss 209 t_pxcb_n<0> vss hvtnfet l=6e-08 w=1.285e-06 $X=14050 $Y=49512 $D=616
M507 200 211 vss vss hvtnfet l=6e-08 w=2e-07 $X=14202 $Y=32533 $D=616
M508 993 dwlb<1> 216 vss hvtnfet l=6e-08 w=4.11e-07 $X=14216 $Y=11276 $D=616
M509 994 dwlb<0> 217 vss hvtnfet l=6e-08 w=4.11e-07 $X=14216 $Y=39446 $D=616
M510 995 210 989 vss hvtnfet l=6e-08 w=5.49e-07 $X=14231 $Y=17417 $D=616
M511 996 210 990 vss hvtnfet l=6e-08 w=5.49e-07 $X=14231 $Y=18966 $D=616
M512 997 210 991 vss hvtnfet l=6e-08 w=5.49e-07 $X=14231 $Y=24337 $D=616
M513 998 210 992 vss hvtnfet l=6e-08 w=5.49e-07 $X=14231 $Y=25886 $D=616
M514 205 ab<12> vss vss hvtnfet l=6e-08 w=2.74e-07 $X=14446 $Y=13476 $D=616
M515 vss 212 993 vss hvtnfet l=6e-08 w=4.11e-07 $X=14476 $Y=11276 $D=616
M516 vss 212 994 vss hvtnfet l=6e-08 w=4.11e-07 $X=14476 $Y=39446 $D=616
M517 192 213 995 vss hvtnfet l=6e-08 w=5.49e-07 $X=14491 $Y=17417 $D=616
M518 193 214 996 vss hvtnfet l=6e-08 w=5.49e-07 $X=14491 $Y=18966 $D=616
M519 194 213 997 vss hvtnfet l=6e-08 w=5.49e-07 $X=14491 $Y=24337 $D=616
M520 195 214 998 vss hvtnfet l=6e-08 w=5.49e-07 $X=14491 $Y=25886 $D=616
M521 b_pxcb_n<1> 218 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=14560 $Y=336 $D=616
M522 218 219 vss vss hvtnfet l=6e-08 w=5e-07 $X=14560 $Y=6701 $D=616
M523 219 190 vss vss hvtnfet l=6e-08 w=3e-07 $X=14560 $Y=7831 $D=616
M524 220 190 vss vss hvtnfet l=6e-08 w=3e-07 $X=14560 $Y=43002 $D=616
M525 221 220 vss vss hvtnfet l=6e-08 w=5e-07 $X=14560 $Y=43932 $D=616
M526 t_pxcb_n<1> 221 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=14560 $Y=49512 $D=616
M527 vss 123 624 vss hvtnfet l=6e-08 w=6e-07 $X=14796 $Y=30668 $D=616
M528 vss 218 b_pxcb_n<1> vss hvtnfet l=6e-08 w=1.285e-06 $X=14820 $Y=336 $D=616
M529 vss 219 218 vss hvtnfet l=6e-08 w=5e-07 $X=14820 $Y=6701 $D=616
M530 vss 190 219 vss hvtnfet l=6e-08 w=3e-07 $X=14820 $Y=7831 $D=616
M531 vss 190 220 vss hvtnfet l=6e-08 w=3e-07 $X=14820 $Y=43002 $D=616
M532 vss 220 221 vss hvtnfet l=6e-08 w=5e-07 $X=14820 $Y=43932 $D=616
M533 vss 221 t_pxcb_n<1> vss hvtnfet l=6e-08 w=1.285e-06 $X=14820 $Y=49512 $D=616
M534 vss 72 58 vss hvtnfet l=6e-08 w=2e-07 $X=14872 $Y=37045 $D=616
M535 48 216 vss vss hvtnfet l=6e-08 w=2e-07 $X=14986 $Y=11276 $D=616
M536 49 217 vss vss hvtnfet l=6e-08 w=2e-07 $X=14986 $Y=39657 $D=616
M537 vss 43 33 vss hvtnfet l=6e-08 w=7e-07 $X=15316 $Y=30668 $D=616
M538 b_pxcb_n<2> 223 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=15330 $Y=336 $D=616
M539 223 224 vss vss hvtnfet l=6e-08 w=5e-07 $X=15330 $Y=6701 $D=616
M540 224 225 vss vss hvtnfet l=6e-08 w=3e-07 $X=15330 $Y=7831 $D=616
M541 226 225 vss vss hvtnfet l=6e-08 w=3e-07 $X=15330 $Y=43002 $D=616
M542 227 226 vss vss hvtnfet l=6e-08 w=5e-07 $X=15330 $Y=43932 $D=616
M543 t_pxcb_n<2> 227 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=15330 $Y=49512 $D=616
M544 629 229 vss vss hvtnfet l=6e-08 w=4e-07 $X=15382 $Y=37045 $D=616
M545 vss ab<11> 210 vss hvtnfet l=6e-08 w=2.74e-07 $X=15456 $Y=13476 $D=616
M546 33 43 vss vss hvtnfet l=6e-08 w=7e-07 $X=15576 $Y=30668 $D=616
M547 vss 223 b_pxcb_n<2> vss hvtnfet l=6e-08 w=1.285e-06 $X=15590 $Y=336 $D=616
M548 vss 224 223 vss hvtnfet l=6e-08 w=5e-07 $X=15590 $Y=6701 $D=616
M549 vss 225 224 vss hvtnfet l=6e-08 w=3e-07 $X=15590 $Y=7831 $D=616
M550 vss 225 226 vss hvtnfet l=6e-08 w=3e-07 $X=15590 $Y=43002 $D=616
M551 vss 226 227 vss hvtnfet l=6e-08 w=5e-07 $X=15590 $Y=43932 $D=616
M552 vss 227 t_pxcb_n<2> vss hvtnfet l=6e-08 w=1.285e-06 $X=15590 $Y=49512 $D=616
M553 vss 228 231 vss hvtnfet l=6e-08 w=2.1e-07 $X=15621 $Y=32688 $D=616
M554 72 172 629 vss hvtnfet l=6e-08 w=4e-07 $X=15642 $Y=37045 $D=616
M555 240 210 vss vss hvtnfet l=6e-08 w=2.74e-07 $X=15716 $Y=13476 $D=616
M556 631 tm<0> vss vss hvtnfet l=6e-08 w=2.74e-07 $X=15880 $Y=39358 $D=616
M557 630 131 vss vss hvtnfet l=6e-08 w=2.1e-07 $X=15881 $Y=32688 $D=616
M558 vss tm<3> 242 vss hvtnfet l=7e-08 w=3.2e-07 $X=16057 $Y=11276 $D=616
M559 b_pxcb_n<3> 235 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=16100 $Y=336 $D=616
M560 235 236 vss vss hvtnfet l=6e-08 w=5e-07 $X=16100 $Y=6701 $D=616
M561 236 237 vss vss hvtnfet l=6e-08 w=3e-07 $X=16100 $Y=7831 $D=616
M562 238 237 vss vss hvtnfet l=6e-08 w=3e-07 $X=16100 $Y=43002 $D=616
M563 239 238 vss vss hvtnfet l=6e-08 w=5e-07 $X=16100 $Y=43932 $D=616
M564 t_pxcb_n<3> 239 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=16100 $Y=49512 $D=616
M565 228 231 630 vss hvtnfet l=6e-08 w=2.1e-07 $X=16141 $Y=32688 $D=616
M566 vss 213 214 vss hvtnfet l=6e-08 w=2.74e-07 $X=16316 $Y=13476 $D=616
M567 635 232 vss vss hvtnfet l=6e-08 w=3.2e-07 $X=16322 $Y=37277 $D=616
M568 243 tm<4> vss vss hvtnfet l=7e-08 w=3.2e-07 $X=16327 $Y=11276 $D=616
M569 999 213 249 vss hvtnfet l=6e-08 w=5.49e-07 $X=16331 $Y=17417 $D=616
M570 1000 214 250 vss hvtnfet l=6e-08 w=5.49e-07 $X=16331 $Y=18966 $D=616
M571 1001 213 251 vss hvtnfet l=6e-08 w=5.49e-07 $X=16331 $Y=24337 $D=616
M572 1002 214 252 vss hvtnfet l=6e-08 w=5.49e-07 $X=16331 $Y=25886 $D=616
M573 vss 123 644 vss hvtnfet l=6e-08 w=6e-07 $X=16346 $Y=30668 $D=616
M574 vss 235 b_pxcb_n<3> vss hvtnfet l=6e-08 w=1.285e-06 $X=16360 $Y=336 $D=616
M575 vss 236 235 vss hvtnfet l=6e-08 w=5e-07 $X=16360 $Y=6701 $D=616
M576 vss 237 236 vss hvtnfet l=6e-08 w=3e-07 $X=16360 $Y=7831 $D=616
M577 vss 237 238 vss hvtnfet l=6e-08 w=3e-07 $X=16360 $Y=43002 $D=616
M578 vss 238 239 vss hvtnfet l=6e-08 w=5e-07 $X=16360 $Y=43932 $D=616
M579 vss 239 t_pxcb_n<3> vss hvtnfet l=6e-08 w=1.285e-06 $X=16360 $Y=49512 $D=616
M580 636 123 228 vss hvtnfet l=6e-08 w=3.2e-07 $X=16401 $Y=32578 $D=616
M581 213 ab<10> vss vss hvtnfet l=6e-08 w=2.74e-07 $X=16576 $Y=13476 $D=616
M582 229 142 635 vss hvtnfet l=6e-08 w=3.2e-07 $X=16582 $Y=37277 $D=616
M583 1003 240 999 vss hvtnfet l=6e-08 w=5.49e-07 $X=16591 $Y=17417 $D=616
M584 1004 240 1000 vss hvtnfet l=6e-08 w=5.49e-07 $X=16591 $Y=18966 $D=616
M585 1005 240 1001 vss hvtnfet l=6e-08 w=5.49e-07 $X=16591 $Y=24337 $D=616
M586 1006 240 1002 vss hvtnfet l=6e-08 w=5.49e-07 $X=16591 $Y=25886 $D=616
M587 644 123 vss vss hvtnfet l=6e-08 w=6e-07 $X=16606 $Y=30668 $D=616
M588 vss 123 636 vss hvtnfet l=6e-08 w=3.2e-07 $X=16661 $Y=32578 $D=616
M589 637 tm<6> vss vss hvtnfet l=6e-08 w=2.74e-07 $X=16680 $Y=39358 $D=616
M590 638 244 229 vss hvtnfet l=6e-08 w=2.1e-07 $X=16842 $Y=37277 $D=616
M591 vss 243 643 vss hvtnfet l=6e-08 w=4.8e-07 $X=16847 $Y=11276 $D=616
M592 1007 204 1003 vss hvtnfet l=6e-08 w=5.49e-07 $X=16851 $Y=17417 $D=616
M593 1008 204 1004 vss hvtnfet l=6e-08 w=5.49e-07 $X=16851 $Y=18966 $D=616
M594 1009 205 1005 vss hvtnfet l=6e-08 w=5.49e-07 $X=16851 $Y=24337 $D=616
M595 1010 205 1006 vss hvtnfet l=6e-08 w=5.49e-07 $X=16851 $Y=25886 $D=616
M596 642 123 644 vss hvtnfet l=6e-08 w=6e-07 $X=16866 $Y=30668 $D=616
M597 b_pxcb_n<4> 245 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=16870 $Y=336 $D=616
M598 245 246 vss vss hvtnfet l=6e-08 w=5e-07 $X=16870 $Y=6701 $D=616
M599 246 187 vss vss hvtnfet l=6e-08 w=3e-07 $X=16870 $Y=7831 $D=616
M600 247 187 vss vss hvtnfet l=6e-08 w=3e-07 $X=16870 $Y=43002 $D=616
M601 248 247 vss vss hvtnfet l=6e-08 w=5e-07 $X=16870 $Y=43932 $D=616
M602 t_pxcb_n<4> 248 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=16870 $Y=49512 $D=616
M603 vss 172 638 vss hvtnfet l=6e-08 w=2.1e-07 $X=17102 $Y=37277 $D=616
M604 643 242 vss vss hvtnfet l=6e-08 w=4.8e-07 $X=17107 $Y=11276 $D=616
M605 vss 43 1007 vss hvtnfet l=6e-08 w=8.23e-07 $X=17121 $Y=17143 $D=616
M606 vss 43 1008 vss hvtnfet l=6e-08 w=8.23e-07 $X=17121 $Y=18966 $D=616
M607 vss 43 1009 vss hvtnfet l=6e-08 w=8.23e-07 $X=17121 $Y=24063 $D=616
M608 vss 43 1010 vss hvtnfet l=6e-08 w=8.23e-07 $X=17121 $Y=25886 $D=616
M609 644 123 642 vss hvtnfet l=6e-08 w=6e-07 $X=17126 $Y=30668 $D=616
M610 vss 245 b_pxcb_n<4> vss hvtnfet l=6e-08 w=1.285e-06 $X=17130 $Y=336 $D=616
M611 vss 246 245 vss hvtnfet l=6e-08 w=5e-07 $X=17130 $Y=6701 $D=616
M612 vss 187 246 vss hvtnfet l=6e-08 w=3e-07 $X=17130 $Y=7831 $D=616
M613 vss 187 247 vss hvtnfet l=6e-08 w=3e-07 $X=17130 $Y=43002 $D=616
M614 vss 247 248 vss hvtnfet l=6e-08 w=5e-07 $X=17130 $Y=43932 $D=616
M615 vss 248 t_pxcb_n<4> vss hvtnfet l=6e-08 w=1.285e-06 $X=17130 $Y=49512 $D=616
M616 244 229 vss vss hvtnfet l=6e-08 w=2.1e-07 $X=17362 $Y=37277 $D=616
M617 253 249 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=17616 $Y=17812 $D=616
M618 254 250 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=17616 $Y=18983 $D=616
M619 225 251 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=17616 $Y=24732 $D=616
M620 237 252 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=17616 $Y=25903 $D=616
M621 647 242 vss vss hvtnfet l=6e-08 w=4.8e-07 $X=17617 $Y=11276 $D=616
M622 1011 33 249 vss hvtnfet l=6e-08 w=1.8e-07 $X=17631 $Y=17143 $D=616
M623 1012 33 250 vss hvtnfet l=6e-08 w=1.8e-07 $X=17631 $Y=19609 $D=616
M624 1013 33 251 vss hvtnfet l=6e-08 w=1.8e-07 $X=17631 $Y=24063 $D=616
M625 1014 33 252 vss hvtnfet l=6e-08 w=1.8e-07 $X=17631 $Y=26529 $D=616
M626 b_pxcb_n<5> 255 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=17640 $Y=336 $D=616
M627 255 256 vss vss hvtnfet l=6e-08 w=5e-07 $X=17640 $Y=6701 $D=616
M628 256 188 vss vss hvtnfet l=6e-08 w=3e-07 $X=17640 $Y=7831 $D=616
M629 257 188 vss vss hvtnfet l=6e-08 w=3e-07 $X=17640 $Y=43002 $D=616
M630 258 257 vss vss hvtnfet l=6e-08 w=5e-07 $X=17640 $Y=43932 $D=616
M631 t_pxcb_n<5> 258 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=17640 $Y=49512 $D=616
M632 23 clkb vss vss hvtnfet l=6e-08 w=4.5e-07 $X=17646 $Y=30668 $D=616
M633 vss 249 253 vss hvtnfet l=6e-08 w=1.37e-07 $X=17876 $Y=17812 $D=616
M634 vss 250 254 vss hvtnfet l=6e-08 w=1.37e-07 $X=17876 $Y=18983 $D=616
M635 vss 251 225 vss hvtnfet l=6e-08 w=1.37e-07 $X=17876 $Y=24732 $D=616
M636 vss 252 237 vss hvtnfet l=6e-08 w=1.37e-07 $X=17876 $Y=25903 $D=616
M637 vss tm<4> 647 vss hvtnfet l=6e-08 w=4.8e-07 $X=17877 $Y=11276 $D=616
M638 vss 253 1011 vss hvtnfet l=6e-08 w=1.8e-07 $X=17891 $Y=17143 $D=616
M639 vss 254 1012 vss hvtnfet l=6e-08 w=1.8e-07 $X=17891 $Y=19609 $D=616
M640 vss 225 1013 vss hvtnfet l=6e-08 w=1.8e-07 $X=17891 $Y=24063 $D=616
M641 vss 237 1014 vss hvtnfet l=6e-08 w=1.8e-07 $X=17891 $Y=26529 $D=616
M642 vss 255 b_pxcb_n<5> vss hvtnfet l=6e-08 w=1.285e-06 $X=17900 $Y=336 $D=616
M643 vss 256 255 vss hvtnfet l=6e-08 w=5e-07 $X=17900 $Y=6701 $D=616
M644 vss 188 256 vss hvtnfet l=6e-08 w=3e-07 $X=17900 $Y=7831 $D=616
M645 vss 188 257 vss hvtnfet l=6e-08 w=3e-07 $X=17900 $Y=43002 $D=616
M646 vss 257 258 vss hvtnfet l=6e-08 w=5e-07 $X=17900 $Y=43932 $D=616
M647 vss 258 t_pxcb_n<5> vss hvtnfet l=6e-08 w=1.285e-06 $X=17900 $Y=49512 $D=616
M648 vss 260 273 vss hvtnfet l=6e-08 w=2.74e-07 $X=18106 $Y=13476 $D=616
M649 vss wenb 232 vss hvtnfet l=6e-08 w=2e-07 $X=18366 $Y=37147 $D=616
M650 648 tm<4> vss vss hvtnfet l=6e-08 w=4.8e-07 $X=18387 $Y=11276 $D=616
M651 b_pxcb_n<6> 265 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=18410 $Y=336 $D=616
M652 265 266 vss vss hvtnfet l=6e-08 w=5e-07 $X=18410 $Y=6701 $D=616
M653 266 253 vss vss hvtnfet l=6e-08 w=3e-07 $X=18410 $Y=7831 $D=616
M654 267 253 vss vss hvtnfet l=6e-08 w=3e-07 $X=18410 $Y=43002 $D=616
M655 268 267 vss vss hvtnfet l=6e-08 w=5e-07 $X=18410 $Y=43932 $D=616
M656 t_pxcb_n<6> 268 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=18410 $Y=49512 $D=616
M657 651 ab<4> vss vss hvtnfet l=6e-08 w=3.2e-07 $X=18460 $Y=30918 $D=616
M658 652 wenb vss vss hvtnfet l=6e-08 w=3.2e-07 $X=18460 $Y=32578 $D=616
M659 vss tm<2> 173 vss hvtnfet l=6e-08 w=2.74e-07 $X=18510 $Y=39358 $D=616
M660 260 ab<1> vss vss hvtnfet l=6e-08 w=2.74e-07 $X=18616 $Y=13476 $D=616
M661 232 264 vss vss hvtnfet l=6e-08 w=2e-07 $X=18626 $Y=37147 $D=616
M662 vss tm<3> 648 vss hvtnfet l=6e-08 w=4.8e-07 $X=18647 $Y=11276 $D=616
M663 vss 265 b_pxcb_n<6> vss hvtnfet l=6e-08 w=1.285e-06 $X=18670 $Y=336 $D=616
M664 vss 266 265 vss hvtnfet l=6e-08 w=5e-07 $X=18670 $Y=6701 $D=616
M665 vss 253 266 vss hvtnfet l=6e-08 w=3e-07 $X=18670 $Y=7831 $D=616
M666 vss 253 267 vss hvtnfet l=6e-08 w=3e-07 $X=18670 $Y=43002 $D=616
M667 vss 267 268 vss hvtnfet l=6e-08 w=5e-07 $X=18670 $Y=43932 $D=616
M668 vss 268 t_pxcb_n<6> vss hvtnfet l=6e-08 w=1.285e-06 $X=18670 $Y=49512 $D=616
M669 154 23 651 vss hvtnfet l=6e-08 w=3.2e-07 $X=18720 $Y=30918 $D=616
M670 274 23 652 vss hvtnfet l=6e-08 w=3.2e-07 $X=18720 $Y=32578 $D=616
M671 1015 269 280 vss hvtnfet l=6e-08 w=5.49e-07 $X=18911 $Y=17143 $D=616
M672 1016 270 281 vss hvtnfet l=6e-08 w=5.49e-07 $X=18911 $Y=19240 $D=616
M673 1017 269 282 vss hvtnfet l=6e-08 w=5.49e-07 $X=18911 $Y=24063 $D=616
M674 1018 270 283 vss hvtnfet l=6e-08 w=5.49e-07 $X=18911 $Y=26160 $D=616
M675 653 271 154 vss hvtnfet l=6e-08 w=2.1e-07 $X=18980 $Y=30918 $D=616
M676 654 272 274 vss hvtnfet l=6e-08 w=2.1e-07 $X=18980 $Y=32688 $D=616
M677 vss 270 269 vss hvtnfet l=6e-08 w=2.74e-07 $X=19126 $Y=13476 $D=616
M678 659 tm<3> vss vss hvtnfet l=6e-08 w=4.8e-07 $X=19157 $Y=11276 $D=616
M679 1019 273 1015 vss hvtnfet l=6e-08 w=5.49e-07 $X=19171 $Y=17143 $D=616
M680 1020 273 1016 vss hvtnfet l=6e-08 w=5.49e-07 $X=19171 $Y=19240 $D=616
M681 1021 260 1017 vss hvtnfet l=6e-08 w=5.49e-07 $X=19171 $Y=24063 $D=616
M682 1022 260 1018 vss hvtnfet l=6e-08 w=5.49e-07 $X=19171 $Y=26160 $D=616
M683 b_pxcb_n<7> 275 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=19180 $Y=336 $D=616
M684 275 276 vss vss hvtnfet l=6e-08 w=5e-07 $X=19180 $Y=6701 $D=616
M685 276 254 vss vss hvtnfet l=6e-08 w=3e-07 $X=19180 $Y=7831 $D=616
M686 277 254 vss vss hvtnfet l=6e-08 w=3e-07 $X=19180 $Y=43002 $D=616
M687 278 277 vss vss hvtnfet l=6e-08 w=5e-07 $X=19180 $Y=43932 $D=616
M688 t_pxcb_n<7> 278 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=19180 $Y=49512 $D=616
M689 vss clkb 653 vss hvtnfet l=6e-08 w=2.1e-07 $X=19240 $Y=30918 $D=616
M690 vss clkb 654 vss hvtnfet l=6e-08 w=2.1e-07 $X=19240 $Y=32688 $D=616
M691 vss 243 659 vss hvtnfet l=6e-08 w=4.8e-07 $X=19417 $Y=11276 $D=616
M692 vss 275 b_pxcb_n<7> vss hvtnfet l=6e-08 w=1.285e-06 $X=19440 $Y=336 $D=616
M693 vss 276 275 vss hvtnfet l=6e-08 w=5e-07 $X=19440 $Y=6701 $D=616
M694 vss 254 276 vss hvtnfet l=6e-08 w=3e-07 $X=19440 $Y=7831 $D=616
M695 vss 254 277 vss hvtnfet l=6e-08 w=3e-07 $X=19440 $Y=43002 $D=616
M696 vss 277 278 vss hvtnfet l=6e-08 w=5e-07 $X=19440 $Y=43932 $D=616
M697 vss 278 t_pxcb_n<7> vss hvtnfet l=6e-08 w=1.285e-06 $X=19440 $Y=49512 $D=616
M698 vss 43 1019 vss hvtnfet l=6e-08 w=8.23e-07 $X=19441 $Y=17143 $D=616
M699 vss 43 1020 vss hvtnfet l=6e-08 w=8.23e-07 $X=19441 $Y=18966 $D=616
M700 vss 43 1021 vss hvtnfet l=6e-08 w=8.23e-07 $X=19441 $Y=24063 $D=616
M701 vss 43 1022 vss hvtnfet l=6e-08 w=8.23e-07 $X=19441 $Y=25886 $D=616
M702 271 154 vss vss hvtnfet l=6e-08 w=2.1e-07 $X=19500 $Y=30918 $D=616
M703 272 274 vss vss hvtnfet l=6e-08 w=2.1e-07 $X=19500 $Y=32688 $D=616
M704 270 ab<0> vss vss hvtnfet l=6e-08 w=2.74e-07 $X=19636 $Y=13476 $D=616
M705 vss 15 r_saeb_n vss hvtnfet l=6e-08 w=8.58e-07 $X=19675 $Y=37027 $D=616
M706 r_saeb_n 15 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=19935 $Y=37027 $D=616
M707 1023 33 280 vss hvtnfet l=6e-08 w=1.8e-07 $X=19951 $Y=17143 $D=616
M708 212 280 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=19951 $Y=17812 $D=616
M709 185 281 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=19951 $Y=18983 $D=616
M710 1024 33 281 vss hvtnfet l=6e-08 w=1.8e-07 $X=19951 $Y=19609 $D=616
M711 1025 33 282 vss hvtnfet l=6e-08 w=1.8e-07 $X=19951 $Y=24063 $D=616
M712 155 282 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=19951 $Y=24732 $D=616
M713 145 283 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=19951 $Y=25903 $D=616
M714 1026 33 283 vss hvtnfet l=6e-08 w=1.8e-07 $X=19951 $Y=26529 $D=616
M715 vss 11 rb_cb<0> vss hvtnfet l=6e-08 w=8.58e-07 $X=20195 $Y=328 $D=616
M716 vss 12 rb_cb<2> vss hvtnfet l=6e-08 w=8.58e-07 $X=20195 $Y=5316 $D=616
M717 vss 13 rb_mb<0> vss hvtnfet l=6e-08 w=8.58e-07 $X=20195 $Y=6788 $D=616
M718 vss 14 rb_mb<2> vss hvtnfet l=6e-08 w=8.58e-07 $X=20195 $Y=11776 $D=616
M719 vss 15 r_saeb_n vss hvtnfet l=6e-08 w=8.58e-07 $X=20195 $Y=37027 $D=616
M720 vss 16 rt_mb<2> vss hvtnfet l=6e-08 w=8.58e-07 $X=20195 $Y=38499 $D=616
M721 vss 17 rt_mb<0> vss hvtnfet l=6e-08 w=8.58e-07 $X=20195 $Y=43487 $D=616
M722 vss 18 rt_cb<2> vss hvtnfet l=6e-08 w=8.58e-07 $X=20195 $Y=44959 $D=616
M723 vss 19 rt_cb<0> vss hvtnfet l=6e-08 w=8.58e-07 $X=20195 $Y=49947 $D=616
M724 vss 212 1023 vss hvtnfet l=6e-08 w=1.8e-07 $X=20211 $Y=17143 $D=616
M725 vss 280 212 vss hvtnfet l=6e-08 w=1.37e-07 $X=20211 $Y=17812 $D=616
M726 vss 281 185 vss hvtnfet l=6e-08 w=1.37e-07 $X=20211 $Y=18983 $D=616
M727 vss 185 1024 vss hvtnfet l=6e-08 w=1.8e-07 $X=20211 $Y=19609 $D=616
M728 vss 155 1025 vss hvtnfet l=6e-08 w=1.8e-07 $X=20211 $Y=24063 $D=616
M729 vss 282 155 vss hvtnfet l=6e-08 w=1.37e-07 $X=20211 $Y=24732 $D=616
M730 vss 283 145 vss hvtnfet l=6e-08 w=1.37e-07 $X=20211 $Y=25903 $D=616
M731 vss 145 1026 vss hvtnfet l=6e-08 w=1.8e-07 $X=20211 $Y=26529 $D=616
M732 rb_cb<0> 11 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=20455 $Y=328 $D=616
M733 rb_cb<2> 12 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=20455 $Y=5316 $D=616
M734 rb_mb<0> 13 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=20455 $Y=6788 $D=616
M735 rb_mb<2> 14 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=20455 $Y=11776 $D=616
M736 r_saeb_n 15 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=20455 $Y=37027 $D=616
M737 rt_mb<2> 16 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=20455 $Y=38499 $D=616
M738 rt_mb<0> 17 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=20455 $Y=43487 $D=616
M739 rt_cb<2> 18 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=20455 $Y=44959 $D=616
M740 rt_cb<0> 19 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=20455 $Y=49947 $D=616
M741 vss 11 rb_cb<0> vss hvtnfet l=6e-08 w=8.58e-07 $X=20715 $Y=328 $D=616
M742 vss 12 rb_cb<2> vss hvtnfet l=6e-08 w=8.58e-07 $X=20715 $Y=5316 $D=616
M743 vss 13 rb_mb<0> vss hvtnfet l=6e-08 w=8.58e-07 $X=20715 $Y=6788 $D=616
M744 vss 14 rb_mb<2> vss hvtnfet l=6e-08 w=8.58e-07 $X=20715 $Y=11776 $D=616
M745 vss 15 r_saeb_n vss hvtnfet l=6e-08 w=8.58e-07 $X=20715 $Y=37027 $D=616
M746 vss 16 rt_mb<2> vss hvtnfet l=6e-08 w=8.58e-07 $X=20715 $Y=38499 $D=616
M747 vss 17 rt_mb<0> vss hvtnfet l=6e-08 w=8.58e-07 $X=20715 $Y=43487 $D=616
M748 vss 18 rt_cb<2> vss hvtnfet l=6e-08 w=8.58e-07 $X=20715 $Y=44959 $D=616
M749 vss 19 rt_cb<0> vss hvtnfet l=6e-08 w=8.58e-07 $X=20715 $Y=49947 $D=616
M750 10 274 vss vss hvtnfet l=6e-08 w=6e-07 $X=20725 $Y=30899 $D=616
M751 rb_cb<1> 34 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=20975 $Y=328 $D=616
M752 rb_cb<3> 35 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=20975 $Y=5316 $D=616
M753 rb_mb<1> 36 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=20975 $Y=6788 $D=616
M754 rb_mb<3> 37 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=20975 $Y=11776 $D=616
M755 r_clk_dqb 8 vss vss hvtnfet l=6e-08 w=1.26e-06 $X=20975 $Y=22041 $D=616
M756 r_clk_dqb_n 9 vss vss hvtnfet l=6e-08 w=1.26e-06 $X=20975 $Y=29007 $D=616
M757 r_sa_preb_n 51 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=20975 $Y=37027 $D=616
M758 rt_mb<3> 39 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=20975 $Y=38499 $D=616
M759 rt_mb<1> 40 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=20975 $Y=43487 $D=616
M760 rt_cb<3> 41 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=20975 $Y=44959 $D=616
M761 rt_cb<1> 42 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=20975 $Y=49947 $D=616
M762 vss 34 rb_cb<1> vss hvtnfet l=6e-08 w=8.58e-07 $X=21235 $Y=328 $D=616
M763 vss 35 rb_cb<3> vss hvtnfet l=6e-08 w=8.58e-07 $X=21235 $Y=5316 $D=616
M764 vss 36 rb_mb<1> vss hvtnfet l=6e-08 w=8.58e-07 $X=21235 $Y=6788 $D=616
M765 vss 37 rb_mb<3> vss hvtnfet l=6e-08 w=8.58e-07 $X=21235 $Y=11776 $D=616
M766 rb_tm_preb_n 20 vss vss hvtnfet l=6e-08 w=1.287e-06 $X=21235 $Y=13280 $D=616
M767 rt_tm_preb_n 21 vss vss hvtnfet l=6e-08 w=1.287e-06 $X=21235 $Y=20124 $D=616
M768 vss 8 r_clk_dqb vss hvtnfet l=6e-08 w=1.26e-06 $X=21235 $Y=22041 $D=616
M769 vss 9 r_clk_dqb_n vss hvtnfet l=6e-08 w=1.26e-06 $X=21235 $Y=29007 $D=616
M770 r_lweb 10 vss vss hvtnfet l=6e-08 w=1.287e-06 $X=21235 $Y=30897 $D=616
M771 vss 51 r_sa_preb_n vss hvtnfet l=6e-08 w=8.58e-07 $X=21235 $Y=37027 $D=616
M772 vss 39 rt_mb<3> vss hvtnfet l=6e-08 w=8.58e-07 $X=21235 $Y=38499 $D=616
M773 vss 40 rt_mb<1> vss hvtnfet l=6e-08 w=8.58e-07 $X=21235 $Y=43487 $D=616
M774 vss 41 rt_cb<3> vss hvtnfet l=6e-08 w=8.58e-07 $X=21235 $Y=44959 $D=616
M775 vss 42 rt_cb<1> vss hvtnfet l=6e-08 w=8.58e-07 $X=21235 $Y=49947 $D=616
M776 rb_cb<1> 34 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=21495 $Y=328 $D=616
M777 rb_cb<3> 35 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=21495 $Y=5316 $D=616
M778 rb_mb<1> 36 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=21495 $Y=6788 $D=616
M779 rb_mb<3> 37 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=21495 $Y=11776 $D=616
M780 vss 20 rb_tm_preb_n vss hvtnfet l=6e-08 w=1.287e-06 $X=21495 $Y=13280 $D=616
M781 vss 21 rt_tm_preb_n vss hvtnfet l=6e-08 w=1.287e-06 $X=21495 $Y=20124 $D=616
M782 r_clk_dqb 8 vss vss hvtnfet l=6e-08 w=1.26e-06 $X=21495 $Y=22041 $D=616
M783 r_clk_dqb_n 9 vss vss hvtnfet l=6e-08 w=1.26e-06 $X=21495 $Y=29007 $D=616
M784 vss 10 r_lweb vss hvtnfet l=6e-08 w=1.287e-06 $X=21495 $Y=30897 $D=616
M785 r_sa_preb_n 51 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=21495 $Y=37027 $D=616
M786 rt_mb<3> 39 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=21495 $Y=38499 $D=616
M787 rt_mb<1> 40 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=21495 $Y=43487 $D=616
M788 rt_cb<3> 41 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=21495 $Y=44959 $D=616
M789 rt_cb<1> 42 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=21495 $Y=49947 $D=616
M790 vss 289 lb_ca<1> vss hvtnfet l=6e-08 w=8.58e-07 $X=22005 $Y=328 $D=616
M791 vss 290 lb_ca<3> vss hvtnfet l=6e-08 w=8.58e-07 $X=22005 $Y=5316 $D=616
M792 vss 291 lb_ma<1> vss hvtnfet l=6e-08 w=8.58e-07 $X=22005 $Y=6788 $D=616
M793 vss 292 lb_ma<3> vss hvtnfet l=6e-08 w=8.58e-07 $X=22005 $Y=11776 $D=616
M794 lb_tm_prea_n 285 vss vss hvtnfet l=6e-08 w=1.287e-06 $X=22005 $Y=13280 $D=616
M795 lt_tm_prea_n 286 vss vss hvtnfet l=6e-08 w=1.287e-06 $X=22005 $Y=20124 $D=616
M796 vss 287 l_clk_dqa vss hvtnfet l=6e-08 w=1.26e-06 $X=22005 $Y=22041 $D=616
M797 vss 288 l_clk_dqa_n vss hvtnfet l=6e-08 w=1.26e-06 $X=22005 $Y=29007 $D=616
M798 l_lwea 284 vss vss hvtnfet l=6e-08 w=1.287e-06 $X=22005 $Y=30897 $D=616
M799 vss 293 l_sa_prea_n vss hvtnfet l=6e-08 w=8.58e-07 $X=22005 $Y=37027 $D=616
M800 vss 294 lt_ma<3> vss hvtnfet l=6e-08 w=8.58e-07 $X=22005 $Y=38499 $D=616
M801 vss 295 lt_ma<1> vss hvtnfet l=6e-08 w=8.58e-07 $X=22005 $Y=43487 $D=616
M802 vss 296 lt_ca<3> vss hvtnfet l=6e-08 w=8.58e-07 $X=22005 $Y=44959 $D=616
M803 vss 297 lt_ca<1> vss hvtnfet l=6e-08 w=8.58e-07 $X=22005 $Y=49947 $D=616
M804 lb_ca<1> 289 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=22265 $Y=328 $D=616
M805 lb_ca<3> 290 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=22265 $Y=5316 $D=616
M806 lb_ma<1> 291 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=22265 $Y=6788 $D=616
M807 lb_ma<3> 292 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=22265 $Y=11776 $D=616
M808 vss 285 lb_tm_prea_n vss hvtnfet l=6e-08 w=1.287e-06 $X=22265 $Y=13280 $D=616
M809 vss 286 lt_tm_prea_n vss hvtnfet l=6e-08 w=1.287e-06 $X=22265 $Y=20124 $D=616
M810 l_clk_dqa 287 vss vss hvtnfet l=6e-08 w=1.26e-06 $X=22265 $Y=22041 $D=616
M811 l_clk_dqa_n 288 vss vss hvtnfet l=6e-08 w=1.26e-06 $X=22265 $Y=29007 $D=616
M812 vss 284 l_lwea vss hvtnfet l=6e-08 w=1.287e-06 $X=22265 $Y=30897 $D=616
M813 l_sa_prea_n 293 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=22265 $Y=37027 $D=616
M814 lt_ma<3> 294 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=22265 $Y=38499 $D=616
M815 lt_ma<1> 295 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=22265 $Y=43487 $D=616
M816 lt_ca<3> 296 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=22265 $Y=44959 $D=616
M817 lt_ca<1> 297 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=22265 $Y=49947 $D=616
M818 vss 289 lb_ca<1> vss hvtnfet l=6e-08 w=8.58e-07 $X=22525 $Y=328 $D=616
M819 vss 290 lb_ca<3> vss hvtnfet l=6e-08 w=8.58e-07 $X=22525 $Y=5316 $D=616
M820 vss 291 lb_ma<1> vss hvtnfet l=6e-08 w=8.58e-07 $X=22525 $Y=6788 $D=616
M821 vss 292 lb_ma<3> vss hvtnfet l=6e-08 w=8.58e-07 $X=22525 $Y=11776 $D=616
M822 vss 287 l_clk_dqa vss hvtnfet l=6e-08 w=1.26e-06 $X=22525 $Y=22041 $D=616
M823 vss 288 l_clk_dqa_n vss hvtnfet l=6e-08 w=1.26e-06 $X=22525 $Y=29007 $D=616
M824 vss 293 l_sa_prea_n vss hvtnfet l=6e-08 w=8.58e-07 $X=22525 $Y=37027 $D=616
M825 vss 294 lt_ma<3> vss hvtnfet l=6e-08 w=8.58e-07 $X=22525 $Y=38499 $D=616
M826 vss 295 lt_ma<1> vss hvtnfet l=6e-08 w=8.58e-07 $X=22525 $Y=43487 $D=616
M827 vss 296 lt_ca<3> vss hvtnfet l=6e-08 w=8.58e-07 $X=22525 $Y=44959 $D=616
M828 vss 297 lt_ca<1> vss hvtnfet l=6e-08 w=8.58e-07 $X=22525 $Y=49947 $D=616
M829 vss 298 284 vss hvtnfet l=6e-08 w=6e-07 $X=22775 $Y=30899 $D=616
M830 lb_ca<0> 299 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=22785 $Y=328 $D=616
M831 lb_ca<2> 300 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=22785 $Y=5316 $D=616
M832 lb_ma<0> 301 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=22785 $Y=6788 $D=616
M833 lb_ma<2> 302 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=22785 $Y=11776 $D=616
M834 l_saea_n 303 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=22785 $Y=37027 $D=616
M835 lt_ma<2> 304 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=22785 $Y=38499 $D=616
M836 lt_ma<0> 305 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=22785 $Y=43487 $D=616
M837 lt_ca<2> 306 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=22785 $Y=44959 $D=616
M838 lt_ca<0> 307 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=22785 $Y=49947 $D=616
M839 vss 299 lb_ca<0> vss hvtnfet l=6e-08 w=8.58e-07 $X=23045 $Y=328 $D=616
M840 vss 300 lb_ca<2> vss hvtnfet l=6e-08 w=8.58e-07 $X=23045 $Y=5316 $D=616
M841 vss 301 lb_ma<0> vss hvtnfet l=6e-08 w=8.58e-07 $X=23045 $Y=6788 $D=616
M842 vss 302 lb_ma<2> vss hvtnfet l=6e-08 w=8.58e-07 $X=23045 $Y=11776 $D=616
M843 vss 303 l_saea_n vss hvtnfet l=6e-08 w=8.58e-07 $X=23045 $Y=37027 $D=616
M844 vss 304 lt_ma<2> vss hvtnfet l=6e-08 w=8.58e-07 $X=23045 $Y=38499 $D=616
M845 vss 305 lt_ma<0> vss hvtnfet l=6e-08 w=8.58e-07 $X=23045 $Y=43487 $D=616
M846 vss 306 lt_ca<2> vss hvtnfet l=6e-08 w=8.58e-07 $X=23045 $Y=44959 $D=616
M847 vss 307 lt_ca<0> vss hvtnfet l=6e-08 w=8.58e-07 $X=23045 $Y=49947 $D=616
M848 1027 308 vss vss hvtnfet l=6e-08 w=1.8e-07 $X=23289 $Y=17143 $D=616
M849 308 312 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=23289 $Y=17812 $D=616
M850 309 313 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=23289 $Y=18983 $D=616
M851 1028 309 vss vss hvtnfet l=6e-08 w=1.8e-07 $X=23289 $Y=19609 $D=616
M852 1029 310 vss vss hvtnfet l=6e-08 w=1.8e-07 $X=23289 $Y=24063 $D=616
M853 310 314 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=23289 $Y=24732 $D=616
M854 311 315 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=23289 $Y=25903 $D=616
M855 1030 311 vss vss hvtnfet l=6e-08 w=1.8e-07 $X=23289 $Y=26529 $D=616
M856 lb_ca<0> 299 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=23305 $Y=328 $D=616
M857 lb_ca<2> 300 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=23305 $Y=5316 $D=616
M858 lb_ma<0> 301 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=23305 $Y=6788 $D=616
M859 lb_ma<2> 302 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=23305 $Y=11776 $D=616
M860 l_saea_n 303 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=23305 $Y=37027 $D=616
M861 lt_ma<2> 304 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=23305 $Y=38499 $D=616
M862 lt_ma<0> 305 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=23305 $Y=43487 $D=616
M863 lt_ca<2> 306 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=23305 $Y=44959 $D=616
M864 lt_ca<0> 307 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=23305 $Y=49947 $D=616
M865 312 317 1027 vss hvtnfet l=6e-08 w=1.8e-07 $X=23549 $Y=17143 $D=616
M866 vss 312 308 vss hvtnfet l=6e-08 w=1.37e-07 $X=23549 $Y=17812 $D=616
M867 vss 313 309 vss hvtnfet l=6e-08 w=1.37e-07 $X=23549 $Y=18983 $D=616
M868 313 317 1028 vss hvtnfet l=6e-08 w=1.8e-07 $X=23549 $Y=19609 $D=616
M869 314 317 1029 vss hvtnfet l=6e-08 w=1.8e-07 $X=23549 $Y=24063 $D=616
M870 vss 314 310 vss hvtnfet l=6e-08 w=1.37e-07 $X=23549 $Y=24732 $D=616
M871 vss 315 311 vss hvtnfet l=6e-08 w=1.37e-07 $X=23549 $Y=25903 $D=616
M872 315 317 1030 vss hvtnfet l=6e-08 w=1.8e-07 $X=23549 $Y=26529 $D=616
M873 vss 303 l_saea_n vss hvtnfet l=6e-08 w=8.58e-07 $X=23565 $Y=37027 $D=616
M874 l_saea_n 303 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=23825 $Y=37027 $D=616
M875 vss aa<0> 327 vss hvtnfet l=6e-08 w=2.74e-07 $X=23864 $Y=13476 $D=616
M876 vss 324 331 vss hvtnfet l=6e-08 w=2.1e-07 $X=24000 $Y=30918 $D=616
M877 vss 298 332 vss hvtnfet l=6e-08 w=2.1e-07 $X=24000 $Y=32688 $D=616
M878 1031 323 vss vss hvtnfet l=6e-08 w=8.23e-07 $X=24059 $Y=17143 $D=616
M879 1032 323 vss vss hvtnfet l=6e-08 w=8.23e-07 $X=24059 $Y=18966 $D=616
M880 1033 323 vss vss hvtnfet l=6e-08 w=8.23e-07 $X=24059 $Y=24063 $D=616
M881 1034 323 vss vss hvtnfet l=6e-08 w=8.23e-07 $X=24059 $Y=25886 $D=616
M882 b_pxca_n<7> 318 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=24060 $Y=336 $D=616
M883 318 319 vss vss hvtnfet l=6e-08 w=5e-07 $X=24060 $Y=6701 $D=616
M884 319 320 vss vss hvtnfet l=6e-08 w=3e-07 $X=24060 $Y=7831 $D=616
M885 321 320 vss vss hvtnfet l=6e-08 w=3e-07 $X=24060 $Y=43002 $D=616
M886 322 321 vss vss hvtnfet l=6e-08 w=5e-07 $X=24060 $Y=43932 $D=616
M887 t_pxca_n<7> 322 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=24060 $Y=49512 $D=616
M888 709 325 vss vss hvtnfet l=6e-08 w=4.8e-07 $X=24083 $Y=11276 $D=616
M889 710 clka vss vss hvtnfet l=6e-08 w=2.1e-07 $X=24260 $Y=30918 $D=616
M890 711 clka vss vss hvtnfet l=6e-08 w=2.1e-07 $X=24260 $Y=32688 $D=616
M891 vss 318 b_pxca_n<7> vss hvtnfet l=6e-08 w=1.285e-06 $X=24320 $Y=336 $D=616
M892 vss 319 318 vss hvtnfet l=6e-08 w=5e-07 $X=24320 $Y=6701 $D=616
M893 vss 320 319 vss hvtnfet l=6e-08 w=3e-07 $X=24320 $Y=7831 $D=616
M894 vss 320 321 vss hvtnfet l=6e-08 w=3e-07 $X=24320 $Y=43002 $D=616
M895 vss 321 322 vss hvtnfet l=6e-08 w=5e-07 $X=24320 $Y=43932 $D=616
M896 vss 322 t_pxca_n<7> vss hvtnfet l=6e-08 w=1.285e-06 $X=24320 $Y=49512 $D=616
M897 1035 328 1031 vss hvtnfet l=6e-08 w=5.49e-07 $X=24329 $Y=17143 $D=616
M898 1036 328 1032 vss hvtnfet l=6e-08 w=5.49e-07 $X=24329 $Y=19240 $D=616
M899 1037 329 1033 vss hvtnfet l=6e-08 w=5.49e-07 $X=24329 $Y=24063 $D=616
M900 1038 329 1034 vss hvtnfet l=6e-08 w=5.49e-07 $X=24329 $Y=26160 $D=616
M901 vss tm<8> 709 vss hvtnfet l=6e-08 w=4.8e-07 $X=24343 $Y=11276 $D=616
M902 334 327 vss vss hvtnfet l=6e-08 w=2.74e-07 $X=24374 $Y=13476 $D=616
M903 vss tm<5> 264 vss hvtnfet l=6e-08 w=2.74e-07 $X=24518 $Y=39358 $D=616
M904 324 331 710 vss hvtnfet l=6e-08 w=2.1e-07 $X=24520 $Y=30918 $D=616
M905 298 332 711 vss hvtnfet l=6e-08 w=2.1e-07 $X=24520 $Y=32688 $D=616
M906 312 334 1035 vss hvtnfet l=6e-08 w=5.49e-07 $X=24589 $Y=17143 $D=616
M907 313 327 1036 vss hvtnfet l=6e-08 w=5.49e-07 $X=24589 $Y=19240 $D=616
M908 314 334 1037 vss hvtnfet l=6e-08 w=5.49e-07 $X=24589 $Y=24063 $D=616
M909 315 327 1038 vss hvtnfet l=6e-08 w=5.49e-07 $X=24589 $Y=26160 $D=616
M910 714 340 324 vss hvtnfet l=6e-08 w=3.2e-07 $X=24780 $Y=30918 $D=616
M911 715 340 298 vss hvtnfet l=6e-08 w=3.2e-07 $X=24780 $Y=32578 $D=616
M912 b_pxca_n<6> 335 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=24830 $Y=336 $D=616
M913 335 336 vss vss hvtnfet l=6e-08 w=5e-07 $X=24830 $Y=6701 $D=616
M914 336 337 vss vss hvtnfet l=6e-08 w=3e-07 $X=24830 $Y=7831 $D=616
M915 338 337 vss vss hvtnfet l=6e-08 w=3e-07 $X=24830 $Y=43002 $D=616
M916 339 338 vss vss hvtnfet l=6e-08 w=5e-07 $X=24830 $Y=43932 $D=616
M917 t_pxca_n<6> 339 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=24830 $Y=49512 $D=616
M918 718 tm<8> vss vss hvtnfet l=6e-08 w=4.8e-07 $X=24853 $Y=11276 $D=616
M919 vss 264 376 vss hvtnfet l=6e-08 w=2e-07 $X=24874 $Y=37147 $D=616
M920 vss aa<1> 329 vss hvtnfet l=6e-08 w=2.74e-07 $X=24884 $Y=13476 $D=616
M921 vss aa<4> 714 vss hvtnfet l=6e-08 w=3.2e-07 $X=25040 $Y=30918 $D=616
M922 vss wena 715 vss hvtnfet l=6e-08 w=3.2e-07 $X=25040 $Y=32578 $D=616
M923 vss 335 b_pxca_n<6> vss hvtnfet l=6e-08 w=1.285e-06 $X=25090 $Y=336 $D=616
M924 vss 336 335 vss hvtnfet l=6e-08 w=5e-07 $X=25090 $Y=6701 $D=616
M925 vss 337 336 vss hvtnfet l=6e-08 w=3e-07 $X=25090 $Y=7831 $D=616
M926 vss 337 338 vss hvtnfet l=6e-08 w=3e-07 $X=25090 $Y=43002 $D=616
M927 vss 338 339 vss hvtnfet l=6e-08 w=5e-07 $X=25090 $Y=43932 $D=616
M928 vss 339 t_pxca_n<6> vss hvtnfet l=6e-08 w=1.285e-06 $X=25090 $Y=49512 $D=616
M929 vss tm<9> 718 vss hvtnfet l=6e-08 w=4.8e-07 $X=25113 $Y=11276 $D=616
M930 376 wena vss vss hvtnfet l=6e-08 w=2e-07 $X=25134 $Y=37147 $D=616
M931 328 329 vss vss hvtnfet l=6e-08 w=2.74e-07 $X=25394 $Y=13476 $D=616
M932 b_pxca_n<5> 345 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=25600 $Y=336 $D=616
M933 345 346 vss vss hvtnfet l=6e-08 w=5e-07 $X=25600 $Y=6701 $D=616
M934 346 347 vss vss hvtnfet l=6e-08 w=3e-07 $X=25600 $Y=7831 $D=616
M935 348 347 vss vss hvtnfet l=6e-08 w=3e-07 $X=25600 $Y=43002 $D=616
M936 349 348 vss vss hvtnfet l=6e-08 w=5e-07 $X=25600 $Y=43932 $D=616
M937 t_pxca_n<5> 349 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=25600 $Y=49512 $D=616
M938 1039 337 vss vss hvtnfet l=6e-08 w=1.8e-07 $X=25609 $Y=17143 $D=616
M939 1040 320 vss vss hvtnfet l=6e-08 w=1.8e-07 $X=25609 $Y=19609 $D=616
M940 1041 350 vss vss hvtnfet l=6e-08 w=1.8e-07 $X=25609 $Y=24063 $D=616
M941 1042 351 vss vss hvtnfet l=6e-08 w=1.8e-07 $X=25609 $Y=26529 $D=616
M942 721 tm<9> vss vss hvtnfet l=6e-08 w=4.8e-07 $X=25623 $Y=11276 $D=616
M943 337 352 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=25624 $Y=17812 $D=616
M944 320 353 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=25624 $Y=18983 $D=616
M945 350 354 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=25624 $Y=24732 $D=616
M946 351 355 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=25624 $Y=25903 $D=616
M947 vss clka 340 vss hvtnfet l=6e-08 w=4.5e-07 $X=25854 $Y=30668 $D=616
M948 vss 345 b_pxca_n<5> vss hvtnfet l=6e-08 w=1.285e-06 $X=25860 $Y=336 $D=616
M949 vss 346 345 vss hvtnfet l=6e-08 w=5e-07 $X=25860 $Y=6701 $D=616
M950 vss 347 346 vss hvtnfet l=6e-08 w=3e-07 $X=25860 $Y=7831 $D=616
M951 vss 347 348 vss hvtnfet l=6e-08 w=3e-07 $X=25860 $Y=43002 $D=616
M952 vss 348 349 vss hvtnfet l=6e-08 w=5e-07 $X=25860 $Y=43932 $D=616
M953 vss 349 t_pxca_n<5> vss hvtnfet l=6e-08 w=1.285e-06 $X=25860 $Y=49512 $D=616
M954 352 317 1039 vss hvtnfet l=6e-08 w=1.8e-07 $X=25869 $Y=17143 $D=616
M955 353 317 1040 vss hvtnfet l=6e-08 w=1.8e-07 $X=25869 $Y=19609 $D=616
M956 354 317 1041 vss hvtnfet l=6e-08 w=1.8e-07 $X=25869 $Y=24063 $D=616
M957 355 317 1042 vss hvtnfet l=6e-08 w=1.8e-07 $X=25869 $Y=26529 $D=616
M958 vss 366 721 vss hvtnfet l=6e-08 w=4.8e-07 $X=25883 $Y=11276 $D=616
M959 vss 352 337 vss hvtnfet l=6e-08 w=1.37e-07 $X=25884 $Y=17812 $D=616
M960 vss 353 320 vss hvtnfet l=6e-08 w=1.37e-07 $X=25884 $Y=18983 $D=616
M961 vss 354 350 vss hvtnfet l=6e-08 w=1.37e-07 $X=25884 $Y=24732 $D=616
M962 vss 355 351 vss hvtnfet l=6e-08 w=1.37e-07 $X=25884 $Y=25903 $D=616
M963 vss 356 363 vss hvtnfet l=6e-08 w=2.1e-07 $X=26138 $Y=37277 $D=616
M964 b_pxca_n<4> 357 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=26370 $Y=336 $D=616
M965 357 358 vss vss hvtnfet l=6e-08 w=5e-07 $X=26370 $Y=6701 $D=616
M966 358 359 vss vss hvtnfet l=6e-08 w=3e-07 $X=26370 $Y=7831 $D=616
M967 360 359 vss vss hvtnfet l=6e-08 w=3e-07 $X=26370 $Y=43002 $D=616
M968 361 360 vss vss hvtnfet l=6e-08 w=5e-07 $X=26370 $Y=43932 $D=616
M969 t_pxca_n<4> 361 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=26370 $Y=49512 $D=616
M970 729 123 733 vss hvtnfet l=6e-08 w=6e-07 $X=26374 $Y=30668 $D=616
M971 1043 323 vss vss hvtnfet l=6e-08 w=8.23e-07 $X=26379 $Y=17143 $D=616
M972 1044 323 vss vss hvtnfet l=6e-08 w=8.23e-07 $X=26379 $Y=18966 $D=616
M973 1045 323 vss vss hvtnfet l=6e-08 w=8.23e-07 $X=26379 $Y=24063 $D=616
M974 1046 323 vss vss hvtnfet l=6e-08 w=8.23e-07 $X=26379 $Y=25886 $D=616
M975 vss 366 727 vss hvtnfet l=6e-08 w=4.8e-07 $X=26393 $Y=11276 $D=616
M976 724 362 vss vss hvtnfet l=6e-08 w=2.1e-07 $X=26398 $Y=37277 $D=616
M977 vss 357 b_pxca_n<4> vss hvtnfet l=6e-08 w=1.285e-06 $X=26630 $Y=336 $D=616
M978 vss 358 357 vss hvtnfet l=6e-08 w=5e-07 $X=26630 $Y=6701 $D=616
M979 vss 359 358 vss hvtnfet l=6e-08 w=3e-07 $X=26630 $Y=7831 $D=616
M980 vss 359 360 vss hvtnfet l=6e-08 w=3e-07 $X=26630 $Y=43002 $D=616
M981 vss 360 361 vss hvtnfet l=6e-08 w=5e-07 $X=26630 $Y=43932 $D=616
M982 vss 361 t_pxca_n<4> vss hvtnfet l=6e-08 w=1.285e-06 $X=26630 $Y=49512 $D=616
M983 733 123 729 vss hvtnfet l=6e-08 w=6e-07 $X=26634 $Y=30668 $D=616
M984 1047 364 1043 vss hvtnfet l=6e-08 w=5.49e-07 $X=26649 $Y=17417 $D=616
M985 1048 364 1044 vss hvtnfet l=6e-08 w=5.49e-07 $X=26649 $Y=18966 $D=616
M986 1049 365 1045 vss hvtnfet l=6e-08 w=5.49e-07 $X=26649 $Y=24337 $D=616
M987 1050 365 1046 vss hvtnfet l=6e-08 w=5.49e-07 $X=26649 $Y=25886 $D=616
M988 727 325 vss vss hvtnfet l=6e-08 w=4.8e-07 $X=26653 $Y=11276 $D=616
M989 356 363 724 vss hvtnfet l=6e-08 w=2.1e-07 $X=26658 $Y=37277 $D=616
M990 vss tm<7> 726 vss hvtnfet l=6e-08 w=2.74e-07 $X=26820 $Y=39358 $D=616
M991 728 123 vss vss hvtnfet l=6e-08 w=3.2e-07 $X=26839 $Y=32578 $D=616
M992 vss 123 733 vss hvtnfet l=6e-08 w=6e-07 $X=26894 $Y=30668 $D=616
M993 1051 369 1047 vss hvtnfet l=6e-08 w=5.49e-07 $X=26909 $Y=17417 $D=616
M994 1052 369 1048 vss hvtnfet l=6e-08 w=5.49e-07 $X=26909 $Y=18966 $D=616
M995 1053 369 1049 vss hvtnfet l=6e-08 w=5.49e-07 $X=26909 $Y=24337 $D=616
M996 1054 369 1050 vss hvtnfet l=6e-08 w=5.49e-07 $X=26909 $Y=25886 $D=616
M997 730 368 356 vss hvtnfet l=6e-08 w=3.2e-07 $X=26918 $Y=37277 $D=616
M998 vss aa<10> 374 vss hvtnfet l=6e-08 w=2.74e-07 $X=26924 $Y=13476 $D=616
M999 379 123 728 vss hvtnfet l=6e-08 w=3.2e-07 $X=27099 $Y=32578 $D=616
M1000 b_pxca_n<3> 370 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=27140 $Y=336 $D=616
M1001 370 371 vss vss hvtnfet l=6e-08 w=5e-07 $X=27140 $Y=6701 $D=616
M1002 371 351 vss vss hvtnfet l=6e-08 w=3e-07 $X=27140 $Y=7831 $D=616
M1003 372 351 vss vss hvtnfet l=6e-08 w=3e-07 $X=27140 $Y=43002 $D=616
M1004 373 372 vss vss hvtnfet l=6e-08 w=5e-07 $X=27140 $Y=43932 $D=616
M1005 t_pxca_n<3> 373 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=27140 $Y=49512 $D=616
M1006 733 123 vss vss hvtnfet l=6e-08 w=6e-07 $X=27154 $Y=30668 $D=616
M1007 vss tm<9> 325 vss hvtnfet l=7e-08 w=3.2e-07 $X=27163 $Y=11276 $D=616
M1008 352 374 1051 vss hvtnfet l=6e-08 w=5.49e-07 $X=27169 $Y=17417 $D=616
M1009 353 375 1052 vss hvtnfet l=6e-08 w=5.49e-07 $X=27169 $Y=18966 $D=616
M1010 354 374 1053 vss hvtnfet l=6e-08 w=5.49e-07 $X=27169 $Y=24337 $D=616
M1011 355 375 1054 vss hvtnfet l=6e-08 w=5.49e-07 $X=27169 $Y=25886 $D=616
M1012 vss 376 730 vss hvtnfet l=6e-08 w=3.2e-07 $X=27178 $Y=37277 $D=616
M1013 375 374 vss vss hvtnfet l=6e-08 w=2.74e-07 $X=27184 $Y=13476 $D=616
M1014 734 377 379 vss hvtnfet l=6e-08 w=2.1e-07 $X=27359 $Y=32688 $D=616
M1015 vss 370 b_pxca_n<3> vss hvtnfet l=6e-08 w=1.285e-06 $X=27400 $Y=336 $D=616
M1016 vss 371 370 vss hvtnfet l=6e-08 w=5e-07 $X=27400 $Y=6701 $D=616
M1017 vss 351 371 vss hvtnfet l=6e-08 w=3e-07 $X=27400 $Y=7831 $D=616
M1018 vss 351 372 vss hvtnfet l=6e-08 w=3e-07 $X=27400 $Y=43002 $D=616
M1019 vss 372 373 vss hvtnfet l=6e-08 w=5e-07 $X=27400 $Y=43932 $D=616
M1020 vss 373 t_pxca_n<3> vss hvtnfet l=6e-08 w=1.285e-06 $X=27400 $Y=49512 $D=616
M1021 366 tm<8> vss vss hvtnfet l=7e-08 w=3.2e-07 $X=27433 $Y=11276 $D=616
M1022 vss 131 734 vss hvtnfet l=6e-08 w=2.1e-07 $X=27619 $Y=32688 $D=616
M1023 vss tm<1> 735 vss hvtnfet l=6e-08 w=2.74e-07 $X=27620 $Y=39358 $D=616
M1024 vss 380 369 vss hvtnfet l=6e-08 w=2.74e-07 $X=27784 $Y=13476 $D=616
M1025 737 362 386 vss hvtnfet l=6e-08 w=4e-07 $X=27858 $Y=37045 $D=616
M1026 377 379 vss vss hvtnfet l=6e-08 w=2.1e-07 $X=27879 $Y=32688 $D=616
M1027 b_pxca_n<2> 381 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=27910 $Y=336 $D=616
M1028 381 382 vss vss hvtnfet l=6e-08 w=5e-07 $X=27910 $Y=6701 $D=616
M1029 382 350 vss vss hvtnfet l=6e-08 w=3e-07 $X=27910 $Y=7831 $D=616
M1030 383 350 vss vss hvtnfet l=6e-08 w=3e-07 $X=27910 $Y=43002 $D=616
M1031 384 383 vss vss hvtnfet l=6e-08 w=5e-07 $X=27910 $Y=43932 $D=616
M1032 t_pxca_n<2> 384 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=27910 $Y=49512 $D=616
M1033 vss 323 317 vss hvtnfet l=6e-08 w=7e-07 $X=27924 $Y=30668 $D=616
M1034 380 aa<11> vss vss hvtnfet l=6e-08 w=2.74e-07 $X=28044 $Y=13476 $D=616
M1035 vss 356 737 vss hvtnfet l=6e-08 w=4e-07 $X=28118 $Y=37045 $D=616
M1036 vss 381 b_pxca_n<2> vss hvtnfet l=6e-08 w=1.285e-06 $X=28170 $Y=336 $D=616
M1037 vss 382 381 vss hvtnfet l=6e-08 w=5e-07 $X=28170 $Y=6701 $D=616
M1038 vss 350 382 vss hvtnfet l=6e-08 w=3e-07 $X=28170 $Y=7831 $D=616
M1039 vss 350 383 vss hvtnfet l=6e-08 w=3e-07 $X=28170 $Y=43002 $D=616
M1040 vss 383 384 vss hvtnfet l=6e-08 w=5e-07 $X=28170 $Y=43932 $D=616
M1041 vss 384 t_pxca_n<2> vss hvtnfet l=6e-08 w=1.285e-06 $X=28170 $Y=49512 $D=616
M1042 317 323 vss vss hvtnfet l=6e-08 w=7e-07 $X=28184 $Y=30668 $D=616
M1043 vss 392 541 vss hvtnfet l=6e-08 w=2e-07 $X=28514 $Y=11276 $D=616
M1044 vss 393 544 vss hvtnfet l=6e-08 w=2e-07 $X=28514 $Y=39657 $D=616
M1045 494 386 vss vss hvtnfet l=6e-08 w=2e-07 $X=28628 $Y=37045 $D=616
M1046 b_pxca_n<1> 387 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=28680 $Y=336 $D=616
M1047 387 388 vss vss hvtnfet l=6e-08 w=5e-07 $X=28680 $Y=6701 $D=616
M1048 388 389 vss vss hvtnfet l=6e-08 w=3e-07 $X=28680 $Y=7831 $D=616
M1049 390 389 vss vss hvtnfet l=6e-08 w=3e-07 $X=28680 $Y=43002 $D=616
M1050 391 390 vss vss hvtnfet l=6e-08 w=5e-07 $X=28680 $Y=43932 $D=616
M1051 t_pxca_n<1> 391 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=28680 $Y=49512 $D=616
M1052 742 123 vss vss hvtnfet l=6e-08 w=6e-07 $X=28704 $Y=30668 $D=616
M1053 vss 387 b_pxca_n<1> vss hvtnfet l=6e-08 w=1.285e-06 $X=28940 $Y=336 $D=616
M1054 vss 388 387 vss hvtnfet l=6e-08 w=5e-07 $X=28940 $Y=6701 $D=616
M1055 vss 389 388 vss hvtnfet l=6e-08 w=3e-07 $X=28940 $Y=7831 $D=616
M1056 vss 389 390 vss hvtnfet l=6e-08 w=3e-07 $X=28940 $Y=43002 $D=616
M1057 vss 390 391 vss hvtnfet l=6e-08 w=5e-07 $X=28940 $Y=43932 $D=616
M1058 vss 391 t_pxca_n<1> vss hvtnfet l=6e-08 w=1.285e-06 $X=28940 $Y=49512 $D=616
M1059 1055 374 407 vss hvtnfet l=6e-08 w=5.49e-07 $X=29009 $Y=17417 $D=616
M1060 1056 375 408 vss hvtnfet l=6e-08 w=5.49e-07 $X=29009 $Y=18966 $D=616
M1061 1057 374 409 vss hvtnfet l=6e-08 w=5.49e-07 $X=29009 $Y=24337 $D=616
M1062 1058 375 410 vss hvtnfet l=6e-08 w=5.49e-07 $X=29009 $Y=25886 $D=616
M1063 1059 308 vss vss hvtnfet l=6e-08 w=4.11e-07 $X=29024 $Y=11276 $D=616
M1064 1060 308 vss vss hvtnfet l=6e-08 w=4.11e-07 $X=29024 $Y=39446 $D=616
M1065 vss aa<12> 365 vss hvtnfet l=6e-08 w=2.74e-07 $X=29054 $Y=13476 $D=616
M1066 1061 380 1055 vss hvtnfet l=6e-08 w=5.49e-07 $X=29269 $Y=17417 $D=616
M1067 1062 380 1056 vss hvtnfet l=6e-08 w=5.49e-07 $X=29269 $Y=18966 $D=616
M1068 1063 380 1057 vss hvtnfet l=6e-08 w=5.49e-07 $X=29269 $Y=24337 $D=616
M1069 1064 380 1058 vss hvtnfet l=6e-08 w=5.49e-07 $X=29269 $Y=25886 $D=616
M1070 392 dwla<1> 1059 vss hvtnfet l=6e-08 w=4.11e-07 $X=29284 $Y=11276 $D=616
M1071 393 dwla<0> 1060 vss hvtnfet l=6e-08 w=4.11e-07 $X=29284 $Y=39446 $D=616
M1072 vss 395 403 vss hvtnfet l=6e-08 w=2e-07 $X=29298 $Y=32533 $D=616
M1073 b_pxca_n<0> 396 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=29450 $Y=336 $D=616
M1074 396 397 vss vss hvtnfet l=6e-08 w=5e-07 $X=29450 $Y=6701 $D=616
M1075 397 398 vss vss hvtnfet l=6e-08 w=3e-07 $X=29450 $Y=7831 $D=616
M1076 399 398 vss vss hvtnfet l=6e-08 w=3e-07 $X=29450 $Y=43002 $D=616
M1077 400 399 vss vss hvtnfet l=6e-08 w=5e-07 $X=29450 $Y=43932 $D=616
M1078 t_pxca_n<0> 400 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=29450 $Y=49512 $D=616
M1079 1065 364 1061 vss hvtnfet l=6e-08 w=5.49e-07 $X=29529 $Y=17417 $D=616
M1080 1066 364 1062 vss hvtnfet l=6e-08 w=5.49e-07 $X=29529 $Y=18966 $D=616
M1081 1067 365 1063 vss hvtnfet l=6e-08 w=5.49e-07 $X=29529 $Y=24337 $D=616
M1082 1068 365 1064 vss hvtnfet l=6e-08 w=5.49e-07 $X=29529 $Y=25886 $D=616
M1083 403 405 vss vss hvtnfet l=6e-08 w=2e-07 $X=29558 $Y=32533 $D=616
M1084 364 365 vss vss hvtnfet l=6e-08 w=2.74e-07 $X=29564 $Y=13476 $D=616
M1085 vss 404 395 vss hvtnfet l=6e-08 w=3.5e-07 $X=29621 $Y=30853 $D=616
M1086 vss 396 b_pxca_n<0> vss hvtnfet l=6e-08 w=1.285e-06 $X=29710 $Y=336 $D=616
M1087 vss 397 396 vss hvtnfet l=6e-08 w=5e-07 $X=29710 $Y=6701 $D=616
M1088 vss 398 397 vss hvtnfet l=6e-08 w=3e-07 $X=29710 $Y=7831 $D=616
M1089 vss 398 399 vss hvtnfet l=6e-08 w=3e-07 $X=29710 $Y=43002 $D=616
M1090 vss 399 400 vss hvtnfet l=6e-08 w=5e-07 $X=29710 $Y=43932 $D=616
M1091 vss 400 t_pxca_n<0> vss hvtnfet l=6e-08 w=1.285e-06 $X=29710 $Y=49512 $D=616
M1092 456 403 vss vss hvtnfet l=6e-08 w=6e-07 $X=29747 $Y=37037 $D=616
M1093 vss 323 1065 vss hvtnfet l=6e-08 w=8.23e-07 $X=29799 $Y=17143 $D=616
M1094 vss 323 1066 vss hvtnfet l=6e-08 w=8.23e-07 $X=29799 $Y=18966 $D=616
M1095 vss 323 1067 vss hvtnfet l=6e-08 w=8.23e-07 $X=29799 $Y=24063 $D=616
M1096 vss 323 1068 vss hvtnfet l=6e-08 w=8.23e-07 $X=29799 $Y=25886 $D=616
M1097 404 406 vss vss hvtnfet l=2.5e-07 w=3.5e-07 $X=29881 $Y=30853 $D=616
M1098 405 tm<7> vss vss hvtnfet l=6e-08 w=2e-07 $X=30068 $Y=32533 $D=616
M1099 dbl_pd_n<3> 131 vss vss hvtnfet l=6e-08 w=2.14e-07 $X=30204 $Y=13361 $D=616
M1100 b_pxba_n<7> 411 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=30220 $Y=336 $D=616
M1101 411 412 vss vss hvtnfet l=6e-08 w=5e-07 $X=30220 $Y=6701 $D=616
M1102 412 413 vss vss hvtnfet l=6e-08 w=3e-07 $X=30220 $Y=7831 $D=616
M1103 414 413 vss vss hvtnfet l=6e-08 w=3e-07 $X=30220 $Y=43002 $D=616
M1104 415 414 vss vss hvtnfet l=6e-08 w=5e-07 $X=30220 $Y=43932 $D=616
M1105 t_pxba_n<7> 415 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=30220 $Y=49512 $D=616
M1106 359 407 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=30294 $Y=17812 $D=616
M1107 347 408 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=30294 $Y=18983 $D=616
M1108 398 409 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=30294 $Y=24732 $D=616
M1109 389 410 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=30294 $Y=25903 $D=616
M1110 1069 317 407 vss hvtnfet l=6e-08 w=1.8e-07 $X=30309 $Y=17143 $D=616
M1111 1070 317 408 vss hvtnfet l=6e-08 w=1.8e-07 $X=30309 $Y=19609 $D=616
M1112 1071 317 409 vss hvtnfet l=6e-08 w=1.8e-07 $X=30309 $Y=24063 $D=616
M1113 1072 317 410 vss hvtnfet l=6e-08 w=1.8e-07 $X=30309 $Y=26529 $D=616
M1114 vss 131 dbl_pd_n<3> vss hvtnfet l=6e-08 w=2.14e-07 $X=30464 $Y=13361 $D=616
M1115 vss 411 b_pxba_n<7> vss hvtnfet l=6e-08 w=1.285e-06 $X=30480 $Y=336 $D=616
M1116 vss 412 411 vss hvtnfet l=6e-08 w=5e-07 $X=30480 $Y=6701 $D=616
M1117 vss 413 412 vss hvtnfet l=6e-08 w=3e-07 $X=30480 $Y=7831 $D=616
M1118 vss 413 414 vss hvtnfet l=6e-08 w=3e-07 $X=30480 $Y=43002 $D=616
M1119 vss 414 415 vss hvtnfet l=6e-08 w=5e-07 $X=30480 $Y=43932 $D=616
M1120 vss 415 t_pxba_n<7> vss hvtnfet l=6e-08 w=1.285e-06 $X=30480 $Y=49512 $D=616
M1121 456 416 vss vss hvtnfet l=6e-08 w=6e-07 $X=30527 $Y=37037 $D=616
M1122 vss 407 359 vss hvtnfet l=6e-08 w=1.37e-07 $X=30554 $Y=17812 $D=616
M1123 vss 408 347 vss hvtnfet l=6e-08 w=1.37e-07 $X=30554 $Y=18983 $D=616
M1124 vss 409 398 vss hvtnfet l=6e-08 w=1.37e-07 $X=30554 $Y=24732 $D=616
M1125 vss 410 389 vss hvtnfet l=6e-08 w=1.37e-07 $X=30554 $Y=25903 $D=616
M1126 vss 359 1069 vss hvtnfet l=6e-08 w=1.8e-07 $X=30569 $Y=17143 $D=616
M1127 vss 347 1070 vss hvtnfet l=6e-08 w=1.8e-07 $X=30569 $Y=19609 $D=616
M1128 vss 398 1071 vss hvtnfet l=6e-08 w=1.8e-07 $X=30569 $Y=24063 $D=616
M1129 vss 389 1072 vss hvtnfet l=6e-08 w=1.8e-07 $X=30569 $Y=26529 $D=616
M1130 1073 dwla<1> 426 vss hvtnfet l=6e-08 w=4.11e-07 $X=30584 $Y=11276 $D=616
M1131 1074 dwla<0> 427 vss hvtnfet l=6e-08 w=4.11e-07 $X=30584 $Y=39446 $D=616
M1132 vss 406 416 vss hvtnfet l=6e-08 w=2e-07 $X=30644 $Y=32533 $D=616
M1133 dbl_pd_n<3> 131 vss vss hvtnfet l=6e-08 w=2.14e-07 $X=30724 $Y=13361 $D=616
M1134 vss 417 406 vss hvtnfet l=6e-08 w=3.5e-07 $X=30741 $Y=30853 $D=616
M1135 vss 309 1073 vss hvtnfet l=6e-08 w=4.11e-07 $X=30844 $Y=11276 $D=616
M1136 vss 309 1074 vss hvtnfet l=6e-08 w=4.11e-07 $X=30844 $Y=39446 $D=616
M1137 416 423 vss vss hvtnfet l=6e-08 w=2e-07 $X=30904 $Y=32533 $D=616
M1138 b_pxba_n<6> 418 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=30990 $Y=336 $D=616
M1139 418 419 vss vss hvtnfet l=6e-08 w=5e-07 $X=30990 $Y=6701 $D=616
M1140 419 420 vss vss hvtnfet l=6e-08 w=3e-07 $X=30990 $Y=7831 $D=616
M1141 421 420 vss vss hvtnfet l=6e-08 w=3e-07 $X=30990 $Y=43002 $D=616
M1142 422 421 vss vss hvtnfet l=6e-08 w=5e-07 $X=30990 $Y=43932 $D=616
M1143 t_pxba_n<6> 422 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=30990 $Y=49512 $D=616
M1144 417 368 vss vss hvtnfet l=2.5e-07 w=3.5e-07 $X=31001 $Y=30853 $D=616
M1145 1075 420 vss vss hvtnfet l=6e-08 w=1.8e-07 $X=31079 $Y=17143 $D=616
M1146 1076 413 vss vss hvtnfet l=6e-08 w=1.8e-07 $X=31079 $Y=19609 $D=616
M1147 1077 424 vss vss hvtnfet l=6e-08 w=1.8e-07 $X=31079 $Y=24063 $D=616
M1148 1078 425 vss vss hvtnfet l=6e-08 w=1.8e-07 $X=31079 $Y=26529 $D=616
M1149 420 428 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=31094 $Y=17812 $D=616
M1150 413 429 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=31094 $Y=18983 $D=616
M1151 424 430 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=31094 $Y=24732 $D=616
M1152 425 431 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=31094 $Y=25903 $D=616
M1153 dbl_pd_n<1> tm<1> vss vss hvtnfet l=6e-08 w=2.14e-07 $X=31234 $Y=13361 $D=616
M1154 vss 418 b_pxba_n<6> vss hvtnfet l=6e-08 w=1.285e-06 $X=31250 $Y=336 $D=616
M1155 vss 419 418 vss hvtnfet l=6e-08 w=5e-07 $X=31250 $Y=6701 $D=616
M1156 vss 420 419 vss hvtnfet l=6e-08 w=3e-07 $X=31250 $Y=7831 $D=616
M1157 vss 420 421 vss hvtnfet l=6e-08 w=3e-07 $X=31250 $Y=43002 $D=616
M1158 vss 421 422 vss hvtnfet l=6e-08 w=5e-07 $X=31250 $Y=43932 $D=616
M1159 vss 422 t_pxba_n<6> vss hvtnfet l=6e-08 w=1.285e-06 $X=31250 $Y=49512 $D=616
M1160 456 362 vss vss hvtnfet l=6e-08 w=6e-07 $X=31307 $Y=37037 $D=616
M1161 428 317 1075 vss hvtnfet l=6e-08 w=1.8e-07 $X=31339 $Y=17143 $D=616
M1162 429 317 1076 vss hvtnfet l=6e-08 w=1.8e-07 $X=31339 $Y=19609 $D=616
M1163 430 317 1077 vss hvtnfet l=6e-08 w=1.8e-07 $X=31339 $Y=24063 $D=616
M1164 431 317 1078 vss hvtnfet l=6e-08 w=1.8e-07 $X=31339 $Y=26529 $D=616
M1165 556 426 vss vss hvtnfet l=6e-08 w=2e-07 $X=31354 $Y=11276 $D=616
M1166 vss 428 420 vss hvtnfet l=6e-08 w=1.37e-07 $X=31354 $Y=17812 $D=616
M1167 vss 429 413 vss hvtnfet l=6e-08 w=1.37e-07 $X=31354 $Y=18983 $D=616
M1168 vss 430 424 vss hvtnfet l=6e-08 w=1.37e-07 $X=31354 $Y=24732 $D=616
M1169 vss 431 425 vss hvtnfet l=6e-08 w=1.37e-07 $X=31354 $Y=25903 $D=616
M1170 558 427 vss vss hvtnfet l=6e-08 w=2e-07 $X=31354 $Y=39657 $D=616
M1171 vss 173 423 vss hvtnfet l=6e-08 w=2e-07 $X=31414 $Y=32533 $D=616
M1172 vss tm<1> dbl_pd_n<1> vss hvtnfet l=6e-08 w=2.14e-07 $X=31494 $Y=13361 $D=616
M1173 dbl_pd_n<1> tm<1> vss vss hvtnfet l=6e-08 w=2.14e-07 $X=31754 $Y=13361 $D=616
M1174 b_pxba_n<5> 432 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=31760 $Y=336 $D=616
M1175 432 433 vss vss hvtnfet l=6e-08 w=5e-07 $X=31760 $Y=6701 $D=616
M1176 433 434 vss vss hvtnfet l=6e-08 w=3e-07 $X=31760 $Y=7831 $D=616
M1177 435 434 vss vss hvtnfet l=6e-08 w=3e-07 $X=31760 $Y=43002 $D=616
M1178 436 435 vss vss hvtnfet l=6e-08 w=5e-07 $X=31760 $Y=43932 $D=616
M1179 t_pxba_n<5> 436 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=31760 $Y=49512 $D=616
M1180 vss 368 362 vss hvtnfet l=6e-08 w=2e-07 $X=31761 $Y=31098 $D=616
M1181 1079 323 vss vss hvtnfet l=6e-08 w=8.23e-07 $X=31849 $Y=17143 $D=616
M1182 1080 323 vss vss hvtnfet l=6e-08 w=8.23e-07 $X=31849 $Y=18966 $D=616
M1183 1081 323 vss vss hvtnfet l=6e-08 w=8.23e-07 $X=31849 $Y=24063 $D=616
M1184 1082 323 vss vss hvtnfet l=6e-08 w=8.23e-07 $X=31849 $Y=25886 $D=616
M1185 vss 437 540 vss hvtnfet l=6e-08 w=2e-07 $X=31864 $Y=11276 $D=616
M1186 vss 438 545 vss hvtnfet l=6e-08 w=2e-07 $X=31864 $Y=39657 $D=616
M1187 vss 432 b_pxba_n<5> vss hvtnfet l=6e-08 w=1.285e-06 $X=32020 $Y=336 $D=616
M1188 vss 433 432 vss hvtnfet l=6e-08 w=5e-07 $X=32020 $Y=6701 $D=616
M1189 vss 434 433 vss hvtnfet l=6e-08 w=3e-07 $X=32020 $Y=7831 $D=616
M1190 vss 434 435 vss hvtnfet l=6e-08 w=3e-07 $X=32020 $Y=43002 $D=616
M1191 vss 435 436 vss hvtnfet l=6e-08 w=5e-07 $X=32020 $Y=43932 $D=616
M1192 vss 436 t_pxba_n<5> vss hvtnfet l=6e-08 w=1.285e-06 $X=32020 $Y=49512 $D=616
M1193 1083 439 1079 vss hvtnfet l=6e-08 w=5.49e-07 $X=32119 $Y=17417 $D=616
M1194 1084 439 1080 vss hvtnfet l=6e-08 w=5.49e-07 $X=32119 $Y=18966 $D=616
M1195 1085 440 1081 vss hvtnfet l=6e-08 w=5.49e-07 $X=32119 $Y=24337 $D=616
M1196 1086 440 1082 vss hvtnfet l=6e-08 w=5.49e-07 $X=32119 $Y=25886 $D=616
M1197 dwla<1> 442 vss vss hvtnfet l=6e-08 w=3e-07 $X=32271 $Y=31098 $D=616
M1198 497 442 vss vss hvtnfet l=6e-08 w=3e-07 $X=32271 $Y=37457 $D=616
M1199 1087 310 vss vss hvtnfet l=6e-08 w=4.11e-07 $X=32374 $Y=11276 $D=616
M1200 1088 310 vss vss hvtnfet l=6e-08 w=4.11e-07 $X=32374 $Y=39446 $D=616
M1201 1089 443 1083 vss hvtnfet l=6e-08 w=5.49e-07 $X=32379 $Y=17417 $D=616
M1202 1090 443 1084 vss hvtnfet l=6e-08 w=5.49e-07 $X=32379 $Y=18966 $D=616
M1203 1091 443 1085 vss hvtnfet l=6e-08 w=5.49e-07 $X=32379 $Y=24337 $D=616
M1204 1092 443 1086 vss hvtnfet l=6e-08 w=5.49e-07 $X=32379 $Y=25886 $D=616
M1205 vss aa<7> 449 vss hvtnfet l=6e-08 w=2.74e-07 $X=32394 $Y=13476 $D=616
M1206 vss 324 442 vss hvtnfet l=6e-08 w=5e-07 $X=32394 $Y=32443 $D=616
M1207 b_pxba_n<4> 444 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=32530 $Y=336 $D=616
M1208 444 445 vss vss hvtnfet l=6e-08 w=5e-07 $X=32530 $Y=6701 $D=616
M1209 445 446 vss vss hvtnfet l=6e-08 w=3e-07 $X=32530 $Y=7831 $D=616
M1210 447 446 vss vss hvtnfet l=6e-08 w=3e-07 $X=32530 $Y=43002 $D=616
M1211 448 447 vss vss hvtnfet l=6e-08 w=5e-07 $X=32530 $Y=43932 $D=616
M1212 t_pxba_n<4> 448 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=32530 $Y=49512 $D=616
M1213 vss 442 dwla<1> vss hvtnfet l=6e-08 w=3e-07 $X=32531 $Y=31098 $D=616
M1214 vss 442 497 vss hvtnfet l=6e-08 w=3e-07 $X=32531 $Y=37457 $D=616
M1215 437 dwla<1> 1087 vss hvtnfet l=6e-08 w=4.11e-07 $X=32634 $Y=11276 $D=616
M1216 438 dwla<0> 1088 vss hvtnfet l=6e-08 w=4.11e-07 $X=32634 $Y=39446 $D=616
M1217 428 449 1089 vss hvtnfet l=6e-08 w=5.49e-07 $X=32639 $Y=17417 $D=616
M1218 429 450 1090 vss hvtnfet l=6e-08 w=5.49e-07 $X=32639 $Y=18966 $D=616
M1219 430 449 1091 vss hvtnfet l=6e-08 w=5.49e-07 $X=32639 $Y=24337 $D=616
M1220 431 450 1092 vss hvtnfet l=6e-08 w=5.49e-07 $X=32639 $Y=25886 $D=616
M1221 450 449 vss vss hvtnfet l=6e-08 w=2.74e-07 $X=32654 $Y=13476 $D=616
M1222 vss 444 b_pxba_n<4> vss hvtnfet l=6e-08 w=1.285e-06 $X=32790 $Y=336 $D=616
M1223 vss 445 444 vss hvtnfet l=6e-08 w=5e-07 $X=32790 $Y=6701 $D=616
M1224 vss 446 445 vss hvtnfet l=6e-08 w=3e-07 $X=32790 $Y=7831 $D=616
M1225 vss 446 447 vss hvtnfet l=6e-08 w=3e-07 $X=32790 $Y=43002 $D=616
M1226 vss 447 448 vss hvtnfet l=6e-08 w=5e-07 $X=32790 $Y=43932 $D=616
M1227 vss 448 t_pxba_n<4> vss hvtnfet l=6e-08 w=1.285e-06 $X=32790 $Y=49512 $D=616
M1228 dwla<1> 368 vss vss hvtnfet l=6e-08 w=3e-07 $X=33041 $Y=31098 $D=616
M1229 497 456 vss vss hvtnfet l=6e-08 w=3e-07 $X=33041 $Y=37457 $D=616
M1230 465 442 vss vss hvtnfet l=6e-08 w=4e-07 $X=33094 $Y=32543 $D=616
M1231 1093 dwla<1> 458 vss hvtnfet l=6e-08 w=4.11e-07 $X=33144 $Y=11276 $D=616
M1232 1094 dwla<0> 459 vss hvtnfet l=6e-08 w=4.11e-07 $X=33144 $Y=39446 $D=616
M1233 vss 455 443 vss hvtnfet l=6e-08 w=2.74e-07 $X=33254 $Y=13476 $D=616
M1234 b_pxba_n<3> 451 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=33300 $Y=336 $D=616
M1235 451 452 vss vss hvtnfet l=6e-08 w=5e-07 $X=33300 $Y=6701 $D=616
M1236 452 425 vss vss hvtnfet l=6e-08 w=3e-07 $X=33300 $Y=7831 $D=616
M1237 453 425 vss vss hvtnfet l=6e-08 w=3e-07 $X=33300 $Y=43002 $D=616
M1238 454 453 vss vss hvtnfet l=6e-08 w=5e-07 $X=33300 $Y=43932 $D=616
M1239 t_pxba_n<3> 454 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=33300 $Y=49512 $D=616
M1240 vss 368 dwla<1> vss hvtnfet l=6e-08 w=3e-07 $X=33301 $Y=31098 $D=616
M1241 vss 456 497 vss hvtnfet l=6e-08 w=3e-07 $X=33301 $Y=37457 $D=616
M1242 vss 311 1093 vss hvtnfet l=6e-08 w=4.11e-07 $X=33404 $Y=11276 $D=616
M1243 vss 311 1094 vss hvtnfet l=6e-08 w=4.11e-07 $X=33404 $Y=39446 $D=616
M1244 455 aa<8> vss vss hvtnfet l=6e-08 w=2.74e-07 $X=33514 $Y=13476 $D=616
M1245 vss 451 b_pxba_n<3> vss hvtnfet l=6e-08 w=1.285e-06 $X=33560 $Y=336 $D=616
M1246 vss 452 451 vss hvtnfet l=6e-08 w=5e-07 $X=33560 $Y=6701 $D=616
M1247 vss 425 452 vss hvtnfet l=6e-08 w=3e-07 $X=33560 $Y=7831 $D=616
M1248 vss 425 453 vss hvtnfet l=6e-08 w=3e-07 $X=33560 $Y=43002 $D=616
M1249 vss 453 454 vss hvtnfet l=6e-08 w=5e-07 $X=33560 $Y=43932 $D=616
M1250 vss 454 t_pxba_n<3> vss hvtnfet l=6e-08 w=1.285e-06 $X=33560 $Y=49512 $D=616
M1251 dwla<0> 368 vss vss hvtnfet l=6e-08 w=3e-07 $X=33811 $Y=31098 $D=616
M1252 498 456 vss vss hvtnfet l=6e-08 w=3e-07 $X=33811 $Y=37457 $D=616
M1253 555 458 vss vss hvtnfet l=6e-08 w=2e-07 $X=33914 $Y=11276 $D=616
M1254 559 459 vss vss hvtnfet l=6e-08 w=2e-07 $X=33914 $Y=39657 $D=616
M1255 b_pxba_n<2> 460 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=34070 $Y=336 $D=616
M1256 460 461 vss vss hvtnfet l=6e-08 w=5e-07 $X=34070 $Y=6701 $D=616
M1257 461 424 vss vss hvtnfet l=6e-08 w=3e-07 $X=34070 $Y=7831 $D=616
M1258 462 424 vss vss hvtnfet l=6e-08 w=3e-07 $X=34070 $Y=43002 $D=616
M1259 463 462 vss vss hvtnfet l=6e-08 w=5e-07 $X=34070 $Y=43932 $D=616
M1260 t_pxba_n<2> 463 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=34070 $Y=49512 $D=616
M1261 vss 368 dwla<0> vss hvtnfet l=6e-08 w=3e-07 $X=34071 $Y=31098 $D=616
M1262 vss 456 498 vss hvtnfet l=6e-08 w=3e-07 $X=34071 $Y=37457 $D=616
M1263 vss 460 b_pxba_n<2> vss hvtnfet l=6e-08 w=1.285e-06 $X=34330 $Y=336 $D=616
M1264 vss 461 460 vss hvtnfet l=6e-08 w=5e-07 $X=34330 $Y=6701 $D=616
M1265 vss 424 461 vss hvtnfet l=6e-08 w=3e-07 $X=34330 $Y=7831 $D=616
M1266 vss 424 462 vss hvtnfet l=6e-08 w=3e-07 $X=34330 $Y=43002 $D=616
M1267 vss 462 463 vss hvtnfet l=6e-08 w=5e-07 $X=34330 $Y=43932 $D=616
M1268 vss 463 t_pxba_n<2> vss hvtnfet l=6e-08 w=1.285e-06 $X=34330 $Y=49512 $D=616
M1269 1095 449 479 vss hvtnfet l=6e-08 w=5.49e-07 $X=34479 $Y=17417 $D=616
M1270 1096 450 480 vss hvtnfet l=6e-08 w=5.49e-07 $X=34479 $Y=18966 $D=616
M1271 1097 449 481 vss hvtnfet l=6e-08 w=5.49e-07 $X=34479 $Y=24337 $D=616
M1272 1098 450 482 vss hvtnfet l=6e-08 w=5.49e-07 $X=34479 $Y=25886 $D=616
M1273 vss aa<9> 440 vss hvtnfet l=6e-08 w=2.74e-07 $X=34524 $Y=13476 $D=616
M1274 dwla<0> 465 vss vss hvtnfet l=6e-08 w=3e-07 $X=34581 $Y=31098 $D=616
M1275 498 465 vss vss hvtnfet l=6e-08 w=3e-07 $X=34581 $Y=37457 $D=616
M1276 1099 vdd vss vss hvtnfet l=6e-08 w=6.4e-07 $X=34621 $Y=32508 $D=616
M1277 123 131 vss vss hvtnfet l=6e-08 w=2e-07 $X=34646 $Y=11546 $D=616
M1278 1100 455 1095 vss hvtnfet l=6e-08 w=5.49e-07 $X=34739 $Y=17417 $D=616
M1279 1101 455 1096 vss hvtnfet l=6e-08 w=5.49e-07 $X=34739 $Y=18966 $D=616
M1280 1102 455 1097 vss hvtnfet l=6e-08 w=5.49e-07 $X=34739 $Y=24337 $D=616
M1281 1103 455 1098 vss hvtnfet l=6e-08 w=5.49e-07 $X=34739 $Y=25886 $D=616
M1282 b_pxba_n<1> 466 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=34840 $Y=336 $D=616
M1283 466 467 vss vss hvtnfet l=6e-08 w=5e-07 $X=34840 $Y=6701 $D=616
M1284 467 468 vss vss hvtnfet l=6e-08 w=3e-07 $X=34840 $Y=7831 $D=616
M1285 469 468 vss vss hvtnfet l=6e-08 w=3e-07 $X=34840 $Y=43002 $D=616
M1286 470 469 vss vss hvtnfet l=6e-08 w=5e-07 $X=34840 $Y=43932 $D=616
M1287 t_pxba_n<1> 470 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=34840 $Y=49512 $D=616
M1288 vss 465 dwla<0> vss hvtnfet l=6e-08 w=3e-07 $X=34841 $Y=31098 $D=616
M1289 vss 465 498 vss hvtnfet l=6e-08 w=3e-07 $X=34841 $Y=37457 $D=616
M1290 535 471 1099 vss hvtnfet l=6e-08 w=6.4e-07 $X=34881 $Y=32508 $D=616
M1291 vss 123 123 vss hvtnfet l=6e-08 w=2e-07 $X=34906 $Y=11546 $D=616
M1292 1104 439 1100 vss hvtnfet l=6e-08 w=5.49e-07 $X=34999 $Y=17417 $D=616
M1293 1105 439 1101 vss hvtnfet l=6e-08 w=5.49e-07 $X=34999 $Y=18966 $D=616
M1294 1106 440 1102 vss hvtnfet l=6e-08 w=5.49e-07 $X=34999 $Y=24337 $D=616
M1295 1107 440 1103 vss hvtnfet l=6e-08 w=5.49e-07 $X=34999 $Y=25886 $D=616
M1296 439 440 vss vss hvtnfet l=6e-08 w=2.74e-07 $X=35034 $Y=13476 $D=616
M1297 vss 466 b_pxba_n<1> vss hvtnfet l=6e-08 w=1.285e-06 $X=35100 $Y=336 $D=616
M1298 vss 467 466 vss hvtnfet l=6e-08 w=5e-07 $X=35100 $Y=6701 $D=616
M1299 vss 468 467 vss hvtnfet l=6e-08 w=3e-07 $X=35100 $Y=7831 $D=616
M1300 vss 468 469 vss hvtnfet l=6e-08 w=3e-07 $X=35100 $Y=43002 $D=616
M1301 vss 469 470 vss hvtnfet l=6e-08 w=5e-07 $X=35100 $Y=43932 $D=616
M1302 vss 470 t_pxba_n<1> vss hvtnfet l=6e-08 w=1.285e-06 $X=35100 $Y=49512 $D=616
M1303 vss 323 1104 vss hvtnfet l=6e-08 w=8.23e-07 $X=35269 $Y=17143 $D=616
M1304 vss 323 1105 vss hvtnfet l=6e-08 w=8.23e-07 $X=35269 $Y=18966 $D=616
M1305 vss 323 1106 vss hvtnfet l=6e-08 w=8.23e-07 $X=35269 $Y=24063 $D=616
M1306 vss 323 1107 vss hvtnfet l=6e-08 w=8.23e-07 $X=35269 $Y=25886 $D=616
M1307 vss 473 484 vss hvtnfet l=6e-08 w=3e-07 $X=35351 $Y=37257 $D=616
M1308 vss 472 471 vss hvtnfet l=6e-08 w=3.5e-07 $X=35446 $Y=32613 $D=616
M1309 b_pxba_n<0> 474 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=35610 $Y=336 $D=616
M1310 474 475 vss vss hvtnfet l=6e-08 w=5e-07 $X=35610 $Y=6701 $D=616
M1311 475 476 vss vss hvtnfet l=6e-08 w=3e-07 $X=35610 $Y=7831 $D=616
M1312 477 476 vss vss hvtnfet l=6e-08 w=3e-07 $X=35610 $Y=43002 $D=616
M1313 478 477 vss vss hvtnfet l=6e-08 w=5e-07 $X=35610 $Y=43932 $D=616
M1314 t_pxba_n<0> 478 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=35610 $Y=49512 $D=616
M1315 472 483 vss vss hvtnfet l=2.5e-07 w=3.5e-07 $X=35706 $Y=32613 $D=616
M1316 446 479 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=35764 $Y=17812 $D=616
M1317 434 480 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=35764 $Y=18983 $D=616
M1318 476 481 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=35764 $Y=24732 $D=616
M1319 468 482 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=35764 $Y=25903 $D=616
M1320 1108 317 479 vss hvtnfet l=6e-08 w=1.8e-07 $X=35779 $Y=17143 $D=616
M1321 1109 317 480 vss hvtnfet l=6e-08 w=1.8e-07 $X=35779 $Y=19609 $D=616
M1322 1110 317 481 vss hvtnfet l=6e-08 w=1.8e-07 $X=35779 $Y=24063 $D=616
M1323 1111 317 482 vss hvtnfet l=6e-08 w=1.8e-07 $X=35779 $Y=26529 $D=616
M1324 473 484 vss vss hvtnfet l=1.2e-07 w=1.5e-07 $X=35861 $Y=37297 $D=616
M1325 vss 474 b_pxba_n<0> vss hvtnfet l=6e-08 w=1.285e-06 $X=35870 $Y=336 $D=616
M1326 vss 475 474 vss hvtnfet l=6e-08 w=5e-07 $X=35870 $Y=6701 $D=616
M1327 vss 476 475 vss hvtnfet l=6e-08 w=3e-07 $X=35870 $Y=7831 $D=616
M1328 vss 476 477 vss hvtnfet l=6e-08 w=3e-07 $X=35870 $Y=43002 $D=616
M1329 vss 477 478 vss hvtnfet l=6e-08 w=5e-07 $X=35870 $Y=43932 $D=616
M1330 vss 478 t_pxba_n<0> vss hvtnfet l=6e-08 w=1.285e-06 $X=35870 $Y=49512 $D=616
M1331 773 495 vss vss hvtnfet l=6e-08 w=8e-07 $X=35945 $Y=30668 $D=616
M1332 vss 479 446 vss hvtnfet l=6e-08 w=1.37e-07 $X=36024 $Y=17812 $D=616
M1333 vss 480 434 vss hvtnfet l=6e-08 w=1.37e-07 $X=36024 $Y=18983 $D=616
M1334 vss 481 476 vss hvtnfet l=6e-08 w=1.37e-07 $X=36024 $Y=24732 $D=616
M1335 vss 482 468 vss hvtnfet l=6e-08 w=1.37e-07 $X=36024 $Y=25903 $D=616
M1336 vss 446 1108 vss hvtnfet l=6e-08 w=1.8e-07 $X=36039 $Y=17143 $D=616
M1337 vss 434 1109 vss hvtnfet l=6e-08 w=1.8e-07 $X=36039 $Y=19609 $D=616
M1338 vss 476 1110 vss hvtnfet l=6e-08 w=1.8e-07 $X=36039 $Y=24063 $D=616
M1339 vss 468 1111 vss hvtnfet l=6e-08 w=1.8e-07 $X=36039 $Y=26529 $D=616
M1340 vss 495 773 vss hvtnfet l=6e-08 w=8e-07 $X=36205 $Y=30668 $D=616
M1341 vss 491 509 vss hvtnfet l=6e-08 w=2.74e-07 $X=36254 $Y=13476 $D=616
M1342 b_pxaa<3> 485 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=36380 $Y=336 $D=616
M1343 485 486 vss vss hvtnfet l=6e-08 w=5e-07 $X=36380 $Y=6701 $D=616
M1344 486 487 vss vss hvtnfet l=6e-08 w=3e-07 $X=36380 $Y=7831 $D=616
M1345 1112 492 vss vss hvtnfet l=6e-08 w=4.11e-07 $X=36380 $Y=11276 $D=616
M1346 1113 492 vss vss hvtnfet l=6e-08 w=4.11e-07 $X=36380 $Y=39446 $D=616
M1347 489 488 vss vss hvtnfet l=6e-08 w=3e-07 $X=36380 $Y=43002 $D=616
M1348 490 489 vss vss hvtnfet l=6e-08 w=5e-07 $X=36380 $Y=43932 $D=616
M1349 t_pxaa<3> 490 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=36380 $Y=49512 $D=616
M1350 vss 494 473 vss hvtnfet l=6e-08 w=3.2e-07 $X=36431 $Y=37292 $D=616
M1351 vss 496 483 vss hvtnfet l=6e-08 w=3.2e-07 $X=36466 $Y=32828 $D=616
M1352 vss 485 b_pxaa<3> vss hvtnfet l=6e-08 w=1.285e-06 $X=36640 $Y=336 $D=616
M1353 vss 486 485 vss hvtnfet l=6e-08 w=5e-07 $X=36640 $Y=6701 $D=616
M1354 vss 487 486 vss hvtnfet l=6e-08 w=3e-07 $X=36640 $Y=7831 $D=616
M1355 487 497 1112 vss hvtnfet l=6e-08 w=4.11e-07 $X=36640 $Y=11276 $D=616
M1356 488 498 1113 vss hvtnfet l=6e-08 w=4.11e-07 $X=36640 $Y=39446 $D=616
M1357 vss 488 489 vss hvtnfet l=6e-08 w=3e-07 $X=36640 $Y=43002 $D=616
M1358 vss 489 490 vss hvtnfet l=6e-08 w=5e-07 $X=36640 $Y=43932 $D=616
M1359 vss 490 t_pxaa<3> vss hvtnfet l=6e-08 w=1.285e-06 $X=36640 $Y=49512 $D=616
M1360 368 clka 773 vss hvtnfet l=6e-08 w=8e-07 $X=36715 $Y=30668 $D=616
M1361 491 aa<6> vss vss hvtnfet l=6e-08 w=2.74e-07 $X=36764 $Y=13476 $D=616
M1362 773 clka 368 vss hvtnfet l=6e-08 w=8e-07 $X=36975 $Y=30668 $D=616
M1363 vss 473 496 vss hvtnfet l=6e-08 w=3.2e-07 $X=36976 $Y=32828 $D=616
M1364 1114 501 519 vss hvtnfet l=6e-08 w=5.49e-07 $X=37059 $Y=17143 $D=616
M1365 1115 502 520 vss hvtnfet l=6e-08 w=5.49e-07 $X=37059 $Y=19240 $D=616
M1366 1116 501 521 vss hvtnfet l=6e-08 w=5.49e-07 $X=37059 $Y=24063 $D=616
M1367 1117 502 522 vss hvtnfet l=6e-08 w=5.49e-07 $X=37059 $Y=26160 $D=616
M1368 b_pxaa<2> 503 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=37150 $Y=336 $D=616
M1369 503 504 vss vss hvtnfet l=6e-08 w=5e-07 $X=37150 $Y=6701 $D=616
M1370 504 505 vss vss hvtnfet l=6e-08 w=3e-07 $X=37150 $Y=7831 $D=616
M1371 1118 497 505 vss hvtnfet l=6e-08 w=4.11e-07 $X=37150 $Y=11276 $D=616
M1372 1119 498 506 vss hvtnfet l=6e-08 w=4.11e-07 $X=37150 $Y=39446 $D=616
M1373 507 506 vss vss hvtnfet l=6e-08 w=3e-07 $X=37150 $Y=43002 $D=616
M1374 508 507 vss vss hvtnfet l=6e-08 w=5e-07 $X=37150 $Y=43932 $D=616
M1375 t_pxaa<2> 508 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=37150 $Y=49512 $D=616
M1376 vss ddqa_n 493 vss hvtnfet l=6e-08 w=2.4e-07 $X=37161 $Y=37292 $D=616
M1377 vss 502 501 vss hvtnfet l=6e-08 w=2.74e-07 $X=37274 $Y=13476 $D=616
M1378 1120 509 1114 vss hvtnfet l=6e-08 w=5.49e-07 $X=37319 $Y=17143 $D=616
M1379 1121 509 1115 vss hvtnfet l=6e-08 w=5.49e-07 $X=37319 $Y=19240 $D=616
M1380 1122 491 1116 vss hvtnfet l=6e-08 w=5.49e-07 $X=37319 $Y=24063 $D=616
M1381 1123 491 1117 vss hvtnfet l=6e-08 w=5.49e-07 $X=37319 $Y=26160 $D=616
M1382 vss 503 b_pxaa<2> vss hvtnfet l=6e-08 w=1.285e-06 $X=37410 $Y=336 $D=616
M1383 vss 504 503 vss hvtnfet l=6e-08 w=5e-07 $X=37410 $Y=6701 $D=616
M1384 vss 505 504 vss hvtnfet l=6e-08 w=3e-07 $X=37410 $Y=7831 $D=616
M1385 vss 510 1118 vss hvtnfet l=6e-08 w=4.11e-07 $X=37410 $Y=11276 $D=616
M1386 vss 510 1119 vss hvtnfet l=6e-08 w=4.11e-07 $X=37410 $Y=39446 $D=616
M1387 vss 506 507 vss hvtnfet l=6e-08 w=3e-07 $X=37410 $Y=43002 $D=616
M1388 vss 507 508 vss hvtnfet l=6e-08 w=5e-07 $X=37410 $Y=43932 $D=616
M1389 vss 508 t_pxaa<2> vss hvtnfet l=6e-08 w=1.285e-06 $X=37410 $Y=49512 $D=616
M1390 493 ddqa vss vss hvtnfet l=6e-08 w=2.4e-07 $X=37421 $Y=37292 $D=616
M1391 vss clka 524 vss hvtnfet l=6e-08 w=6e-07 $X=37485 $Y=30668 $D=616
M1392 vss 323 1120 vss hvtnfet l=6e-08 w=8.23e-07 $X=37589 $Y=17143 $D=616
M1393 vss 323 1121 vss hvtnfet l=6e-08 w=8.23e-07 $X=37589 $Y=18966 $D=616
M1394 vss 323 1122 vss hvtnfet l=6e-08 w=8.23e-07 $X=37589 $Y=24063 $D=616
M1395 vss 323 1123 vss hvtnfet l=6e-08 w=8.23e-07 $X=37589 $Y=25886 $D=616
M1396 1124 496 557 vss hvtnfet l=6e-08 w=6.4e-07 $X=37661 $Y=32508 $D=616
M1397 502 aa<5> vss vss hvtnfet l=6e-08 w=2.74e-07 $X=37784 $Y=13476 $D=616
M1398 b_pxaa<1> 512 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=37920 $Y=336 $D=616
M1399 512 513 vss vss hvtnfet l=6e-08 w=5e-07 $X=37920 $Y=6701 $D=616
M1400 513 514 vss vss hvtnfet l=6e-08 w=3e-07 $X=37920 $Y=7831 $D=616
M1401 1125 523 vss vss hvtnfet l=6e-08 w=4.11e-07 $X=37920 $Y=11276 $D=616
M1402 1126 523 vss vss hvtnfet l=6e-08 w=4.11e-07 $X=37920 $Y=39446 $D=616
M1403 516 515 vss vss hvtnfet l=6e-08 w=3e-07 $X=37920 $Y=43002 $D=616
M1404 517 516 vss vss hvtnfet l=6e-08 w=5e-07 $X=37920 $Y=43932 $D=616
M1405 t_pxaa<1> 517 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=37920 $Y=49512 $D=616
M1406 vss 386 1124 vss hvtnfet l=6e-08 w=6.4e-07 $X=37921 $Y=32508 $D=616
M1407 1127 317 519 vss hvtnfet l=6e-08 w=1.8e-07 $X=38099 $Y=17143 $D=616
M1408 492 519 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=38099 $Y=17812 $D=616
M1409 510 520 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=38099 $Y=18983 $D=616
M1410 1128 317 520 vss hvtnfet l=6e-08 w=1.8e-07 $X=38099 $Y=19609 $D=616
M1411 1129 317 521 vss hvtnfet l=6e-08 w=1.8e-07 $X=38099 $Y=24063 $D=616
M1412 523 521 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=38099 $Y=24732 $D=616
M1413 525 522 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=38099 $Y=25903 $D=616
M1414 1130 317 522 vss hvtnfet l=6e-08 w=1.8e-07 $X=38099 $Y=26529 $D=616
M1415 vss 493 526 vss hvtnfet l=1.4e-07 w=3.2e-07 $X=38141 $Y=37127 $D=616
M1416 vss 512 b_pxaa<1> vss hvtnfet l=6e-08 w=1.285e-06 $X=38180 $Y=336 $D=616
M1417 vss 513 512 vss hvtnfet l=6e-08 w=5e-07 $X=38180 $Y=6701 $D=616
M1418 vss 514 513 vss hvtnfet l=6e-08 w=3e-07 $X=38180 $Y=7831 $D=616
M1419 514 497 1125 vss hvtnfet l=6e-08 w=4.11e-07 $X=38180 $Y=11276 $D=616
M1420 515 498 1126 vss hvtnfet l=6e-08 w=4.11e-07 $X=38180 $Y=39446 $D=616
M1421 vss 515 516 vss hvtnfet l=6e-08 w=3e-07 $X=38180 $Y=43002 $D=616
M1422 vss 516 517 vss hvtnfet l=6e-08 w=5e-07 $X=38180 $Y=43932 $D=616
M1423 vss 517 t_pxaa<1> vss hvtnfet l=6e-08 w=1.285e-06 $X=38180 $Y=49512 $D=616
M1424 vss 524 534 vss hvtnfet l=6e-08 w=5.49e-07 $X=38255 $Y=30668 $D=616
M1425 vss 492 1127 vss hvtnfet l=6e-08 w=1.8e-07 $X=38359 $Y=17143 $D=616
M1426 vss 519 492 vss hvtnfet l=6e-08 w=1.37e-07 $X=38359 $Y=17812 $D=616
M1427 vss 520 510 vss hvtnfet l=6e-08 w=1.37e-07 $X=38359 $Y=18983 $D=616
M1428 vss 510 1128 vss hvtnfet l=6e-08 w=1.8e-07 $X=38359 $Y=19609 $D=616
M1429 vss 523 1129 vss hvtnfet l=6e-08 w=1.8e-07 $X=38359 $Y=24063 $D=616
M1430 vss 521 523 vss hvtnfet l=6e-08 w=1.37e-07 $X=38359 $Y=24732 $D=616
M1431 vss 522 525 vss hvtnfet l=6e-08 w=1.37e-07 $X=38359 $Y=25903 $D=616
M1432 vss 525 1130 vss hvtnfet l=6e-08 w=1.8e-07 $X=38359 $Y=26529 $D=616
M1433 779 494 vss vss hvtnfet l=6e-08 w=3.2e-07 $X=38431 $Y=32828 $D=616
M1434 780 526 vss vss hvtnfet l=1.4e-07 w=3.2e-07 $X=38481 $Y=37127 $D=616
M1435 534 495 vss vss hvtnfet l=6e-08 w=5.49e-07 $X=38515 $Y=30668 $D=616
M1436 vss 533 546 vss hvtnfet l=6e-08 w=2.74e-07 $X=38574 $Y=13476 $D=616
M1437 b_pxaa<0> 527 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=38690 $Y=336 $D=616
M1438 527 528 vss vss hvtnfet l=6e-08 w=5e-07 $X=38690 $Y=6701 $D=616
M1439 528 529 vss vss hvtnfet l=6e-08 w=3e-07 $X=38690 $Y=7831 $D=616
M1440 1131 497 529 vss hvtnfet l=6e-08 w=4.11e-07 $X=38690 $Y=11276 $D=616
M1441 1132 498 530 vss hvtnfet l=6e-08 w=4.11e-07 $X=38690 $Y=39446 $D=616
M1442 531 530 vss vss hvtnfet l=6e-08 w=3e-07 $X=38690 $Y=43002 $D=616
M1443 532 531 vss vss hvtnfet l=6e-08 w=5e-07 $X=38690 $Y=43932 $D=616
M1444 t_pxaa<0> 532 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=38690 $Y=49512 $D=616
M1445 vss 527 b_pxaa<0> vss hvtnfet l=6e-08 w=1.285e-06 $X=38950 $Y=336 $D=616
M1446 vss 528 527 vss hvtnfet l=6e-08 w=5e-07 $X=38950 $Y=6701 $D=616
M1447 vss 529 528 vss hvtnfet l=6e-08 w=3e-07 $X=38950 $Y=7831 $D=616
M1448 vss 525 1131 vss hvtnfet l=6e-08 w=4.11e-07 $X=38950 $Y=11276 $D=616
M1449 vss 525 1132 vss hvtnfet l=6e-08 w=4.11e-07 $X=38950 $Y=39446 $D=616
M1450 vss 530 531 vss hvtnfet l=6e-08 w=3e-07 $X=38950 $Y=43002 $D=616
M1451 vss 531 532 vss hvtnfet l=6e-08 w=5e-07 $X=38950 $Y=43932 $D=616
M1452 vss 532 t_pxaa<0> vss hvtnfet l=6e-08 w=1.285e-06 $X=38950 $Y=49512 $D=616
M1453 vss 534 495 vss hvtnfet l=6e-08 w=5.49e-07 $X=39025 $Y=30668 $D=616
M1454 533 aa<3> vss vss hvtnfet l=6e-08 w=2.74e-07 $X=39084 $Y=13476 $D=616
M1455 vss clka 323 vss hvtnfet l=6e-08 w=6e-07 $X=39174 $Y=32403 $D=616
M1456 293 535 vss vss hvtnfet l=6e-08 w=6e-07 $X=39185 $Y=37277 $D=616
M1457 495 539 vss vss hvtnfet l=6e-08 w=5.49e-07 $X=39285 $Y=30668 $D=616
M1458 1133 537 549 vss hvtnfet l=6e-08 w=5.49e-07 $X=39379 $Y=17143 $D=616
M1459 1134 538 550 vss hvtnfet l=6e-08 w=5.49e-07 $X=39379 $Y=19240 $D=616
M1460 1135 537 551 vss hvtnfet l=6e-08 w=5.49e-07 $X=39379 $Y=24063 $D=616
M1461 1136 538 552 vss hvtnfet l=6e-08 w=5.49e-07 $X=39379 $Y=26160 $D=616
M1462 323 clka vss vss hvtnfet l=6e-08 w=6e-07 $X=39434 $Y=32403 $D=616
M1463 vss 538 537 vss hvtnfet l=6e-08 w=2.74e-07 $X=39594 $Y=13476 $D=616
M1464 1137 546 1133 vss hvtnfet l=6e-08 w=5.49e-07 $X=39639 $Y=17143 $D=616
M1465 1138 546 1134 vss hvtnfet l=6e-08 w=5.49e-07 $X=39639 $Y=19240 $D=616
M1466 1139 533 1135 vss hvtnfet l=6e-08 w=5.49e-07 $X=39639 $Y=24063 $D=616
M1467 1140 533 1136 vss hvtnfet l=6e-08 w=5.49e-07 $X=39639 $Y=26160 $D=616
M1468 r_sa_prea_n 293 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=39695 $Y=37027 $D=616
M1469 289 540 vss vss hvtnfet l=6e-08 w=6e-07 $X=39705 $Y=336 $D=616
M1470 290 541 vss vss hvtnfet l=6e-08 w=6e-07 $X=39705 $Y=5566 $D=616
M1471 291 542 vss vss hvtnfet l=6e-08 w=6e-07 $X=39705 $Y=6796 $D=616
M1472 292 543 vss vss hvtnfet l=6e-08 w=6e-07 $X=39705 $Y=12026 $D=616
M1473 294 543 vss vss hvtnfet l=6e-08 w=6e-07 $X=39705 $Y=38507 $D=616
M1474 295 542 vss vss hvtnfet l=6e-08 w=6e-07 $X=39705 $Y=43737 $D=616
M1475 296 544 vss vss hvtnfet l=6e-08 w=6e-07 $X=39705 $Y=44967 $D=616
M1476 297 545 vss vss hvtnfet l=6e-08 w=6e-07 $X=39705 $Y=50197 $D=616
M1477 vss stclka 539 vss hvtnfet l=6e-08 w=2.74e-07 $X=39795 $Y=30668 $D=616
M1478 vss 323 1137 vss hvtnfet l=6e-08 w=8.23e-07 $X=39909 $Y=17143 $D=616
M1479 vss 323 1138 vss hvtnfet l=6e-08 w=8.23e-07 $X=39909 $Y=18966 $D=616
M1480 vss 323 1139 vss hvtnfet l=6e-08 w=8.23e-07 $X=39909 $Y=24063 $D=616
M1481 vss 323 1140 vss hvtnfet l=6e-08 w=8.23e-07 $X=39909 $Y=25886 $D=616
M1482 vss 293 r_sa_prea_n vss hvtnfet l=6e-08 w=8.58e-07 $X=39955 $Y=37027 $D=616
M1483 538 aa<2> vss vss hvtnfet l=6e-08 w=2.74e-07 $X=40104 $Y=13476 $D=616
M1484 rb_ca<1> 289 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=40215 $Y=328 $D=616
M1485 rb_ca<3> 290 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=40215 $Y=5316 $D=616
M1486 rb_ma<1> 291 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=40215 $Y=6788 $D=616
M1487 rb_ma<3> 292 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=40215 $Y=11776 $D=616
M1488 r_sa_prea_n 293 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=40215 $Y=37027 $D=616
M1489 rt_ma<3> 294 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=40215 $Y=38499 $D=616
M1490 rt_ma<1> 295 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=40215 $Y=43487 $D=616
M1491 rt_ca<3> 296 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=40215 $Y=44959 $D=616
M1492 rt_ca<1> 297 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=40215 $Y=49947 $D=616
M1493 1141 317 549 vss hvtnfet l=6e-08 w=1.8e-07 $X=40419 $Y=17143 $D=616
M1494 543 549 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=40419 $Y=17812 $D=616
M1495 553 550 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=40419 $Y=18983 $D=616
M1496 1142 317 550 vss hvtnfet l=6e-08 w=1.8e-07 $X=40419 $Y=19609 $D=616
M1497 1143 317 551 vss hvtnfet l=6e-08 w=1.8e-07 $X=40419 $Y=24063 $D=616
M1498 542 551 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=40419 $Y=24732 $D=616
M1499 554 552 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=40419 $Y=25903 $D=616
M1500 1144 317 552 vss hvtnfet l=6e-08 w=1.8e-07 $X=40419 $Y=26529 $D=616
M1501 vss 289 rb_ca<1> vss hvtnfet l=6e-08 w=8.58e-07 $X=40475 $Y=328 $D=616
M1502 vss 290 rb_ca<3> vss hvtnfet l=6e-08 w=8.58e-07 $X=40475 $Y=5316 $D=616
M1503 vss 291 rb_ma<1> vss hvtnfet l=6e-08 w=8.58e-07 $X=40475 $Y=6788 $D=616
M1504 vss 292 rb_ma<3> vss hvtnfet l=6e-08 w=8.58e-07 $X=40475 $Y=11776 $D=616
M1505 vss 294 rt_ma<3> vss hvtnfet l=6e-08 w=8.58e-07 $X=40475 $Y=38499 $D=616
M1506 vss 295 rt_ma<1> vss hvtnfet l=6e-08 w=8.58e-07 $X=40475 $Y=43487 $D=616
M1507 vss 296 rt_ca<3> vss hvtnfet l=6e-08 w=8.58e-07 $X=40475 $Y=44959 $D=616
M1508 vss 297 rt_ca<1> vss hvtnfet l=6e-08 w=8.58e-07 $X=40475 $Y=49947 $D=616
M1509 vss 543 1141 vss hvtnfet l=6e-08 w=1.8e-07 $X=40679 $Y=17143 $D=616
M1510 vss 549 543 vss hvtnfet l=6e-08 w=1.37e-07 $X=40679 $Y=17812 $D=616
M1511 vss 550 553 vss hvtnfet l=6e-08 w=1.37e-07 $X=40679 $Y=18983 $D=616
M1512 vss 553 1142 vss hvtnfet l=6e-08 w=1.8e-07 $X=40679 $Y=19609 $D=616
M1513 vss 542 1143 vss hvtnfet l=6e-08 w=1.8e-07 $X=40679 $Y=24063 $D=616
M1514 vss 551 542 vss hvtnfet l=6e-08 w=1.37e-07 $X=40679 $Y=24732 $D=616
M1515 vss 552 554 vss hvtnfet l=6e-08 w=1.37e-07 $X=40679 $Y=25903 $D=616
M1516 vss 554 1144 vss hvtnfet l=6e-08 w=1.8e-07 $X=40679 $Y=26529 $D=616
M1517 vss 303 r_saea_n vss hvtnfet l=6e-08 w=8.58e-07 $X=40725 $Y=37027 $D=616
M1518 rb_ca<1> 289 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=40735 $Y=328 $D=616
M1519 rb_ca<3> 290 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=40735 $Y=5316 $D=616
M1520 rb_ma<1> 291 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=40735 $Y=6788 $D=616
M1521 rb_ma<3> 292 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=40735 $Y=11776 $D=616
M1522 rt_ma<3> 294 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=40735 $Y=38499 $D=616
M1523 rt_ma<1> 295 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=40735 $Y=43487 $D=616
M1524 rt_ca<3> 296 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=40735 $Y=44959 $D=616
M1525 rt_ca<1> 297 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=40735 $Y=49947 $D=616
M1526 r_saea_n 303 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=40985 $Y=37027 $D=616
M1527 vss 299 rb_ca<0> vss hvtnfet l=6e-08 w=8.58e-07 $X=41245 $Y=328 $D=616
M1528 vss 300 rb_ca<2> vss hvtnfet l=6e-08 w=8.58e-07 $X=41245 $Y=5316 $D=616
M1529 vss 301 rb_ma<0> vss hvtnfet l=6e-08 w=8.58e-07 $X=41245 $Y=6788 $D=616
M1530 vss 302 rb_ma<2> vss hvtnfet l=6e-08 w=8.58e-07 $X=41245 $Y=11776 $D=616
M1531 vss 303 r_saea_n vss hvtnfet l=6e-08 w=8.58e-07 $X=41245 $Y=37027 $D=616
M1532 vss 304 rt_ma<2> vss hvtnfet l=6e-08 w=8.58e-07 $X=41245 $Y=38499 $D=616
M1533 vss 305 rt_ma<0> vss hvtnfet l=6e-08 w=8.58e-07 $X=41245 $Y=43487 $D=616
M1534 vss 306 rt_ca<2> vss hvtnfet l=6e-08 w=8.58e-07 $X=41245 $Y=44959 $D=616
M1535 vss 307 rt_ca<0> vss hvtnfet l=6e-08 w=8.58e-07 $X=41245 $Y=49947 $D=616
M1536 vss clka 287 vss hvtnfet l=6e-08 w=1.05e-06 $X=41495 $Y=22251 $D=616
M1537 vss 340 288 vss hvtnfet l=6e-08 w=1.05e-06 $X=41495 $Y=29007 $D=616
M1538 rb_ca<0> 299 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=41505 $Y=328 $D=616
M1539 rb_ca<2> 300 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=41505 $Y=5316 $D=616
M1540 rb_ma<0> 301 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=41505 $Y=6788 $D=616
M1541 rb_ma<2> 302 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=41505 $Y=11776 $D=616
M1542 285 497 vss vss hvtnfet l=6e-08 w=6e-07 $X=41505 $Y=13282 $D=616
M1543 286 498 vss vss hvtnfet l=6e-08 w=6e-07 $X=41505 $Y=20809 $D=616
M1544 r_saea_n 303 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=41505 $Y=37027 $D=616
M1545 rt_ma<2> 304 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=41505 $Y=38499 $D=616
M1546 rt_ma<0> 305 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=41505 $Y=43487 $D=616
M1547 rt_ca<2> 306 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=41505 $Y=44959 $D=616
M1548 rt_ca<0> 307 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=41505 $Y=49947 $D=616
M1549 r_clk_dqa 287 vss vss hvtnfet l=6e-08 w=1.26e-06 $X=41755 $Y=22041 $D=616
M1550 r_clk_dqa_n 288 vss vss hvtnfet l=6e-08 w=1.26e-06 $X=41755 $Y=29007 $D=616
M1551 vss 299 rb_ca<0> vss hvtnfet l=6e-08 w=8.58e-07 $X=41765 $Y=328 $D=616
M1552 vss 300 rb_ca<2> vss hvtnfet l=6e-08 w=8.58e-07 $X=41765 $Y=5316 $D=616
M1553 vss 301 rb_ma<0> vss hvtnfet l=6e-08 w=8.58e-07 $X=41765 $Y=6788 $D=616
M1554 vss 302 rb_ma<2> vss hvtnfet l=6e-08 w=8.58e-07 $X=41765 $Y=11776 $D=616
M1555 vss 303 r_saea_n vss hvtnfet l=6e-08 w=8.58e-07 $X=41765 $Y=37027 $D=616
M1556 vss 304 rt_ma<2> vss hvtnfet l=6e-08 w=8.58e-07 $X=41765 $Y=38499 $D=616
M1557 vss 305 rt_ma<0> vss hvtnfet l=6e-08 w=8.58e-07 $X=41765 $Y=43487 $D=616
M1558 vss 306 rt_ca<2> vss hvtnfet l=6e-08 w=8.58e-07 $X=41765 $Y=44959 $D=616
M1559 vss 307 rt_ca<0> vss hvtnfet l=6e-08 w=8.58e-07 $X=41765 $Y=49947 $D=616
M1560 rb_tm_prea_n 285 vss vss hvtnfet l=6e-08 w=1.287e-06 $X=42015 $Y=13280 $D=616
M1561 rt_tm_prea_n 286 vss vss hvtnfet l=6e-08 w=1.287e-06 $X=42015 $Y=20124 $D=616
M1562 vss 287 r_clk_dqa vss hvtnfet l=6e-08 w=1.26e-06 $X=42015 $Y=22041 $D=616
M1563 vss 288 r_clk_dqa_n vss hvtnfet l=6e-08 w=1.26e-06 $X=42015 $Y=29007 $D=616
M1564 r_lwea 284 vss vss hvtnfet l=6e-08 w=1.287e-06 $X=42015 $Y=30897 $D=616
M1565 vss 555 299 vss hvtnfet l=6e-08 w=6e-07 $X=42275 $Y=336 $D=616
M1566 vss 556 300 vss hvtnfet l=6e-08 w=6e-07 $X=42275 $Y=5566 $D=616
M1567 vss 554 301 vss hvtnfet l=6e-08 w=6e-07 $X=42275 $Y=6796 $D=616
M1568 vss 553 302 vss hvtnfet l=6e-08 w=6e-07 $X=42275 $Y=12026 $D=616
M1569 vss 285 rb_tm_prea_n vss hvtnfet l=6e-08 w=1.287e-06 $X=42275 $Y=13280 $D=616
M1570 vss 286 rt_tm_prea_n vss hvtnfet l=6e-08 w=1.287e-06 $X=42275 $Y=20124 $D=616
M1571 r_clk_dqa 287 vss vss hvtnfet l=6e-08 w=1.26e-06 $X=42275 $Y=22041 $D=616
M1572 r_clk_dqa_n 288 vss vss hvtnfet l=6e-08 w=1.26e-06 $X=42275 $Y=29007 $D=616
M1573 vss 284 r_lwea vss hvtnfet l=6e-08 w=1.287e-06 $X=42275 $Y=30897 $D=616
M1574 vss 557 303 vss hvtnfet l=6e-08 w=6e-07 $X=42275 $Y=37277 $D=616
M1575 vss 553 304 vss hvtnfet l=6e-08 w=6e-07 $X=42275 $Y=38507 $D=616
M1576 vss 554 305 vss hvtnfet l=6e-08 w=6e-07 $X=42275 $Y=43737 $D=616
M1577 vss 558 306 vss hvtnfet l=6e-08 w=6e-07 $X=42275 $Y=44967 $D=616
M1578 vss 559 307 vss hvtnfet l=6e-08 w=6e-07 $X=42275 $Y=50197 $D=616
M1579 303 557 vss vss hvtnfet l=6e-08 w=6e-07 $X=42535 $Y=37277 $D=616
M1580 vdd 5 15 vdd hvtpfet l=6e-08 w=1.2e-06 $X=965 $Y=35277 $D=636
M1581 11 1 vdd vdd hvtpfet l=6e-08 w=1.2e-06 $X=1225 $Y=1736 $D=636
M1582 12 2 vdd vdd hvtpfet l=6e-08 w=1.2e-06 $X=1225 $Y=3566 $D=636
M1583 13 3 vdd vdd hvtpfet l=6e-08 w=1.2e-06 $X=1225 $Y=8196 $D=636
M1584 14 4 vdd vdd hvtpfet l=6e-08 w=1.2e-06 $X=1225 $Y=10026 $D=636
M1585 lb_tm_preb_n 20 vdd vdd hvtpfet l=6e-08 w=2.145e-06 $X=1225 $Y=14887 $D=636
M1586 lt_tm_preb_n 21 vdd vdd hvtpfet l=6e-08 w=2.145e-06 $X=1225 $Y=17659 $D=636
M1587 vdd 8 l_clk_dqb vdd hvtpfet l=6e-08 w=2.1e-06 $X=1225 $Y=23621 $D=636
M1588 vdd 9 l_clk_dqb_n vdd hvtpfet l=6e-08 w=2.1e-06 $X=1225 $Y=26587 $D=636
M1589 l_lweb 10 vdd vdd hvtpfet l=6e-08 w=2.145e-06 $X=1225 $Y=32504 $D=636
M1590 15 5 vdd vdd hvtpfet l=6e-08 w=1.2e-06 $X=1225 $Y=35277 $D=636
M1591 16 4 vdd vdd hvtpfet l=6e-08 w=1.2e-06 $X=1225 $Y=39907 $D=636
M1592 17 3 vdd vdd hvtpfet l=6e-08 w=1.2e-06 $X=1225 $Y=41737 $D=636
M1593 18 6 vdd vdd hvtpfet l=6e-08 w=1.2e-06 $X=1225 $Y=46367 $D=636
M1594 19 7 vdd vdd hvtpfet l=6e-08 w=1.2e-06 $X=1225 $Y=48197 $D=636
M1595 vdd 20 lb_tm_preb_n vdd hvtpfet l=6e-08 w=2.145e-06 $X=1485 $Y=14887 $D=636
M1596 vdd 21 lt_tm_preb_n vdd hvtpfet l=6e-08 w=2.145e-06 $X=1485 $Y=17659 $D=636
M1597 l_clk_dqb 8 vdd vdd hvtpfet l=6e-08 w=2.1e-06 $X=1485 $Y=23621 $D=636
M1598 l_clk_dqb_n 9 vdd vdd hvtpfet l=6e-08 w=2.1e-06 $X=1485 $Y=26587 $D=636
M1599 vdd 10 l_lweb vdd hvtpfet l=6e-08 w=2.145e-06 $X=1485 $Y=32504 $D=636
M1600 lb_cb<0> 11 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=1735 $Y=1506 $D=636
M1601 lb_cb<2> 12 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=1735 $Y=3566 $D=636
M1602 lb_mb<0> 13 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=1735 $Y=7966 $D=636
M1603 lb_mb<2> 14 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=1735 $Y=10026 $D=636
M1604 l_saeb_n 15 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=1735 $Y=35277 $D=636
M1605 lt_mb<2> 16 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=1735 $Y=39677 $D=636
M1606 lt_mb<0> 17 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=1735 $Y=41737 $D=636
M1607 lt_cb<2> 18 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=1735 $Y=46137 $D=636
M1608 lt_cb<0> 19 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=1735 $Y=48197 $D=636
M1609 vdd 8 l_clk_dqb vdd hvtpfet l=6e-08 w=2.1e-06 $X=1745 $Y=23621 $D=636
M1610 vdd 9 l_clk_dqb_n vdd hvtpfet l=6e-08 w=2.1e-06 $X=1745 $Y=26587 $D=636
M1611 vdd 11 lb_cb<0> vdd hvtpfet l=6e-08 w=1.43e-06 $X=1995 $Y=1506 $D=636
M1612 vdd 12 lb_cb<2> vdd hvtpfet l=6e-08 w=1.43e-06 $X=1995 $Y=3566 $D=636
M1613 vdd 13 lb_mb<0> vdd hvtpfet l=6e-08 w=1.43e-06 $X=1995 $Y=7966 $D=636
M1614 vdd 14 lb_mb<2> vdd hvtpfet l=6e-08 w=1.43e-06 $X=1995 $Y=10026 $D=636
M1615 vdd 24 20 vdd hvtpfet l=6e-08 w=1.2e-06 $X=1995 $Y=15067 $D=636
M1616 vdd 25 21 vdd hvtpfet l=6e-08 w=1.2e-06 $X=1995 $Y=18424 $D=636
M1617 vdd 15 l_saeb_n vdd hvtpfet l=6e-08 w=1.43e-06 $X=1995 $Y=35277 $D=636
M1618 vdd 16 lt_mb<2> vdd hvtpfet l=6e-08 w=1.43e-06 $X=1995 $Y=39677 $D=636
M1619 vdd 17 lt_mb<0> vdd hvtpfet l=6e-08 w=1.43e-06 $X=1995 $Y=41737 $D=636
M1620 vdd 18 lt_cb<2> vdd hvtpfet l=6e-08 w=1.43e-06 $X=1995 $Y=46137 $D=636
M1621 vdd 19 lt_cb<0> vdd hvtpfet l=6e-08 w=1.43e-06 $X=1995 $Y=48197 $D=636
M1622 8 clkb vdd vdd hvtpfet l=6e-08 w=2.1e-06 $X=2005 $Y=23621 $D=636
M1623 9 23 vdd vdd hvtpfet l=6e-08 w=2.1e-06 $X=2005 $Y=26587 $D=636
M1624 lb_cb<0> 11 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=2255 $Y=1506 $D=636
M1625 lb_cb<2> 12 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=2255 $Y=3566 $D=636
M1626 lb_mb<0> 13 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=2255 $Y=7966 $D=636
M1627 lb_mb<2> 14 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=2255 $Y=10026 $D=636
M1628 l_saeb_n 15 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=2255 $Y=35277 $D=636
M1629 lt_mb<2> 16 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=2255 $Y=39677 $D=636
M1630 lt_mb<0> 17 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=2255 $Y=41737 $D=636
M1631 lt_cb<2> 18 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=2255 $Y=46137 $D=636
M1632 lt_cb<0> 19 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=2255 $Y=48197 $D=636
M1633 vdd 15 l_saeb_n vdd hvtpfet l=6e-08 w=1.43e-06 $X=2515 $Y=35277 $D=636
M1634 vdd 34 lb_cb<1> vdd hvtpfet l=6e-08 w=1.43e-06 $X=2765 $Y=1506 $D=636
M1635 vdd 35 lb_cb<3> vdd hvtpfet l=6e-08 w=1.43e-06 $X=2765 $Y=3566 $D=636
M1636 vdd 36 lb_mb<1> vdd hvtpfet l=6e-08 w=1.43e-06 $X=2765 $Y=7966 $D=636
M1637 vdd 37 lb_mb<3> vdd hvtpfet l=6e-08 w=1.43e-06 $X=2765 $Y=10026 $D=636
M1638 vdd 39 lt_mb<3> vdd hvtpfet l=6e-08 w=1.43e-06 $X=2765 $Y=39677 $D=636
M1639 vdd 40 lt_mb<1> vdd hvtpfet l=6e-08 w=1.43e-06 $X=2765 $Y=41737 $D=636
M1640 vdd 41 lt_cb<3> vdd hvtpfet l=6e-08 w=1.43e-06 $X=2765 $Y=46137 $D=636
M1641 vdd 42 lt_cb<1> vdd hvtpfet l=6e-08 w=1.43e-06 $X=2765 $Y=48197 $D=636
M1642 l_saeb_n 15 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=2775 $Y=35277 $D=636
M1643 26 28 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=2821 $Y=15321 $D=636
M1644 1145 26 vdd vdd hvtpfet l=6e-08 w=2.74e-07 $X=2821 $Y=16069 $D=636
M1645 1146 4 vdd vdd hvtpfet l=6e-08 w=2.74e-07 $X=2821 $Y=20589 $D=636
M1646 4 29 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=2821 $Y=21405 $D=636
M1647 27 30 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=2821 $Y=22241 $D=636
M1648 1147 27 vdd vdd hvtpfet l=6e-08 w=2.74e-07 $X=2821 $Y=22989 $D=636
M1649 1148 3 vdd vdd hvtpfet l=6e-08 w=2.74e-07 $X=2821 $Y=27509 $D=636
M1650 3 31 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=2821 $Y=28325 $D=636
M1651 lb_cb<1> 34 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=3025 $Y=1506 $D=636
M1652 lb_cb<3> 35 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=3025 $Y=3566 $D=636
M1653 lb_mb<1> 36 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=3025 $Y=7966 $D=636
M1654 lb_mb<3> 37 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=3025 $Y=10026 $D=636
M1655 lt_mb<3> 39 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=3025 $Y=39677 $D=636
M1656 lt_mb<1> 40 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=3025 $Y=41737 $D=636
M1657 lt_cb<3> 41 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=3025 $Y=46137 $D=636
M1658 lt_cb<1> 42 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=3025 $Y=48197 $D=636
M1659 vdd 28 26 vdd hvtpfet l=6e-08 w=2.06e-07 $X=3081 $Y=15321 $D=636
M1660 28 43 1145 vdd hvtpfet l=6e-08 w=2.74e-07 $X=3081 $Y=16069 $D=636
M1661 29 43 1146 vdd hvtpfet l=6e-08 w=2.74e-07 $X=3081 $Y=20589 $D=636
M1662 vdd 29 4 vdd hvtpfet l=6e-08 w=2.06e-07 $X=3081 $Y=21405 $D=636
M1663 vdd 30 27 vdd hvtpfet l=6e-08 w=2.06e-07 $X=3081 $Y=22241 $D=636
M1664 30 43 1147 vdd hvtpfet l=6e-08 w=2.74e-07 $X=3081 $Y=22989 $D=636
M1665 31 43 1148 vdd hvtpfet l=6e-08 w=2.74e-07 $X=3081 $Y=27509 $D=636
M1666 vdd 31 3 vdd hvtpfet l=6e-08 w=2.06e-07 $X=3081 $Y=28325 $D=636
M1667 vdd 34 lb_cb<1> vdd hvtpfet l=6e-08 w=1.43e-06 $X=3285 $Y=1506 $D=636
M1668 vdd 35 lb_cb<3> vdd hvtpfet l=6e-08 w=1.43e-06 $X=3285 $Y=3566 $D=636
M1669 vdd 36 lb_mb<1> vdd hvtpfet l=6e-08 w=1.43e-06 $X=3285 $Y=7966 $D=636
M1670 vdd 37 lb_mb<3> vdd hvtpfet l=6e-08 w=1.43e-06 $X=3285 $Y=10026 $D=636
M1671 vdd 51 l_sa_preb_n vdd hvtpfet l=6e-08 w=1.43e-06 $X=3285 $Y=35277 $D=636
M1672 vdd 39 lt_mb<3> vdd hvtpfet l=6e-08 w=1.43e-06 $X=3285 $Y=39677 $D=636
M1673 vdd 40 lt_mb<1> vdd hvtpfet l=6e-08 w=1.43e-06 $X=3285 $Y=41737 $D=636
M1674 vdd 41 lt_cb<3> vdd hvtpfet l=6e-08 w=1.43e-06 $X=3285 $Y=46137 $D=636
M1675 vdd 42 lt_cb<1> vdd hvtpfet l=6e-08 w=1.43e-06 $X=3285 $Y=48197 $D=636
M1676 vdd ab<2> 44 vdd hvtpfet l=6e-08 w=4.11e-07 $X=3396 $Y=14280 $D=636
M1677 l_sa_preb_n 51 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=3545 $Y=35277 $D=636
M1678 vdd clkb 43 vdd hvtpfet l=6e-08 w=6e-07 $X=3546 $Y=33747 $D=636
M1679 1149 33 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=3591 $Y=15520 $D=636
M1680 1150 33 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=3591 $Y=20589 $D=636
M1681 1151 33 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=3591 $Y=22440 $D=636
M1682 1152 33 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=3591 $Y=27509 $D=636
M1683 52 stclkb vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=3705 $Y=29937 $D=636
M1684 vdd 47 34 vdd hvtpfet l=6e-08 w=1.2e-06 $X=3795 $Y=1736 $D=636
M1685 vdd 48 35 vdd hvtpfet l=6e-08 w=1.2e-06 $X=3795 $Y=3566 $D=636
M1686 vdd 27 36 vdd hvtpfet l=6e-08 w=1.2e-06 $X=3795 $Y=8196 $D=636
M1687 vdd 26 37 vdd hvtpfet l=6e-08 w=1.2e-06 $X=3795 $Y=10026 $D=636
M1688 vdd 26 39 vdd hvtpfet l=6e-08 w=1.2e-06 $X=3795 $Y=39907 $D=636
M1689 vdd 27 40 vdd hvtpfet l=6e-08 w=1.2e-06 $X=3795 $Y=41737 $D=636
M1690 vdd 49 41 vdd hvtpfet l=6e-08 w=1.2e-06 $X=3795 $Y=46367 $D=636
M1691 vdd 50 42 vdd hvtpfet l=6e-08 w=1.2e-06 $X=3795 $Y=48197 $D=636
M1692 vdd 51 l_sa_preb_n vdd hvtpfet l=6e-08 w=1.43e-06 $X=3805 $Y=35277 $D=636
M1693 43 clkb vdd vdd hvtpfet l=6e-08 w=6e-07 $X=3806 $Y=33747 $D=636
M1694 28 45 1149 vdd hvtpfet l=6e-08 w=4.11e-07 $X=3861 $Y=15932 $D=636
M1695 29 45 1150 vdd hvtpfet l=6e-08 w=4.11e-07 $X=3861 $Y=20589 $D=636
M1696 30 46 1151 vdd hvtpfet l=6e-08 w=4.11e-07 $X=3861 $Y=22852 $D=636
M1697 31 46 1152 vdd hvtpfet l=6e-08 w=4.11e-07 $X=3861 $Y=27509 $D=636
M1698 53 44 vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=3906 $Y=14280 $D=636
M1699 vdd clkb 43 vdd hvtpfet l=6e-08 w=6e-07 $X=4066 $Y=33747 $D=636
M1700 1153 53 28 vdd hvtpfet l=6e-08 w=4.11e-07 $X=4121 $Y=15932 $D=636
M1701 1154 44 29 vdd hvtpfet l=6e-08 w=4.11e-07 $X=4121 $Y=20589 $D=636
M1702 1155 53 30 vdd hvtpfet l=6e-08 w=4.11e-07 $X=4121 $Y=22852 $D=636
M1703 1156 44 31 vdd hvtpfet l=6e-08 w=4.11e-07 $X=4121 $Y=27509 $D=636
M1704 1157 52 59 vdd hvtpfet l=6e-08 w=8.23e-07 $X=4215 $Y=29525 $D=636
M1705 vdd 55 51 vdd hvtpfet l=6e-08 w=1.2e-06 $X=4315 $Y=35277 $D=636
M1706 43 clkb vdd vdd hvtpfet l=6e-08 w=6e-07 $X=4326 $Y=33747 $D=636
M1707 vdd 33 1153 vdd hvtpfet l=6e-08 w=8.23e-07 $X=4391 $Y=15520 $D=636
M1708 vdd 33 1154 vdd hvtpfet l=6e-08 w=8.23e-07 $X=4391 $Y=20589 $D=636
M1709 vdd 33 1155 vdd hvtpfet l=6e-08 w=8.23e-07 $X=4391 $Y=22440 $D=636
M1710 vdd 33 1156 vdd hvtpfet l=6e-08 w=8.23e-07 $X=4391 $Y=27509 $D=636
M1711 vdd ab<3> 46 vdd hvtpfet l=6e-08 w=4.11e-07 $X=4416 $Y=14280 $D=636
M1712 vdd 56 1157 vdd hvtpfet l=6e-08 w=8.23e-07 $X=4475 $Y=29525 $D=636
M1713 b_pxab<0> 60 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=4550 $Y=1941 $D=636
M1714 60 61 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=4550 $Y=5141 $D=636
M1715 61 62 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=4550 $Y=8691 $D=636
M1716 vdd 57 62 vdd hvtpfet l=6e-08 w=4.11e-07 $X=4550 $Y=10156 $D=636
M1717 vdd 57 63 vdd hvtpfet l=6e-08 w=4.11e-07 $X=4550 $Y=40566 $D=636
M1718 64 63 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=4550 $Y=41842 $D=636
M1719 65 64 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=4550 $Y=44992 $D=636
M1720 t_pxab<0> 65 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=4550 $Y=46622 $D=636
M1721 vdd 60 b_pxab<0> vdd hvtpfet l=6e-08 w=2.57e-06 $X=4810 $Y=1941 $D=636
M1722 vdd 61 60 vdd hvtpfet l=6e-08 w=1e-06 $X=4810 $Y=5141 $D=636
M1723 vdd 62 61 vdd hvtpfet l=6e-08 w=6e-07 $X=4810 $Y=8691 $D=636
M1724 62 24 vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=4810 $Y=10156 $D=636
M1725 63 25 vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=4810 $Y=40566 $D=636
M1726 vdd 63 64 vdd hvtpfet l=6e-08 w=6e-07 $X=4810 $Y=41842 $D=636
M1727 vdd 64 65 vdd hvtpfet l=6e-08 w=1e-06 $X=4810 $Y=44992 $D=636
M1728 vdd 65 t_pxab<0> vdd hvtpfet l=6e-08 w=2.57e-06 $X=4810 $Y=46622 $D=636
M1729 45 46 vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=4926 $Y=14280 $D=636
M1730 vdd 66 586 vdd hvtpfet l=1.4e-07 w=6.4e-07 $X=4939 $Y=36067 $D=636
M1731 1158 59 56 vdd hvtpfet l=6e-08 w=8.23e-07 $X=4985 $Y=29525 $D=636
M1732 vdd 58 587 vdd hvtpfet l=6e-08 w=6.4e-07 $X=5069 $Y=33468 $D=636
M1733 67 73 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=5141 $Y=15321 $D=636
M1734 1159 67 vdd vdd hvtpfet l=6e-08 w=2.74e-07 $X=5141 $Y=16069 $D=636
M1735 1160 68 vdd vdd hvtpfet l=6e-08 w=2.74e-07 $X=5141 $Y=20589 $D=636
M1736 68 74 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=5141 $Y=21405 $D=636
M1737 69 75 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=5141 $Y=22241 $D=636
M1738 1161 69 vdd vdd hvtpfet l=6e-08 w=2.74e-07 $X=5141 $Y=22989 $D=636
M1739 1162 57 vdd vdd hvtpfet l=6e-08 w=2.74e-07 $X=5141 $Y=27509 $D=636
M1740 57 76 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=5141 $Y=28325 $D=636
M1741 vdd 70 1158 vdd hvtpfet l=6e-08 w=8.23e-07 $X=5245 $Y=29525 $D=636
M1742 66 71 vdd vdd hvtpfet l=1.4e-07 w=6.4e-07 $X=5279 $Y=36067 $D=636
M1743 b_pxab<1> 78 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=5320 $Y=1941 $D=636
M1744 78 79 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=5320 $Y=5141 $D=636
M1745 79 80 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=5320 $Y=8691 $D=636
M1746 vdd 24 80 vdd hvtpfet l=6e-08 w=4.11e-07 $X=5320 $Y=10156 $D=636
M1747 vdd 25 81 vdd hvtpfet l=6e-08 w=4.11e-07 $X=5320 $Y=40566 $D=636
M1748 82 81 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=5320 $Y=41842 $D=636
M1749 83 82 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=5320 $Y=44992 $D=636
M1750 t_pxab<1> 83 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=5320 $Y=46622 $D=636
M1751 vdd 73 67 vdd hvtpfet l=6e-08 w=2.06e-07 $X=5401 $Y=15321 $D=636
M1752 73 43 1159 vdd hvtpfet l=6e-08 w=2.74e-07 $X=5401 $Y=16069 $D=636
M1753 74 43 1160 vdd hvtpfet l=6e-08 w=2.74e-07 $X=5401 $Y=20589 $D=636
M1754 vdd 74 68 vdd hvtpfet l=6e-08 w=2.06e-07 $X=5401 $Y=21405 $D=636
M1755 vdd 75 69 vdd hvtpfet l=6e-08 w=2.06e-07 $X=5401 $Y=22241 $D=636
M1756 75 43 1161 vdd hvtpfet l=6e-08 w=2.74e-07 $X=5401 $Y=22989 $D=636
M1757 76 43 1162 vdd hvtpfet l=6e-08 w=2.74e-07 $X=5401 $Y=27509 $D=636
M1758 vdd 76 57 vdd hvtpfet l=6e-08 w=2.06e-07 $X=5401 $Y=28325 $D=636
M1759 vdd 72 5 vdd hvtpfet l=6e-08 w=6.4e-07 $X=5579 $Y=33693 $D=636
M1760 vdd 78 b_pxab<1> vdd hvtpfet l=6e-08 w=2.57e-06 $X=5580 $Y=1941 $D=636
M1761 vdd 79 78 vdd hvtpfet l=6e-08 w=1e-06 $X=5580 $Y=5141 $D=636
M1762 vdd 80 79 vdd hvtpfet l=6e-08 w=6e-07 $X=5580 $Y=8691 $D=636
M1763 80 69 vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=5580 $Y=10156 $D=636
M1764 81 69 vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=5580 $Y=40566 $D=636
M1765 vdd 81 82 vdd hvtpfet l=6e-08 w=6e-07 $X=5580 $Y=41842 $D=636
M1766 vdd 82 83 vdd hvtpfet l=6e-08 w=1e-06 $X=5580 $Y=44992 $D=636
M1767 vdd 83 t_pxab<1> vdd hvtpfet l=6e-08 w=2.57e-06 $X=5580 $Y=46622 $D=636
M1768 vdd ab<5> 86 vdd hvtpfet l=6e-08 w=4.11e-07 $X=5716 $Y=14280 $D=636
M1769 5 85 vdd vdd hvtpfet l=6e-08 w=6.4e-07 $X=5839 $Y=33693 $D=636
M1770 1163 33 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=5911 $Y=15520 $D=636
M1771 1164 33 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=5911 $Y=20589 $D=636
M1772 1165 33 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=5911 $Y=22440 $D=636
M1773 1166 33 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=5911 $Y=27509 $D=636
M1774 70 clkb vdd vdd hvtpfet l=6e-08 w=1.2e-06 $X=6015 $Y=29148 $D=636
M1775 592 ddqb 71 vdd hvtpfet l=6e-08 w=6.4e-07 $X=6079 $Y=35802 $D=636
M1776 b_pxab<2> 90 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=6090 $Y=1941 $D=636
M1777 90 91 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=6090 $Y=5141 $D=636
M1778 91 92 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=6090 $Y=8691 $D=636
M1779 vdd 68 92 vdd hvtpfet l=6e-08 w=4.11e-07 $X=6090 $Y=10156 $D=636
M1780 vdd 68 93 vdd hvtpfet l=6e-08 w=4.11e-07 $X=6090 $Y=40566 $D=636
M1781 94 93 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=6090 $Y=41842 $D=636
M1782 95 94 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=6090 $Y=44992 $D=636
M1783 t_pxab<2> 95 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=6090 $Y=46622 $D=636
M1784 73 87 1163 vdd hvtpfet l=6e-08 w=4.11e-07 $X=6181 $Y=15932 $D=636
M1785 74 87 1164 vdd hvtpfet l=6e-08 w=4.11e-07 $X=6181 $Y=20589 $D=636
M1786 75 88 1165 vdd hvtpfet l=6e-08 w=4.11e-07 $X=6181 $Y=22852 $D=636
M1787 76 88 1166 vdd hvtpfet l=6e-08 w=4.11e-07 $X=6181 $Y=27509 $D=636
M1788 97 86 vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=6226 $Y=14280 $D=636
M1789 vdd ddqb_n 592 vdd hvtpfet l=6e-08 w=6.4e-07 $X=6339 $Y=35802 $D=636
M1790 vdd 90 b_pxab<2> vdd hvtpfet l=6e-08 w=2.57e-06 $X=6350 $Y=1941 $D=636
M1791 vdd 91 90 vdd hvtpfet l=6e-08 w=1e-06 $X=6350 $Y=5141 $D=636
M1792 vdd 92 91 vdd hvtpfet l=6e-08 w=6e-07 $X=6350 $Y=8691 $D=636
M1793 92 24 vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=6350 $Y=10156 $D=636
M1794 93 25 vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=6350 $Y=40566 $D=636
M1795 vdd 93 94 vdd hvtpfet l=6e-08 w=6e-07 $X=6350 $Y=41842 $D=636
M1796 vdd 94 95 vdd hvtpfet l=6e-08 w=1e-06 $X=6350 $Y=44992 $D=636
M1797 vdd 95 t_pxab<2> vdd hvtpfet l=6e-08 w=2.57e-06 $X=6350 $Y=46622 $D=636
M1798 1167 97 73 vdd hvtpfet l=6e-08 w=4.11e-07 $X=6441 $Y=15932 $D=636
M1799 1168 86 74 vdd hvtpfet l=6e-08 w=4.11e-07 $X=6441 $Y=20589 $D=636
M1800 1169 97 75 vdd hvtpfet l=6e-08 w=4.11e-07 $X=6441 $Y=22852 $D=636
M1801 1170 86 76 vdd hvtpfet l=6e-08 w=4.11e-07 $X=6441 $Y=27509 $D=636
M1802 85 89 vdd vdd hvtpfet l=6e-08 w=6.4e-07 $X=6524 $Y=33693 $D=636
M1803 142 clkb vdd vdd hvtpfet l=6e-08 w=8e-07 $X=6525 $Y=29548 $D=636
M1804 vdd 33 1167 vdd hvtpfet l=6e-08 w=8.23e-07 $X=6711 $Y=15520 $D=636
M1805 vdd 33 1168 vdd hvtpfet l=6e-08 w=8.23e-07 $X=6711 $Y=20589 $D=636
M1806 vdd 33 1169 vdd hvtpfet l=6e-08 w=8.23e-07 $X=6711 $Y=22440 $D=636
M1807 vdd 33 1170 vdd hvtpfet l=6e-08 w=8.23e-07 $X=6711 $Y=27509 $D=636
M1808 vdd ab<6> 88 vdd hvtpfet l=6e-08 w=4.11e-07 $X=6736 $Y=14280 $D=636
M1809 vdd clkb 142 vdd hvtpfet l=6e-08 w=8e-07 $X=6785 $Y=29548 $D=636
M1810 b_pxab<3> 99 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=6860 $Y=1941 $D=636
M1811 99 100 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=6860 $Y=5141 $D=636
M1812 100 101 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=6860 $Y=8691 $D=636
M1813 vdd 24 101 vdd hvtpfet l=6e-08 w=4.11e-07 $X=6860 $Y=10156 $D=636
M1814 vdd 25 102 vdd hvtpfet l=6e-08 w=4.11e-07 $X=6860 $Y=40566 $D=636
M1815 103 102 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=6860 $Y=41842 $D=636
M1816 104 103 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=6860 $Y=44992 $D=636
M1817 t_pxab<3> 104 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=6860 $Y=46622 $D=636
M1818 109 85 vdd vdd hvtpfet l=6e-08 w=6.4e-07 $X=7034 $Y=33468 $D=636
M1819 89 71 vdd vdd hvtpfet l=6e-08 w=6.4e-07 $X=7069 $Y=35802 $D=636
M1820 vdd 99 b_pxab<3> vdd hvtpfet l=6e-08 w=2.57e-06 $X=7120 $Y=1941 $D=636
M1821 vdd 100 99 vdd hvtpfet l=6e-08 w=1e-06 $X=7120 $Y=5141 $D=636
M1822 vdd 101 100 vdd hvtpfet l=6e-08 w=6e-07 $X=7120 $Y=8691 $D=636
M1823 101 67 vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=7120 $Y=10156 $D=636
M1824 102 67 vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=7120 $Y=40566 $D=636
M1825 vdd 102 103 vdd hvtpfet l=6e-08 w=6e-07 $X=7120 $Y=41842 $D=636
M1826 vdd 103 104 vdd hvtpfet l=6e-08 w=1e-06 $X=7120 $Y=44992 $D=636
M1827 vdd 104 t_pxab<3> vdd hvtpfet l=6e-08 w=2.57e-06 $X=7120 $Y=46622 $D=636
M1828 87 88 vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=7246 $Y=14280 $D=636
M1829 142 59 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=7295 $Y=29548 $D=636
M1830 105 111 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=7461 $Y=15321 $D=636
M1831 1171 105 vdd vdd hvtpfet l=6e-08 w=2.74e-07 $X=7461 $Y=16069 $D=636
M1832 1172 106 vdd vdd hvtpfet l=6e-08 w=2.74e-07 $X=7461 $Y=20589 $D=636
M1833 106 112 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=7461 $Y=21405 $D=636
M1834 107 113 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=7461 $Y=22241 $D=636
M1835 1173 107 vdd vdd hvtpfet l=6e-08 w=2.74e-07 $X=7461 $Y=22989 $D=636
M1836 1174 108 vdd vdd hvtpfet l=6e-08 w=2.74e-07 $X=7461 $Y=27509 $D=636
M1837 108 114 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=7461 $Y=28325 $D=636
M1838 vdd 59 142 vdd hvtpfet l=6e-08 w=8e-07 $X=7555 $Y=29548 $D=636
M1839 vdd 110 89 vdd hvtpfet l=1.2e-07 w=3e-07 $X=7579 $Y=36382 $D=636
M1840 b_pxbb_n<0> 115 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=7630 $Y=1941 $D=636
M1841 115 116 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=7630 $Y=5141 $D=636
M1842 116 107 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=7630 $Y=8691 $D=636
M1843 117 107 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=7630 $Y=41842 $D=636
M1844 118 117 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=7630 $Y=44992 $D=636
M1845 t_pxbb_n<0> 118 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=7630 $Y=46622 $D=636
M1846 vdd 109 119 vdd hvtpfet l=6e-08 w=5e-07 $X=7634 $Y=33503 $D=636
M1847 vdd 111 105 vdd hvtpfet l=6e-08 w=2.06e-07 $X=7721 $Y=15321 $D=636
M1848 111 43 1171 vdd hvtpfet l=6e-08 w=2.74e-07 $X=7721 $Y=16069 $D=636
M1849 112 43 1172 vdd hvtpfet l=6e-08 w=2.74e-07 $X=7721 $Y=20589 $D=636
M1850 vdd 112 106 vdd hvtpfet l=6e-08 w=2.06e-07 $X=7721 $Y=21405 $D=636
M1851 vdd 113 107 vdd hvtpfet l=6e-08 w=2.06e-07 $X=7721 $Y=22241 $D=636
M1852 113 43 1173 vdd hvtpfet l=6e-08 w=2.74e-07 $X=7721 $Y=22989 $D=636
M1853 114 43 1174 vdd hvtpfet l=6e-08 w=2.74e-07 $X=7721 $Y=27509 $D=636
M1854 vdd 114 108 vdd hvtpfet l=6e-08 w=2.06e-07 $X=7721 $Y=28325 $D=636
M1855 vdd 115 b_pxbb_n<0> vdd hvtpfet l=6e-08 w=2.57e-06 $X=7890 $Y=1941 $D=636
M1856 vdd 116 115 vdd hvtpfet l=6e-08 w=1e-06 $X=7890 $Y=5141 $D=636
M1857 vdd 107 116 vdd hvtpfet l=6e-08 w=6e-07 $X=7890 $Y=8691 $D=636
M1858 vdd 107 117 vdd hvtpfet l=6e-08 w=6e-07 $X=7890 $Y=41842 $D=636
M1859 vdd 117 118 vdd hvtpfet l=6e-08 w=1e-06 $X=7890 $Y=44992 $D=636
M1860 vdd 118 t_pxbb_n<0> vdd hvtpfet l=6e-08 w=2.57e-06 $X=7890 $Y=46622 $D=636
M1861 120 119 vdd vdd hvtpfet l=2.5e-07 w=5e-07 $X=7894 $Y=33503 $D=636
M1862 110 89 vdd vdd hvtpfet l=6e-08 w=3e-07 $X=8149 $Y=36377 $D=636
M1863 1175 33 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=8231 $Y=15520 $D=636
M1864 1176 33 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=8231 $Y=20589 $D=636
M1865 1177 33 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=8231 $Y=22440 $D=636
M1866 1178 33 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=8231 $Y=27509 $D=636
M1867 b_pxbb_n<1> 125 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=8400 $Y=1941 $D=636
M1868 125 126 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=8400 $Y=5141 $D=636
M1869 126 108 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=8400 $Y=8691 $D=636
M1870 127 108 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=8400 $Y=41842 $D=636
M1871 128 127 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=8400 $Y=44992 $D=636
M1872 t_pxbb_n<1> 128 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=8400 $Y=46622 $D=636
M1873 vdd 122 121 vdd hvtpfet l=6e-08 w=4.11e-07 $X=8466 $Y=14280 $D=636
M1874 111 121 1175 vdd hvtpfet l=6e-08 w=4.11e-07 $X=8501 $Y=15932 $D=636
M1875 112 121 1176 vdd hvtpfet l=6e-08 w=4.11e-07 $X=8501 $Y=20589 $D=636
M1876 113 122 1177 vdd hvtpfet l=6e-08 w=4.11e-07 $X=8501 $Y=22852 $D=636
M1877 114 122 1178 vdd hvtpfet l=6e-08 w=4.11e-07 $X=8501 $Y=27509 $D=636
M1878 131 123 vdd vdd hvtpfet l=6e-08 w=2e-07 $X=8594 $Y=10756 $D=636
M1879 vdd 120 55 vdd hvtpfet l=6e-08 w=6.4e-07 $X=8619 $Y=33468 $D=636
M1880 602 124 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=8659 $Y=29348 $D=636
M1881 603 124 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=8659 $Y=35707 $D=636
M1882 vdd 125 b_pxbb_n<1> vdd hvtpfet l=6e-08 w=2.57e-06 $X=8660 $Y=1941 $D=636
M1883 vdd 126 125 vdd hvtpfet l=6e-08 w=1e-06 $X=8660 $Y=5141 $D=636
M1884 vdd 108 126 vdd hvtpfet l=6e-08 w=6e-07 $X=8660 $Y=8691 $D=636
M1885 vdd 108 127 vdd hvtpfet l=6e-08 w=6e-07 $X=8660 $Y=41842 $D=636
M1886 vdd 127 128 vdd hvtpfet l=6e-08 w=1e-06 $X=8660 $Y=44992 $D=636
M1887 vdd 128 t_pxbb_n<1> vdd hvtpfet l=6e-08 w=2.57e-06 $X=8660 $Y=46622 $D=636
M1888 1179 129 111 vdd hvtpfet l=6e-08 w=4.11e-07 $X=8761 $Y=15932 $D=636
M1889 1180 129 112 vdd hvtpfet l=6e-08 w=4.11e-07 $X=8761 $Y=20589 $D=636
M1890 1181 129 113 vdd hvtpfet l=6e-08 w=4.11e-07 $X=8761 $Y=22852 $D=636
M1891 1182 129 114 vdd hvtpfet l=6e-08 w=4.11e-07 $X=8761 $Y=27509 $D=636
M1892 55 vdd vdd vdd hvtpfet l=6e-08 w=6.4e-07 $X=8879 $Y=33468 $D=636
M1893 vdd 124 602 vdd hvtpfet l=6e-08 w=1e-06 $X=8919 $Y=29348 $D=636
M1894 vdd 124 603 vdd hvtpfet l=6e-08 w=1e-06 $X=8919 $Y=35707 $D=636
M1895 122 ab<9> vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=8976 $Y=14280 $D=636
M1896 vdd 33 1179 vdd hvtpfet l=6e-08 w=8.23e-07 $X=9031 $Y=15520 $D=636
M1897 vdd 33 1180 vdd hvtpfet l=6e-08 w=8.23e-07 $X=9031 $Y=20589 $D=636
M1898 vdd 33 1181 vdd hvtpfet l=6e-08 w=8.23e-07 $X=9031 $Y=22440 $D=636
M1899 vdd 33 1182 vdd hvtpfet l=6e-08 w=8.23e-07 $X=9031 $Y=27509 $D=636
M1900 b_pxbb_n<2> 135 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=9170 $Y=1941 $D=636
M1901 135 136 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=9170 $Y=5141 $D=636
M1902 136 137 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=9170 $Y=8691 $D=636
M1903 138 137 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=9170 $Y=41842 $D=636
M1904 139 138 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=9170 $Y=44992 $D=636
M1905 t_pxbb_n<2> 139 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=9170 $Y=46622 $D=636
M1906 dwlb<0> 142 602 vdd hvtpfet l=6e-08 w=1e-06 $X=9429 $Y=29348 $D=636
M1907 25 143 603 vdd hvtpfet l=6e-08 w=1e-06 $X=9429 $Y=35707 $D=636
M1908 vdd 135 b_pxbb_n<2> vdd hvtpfet l=6e-08 w=2.57e-06 $X=9430 $Y=1941 $D=636
M1909 vdd 136 135 vdd hvtpfet l=6e-08 w=1e-06 $X=9430 $Y=5141 $D=636
M1910 vdd 137 136 vdd hvtpfet l=6e-08 w=6e-07 $X=9430 $Y=8691 $D=636
M1911 vdd 137 138 vdd hvtpfet l=6e-08 w=6e-07 $X=9430 $Y=41842 $D=636
M1912 vdd 138 139 vdd hvtpfet l=6e-08 w=1e-06 $X=9430 $Y=44992 $D=636
M1913 vdd 139 t_pxbb_n<2> vdd hvtpfet l=6e-08 w=2.57e-06 $X=9430 $Y=46622 $D=636
M1914 1183 132 111 vdd hvtpfet l=6e-08 w=4.11e-07 $X=9541 $Y=15932 $D=636
M1915 1184 133 112 vdd hvtpfet l=6e-08 w=4.11e-07 $X=9541 $Y=20589 $D=636
M1916 1185 132 113 vdd hvtpfet l=6e-08 w=4.11e-07 $X=9541 $Y=22852 $D=636
M1917 1186 133 114 vdd hvtpfet l=6e-08 w=4.11e-07 $X=9541 $Y=27509 $D=636
M1918 vdd 140 1 vdd hvtpfet l=6e-08 w=4e-07 $X=9586 $Y=10167 $D=636
M1919 vdd 141 7 vdd hvtpfet l=6e-08 w=4e-07 $X=9586 $Y=40566 $D=636
M1920 602 142 dwlb<0> vdd hvtpfet l=6e-08 w=1e-06 $X=9689 $Y=29348 $D=636
M1921 603 143 25 vdd hvtpfet l=6e-08 w=1e-06 $X=9689 $Y=35707 $D=636
M1922 vdd 33 1183 vdd hvtpfet l=6e-08 w=8.23e-07 $X=9811 $Y=15520 $D=636
M1923 vdd 33 1184 vdd hvtpfet l=6e-08 w=8.23e-07 $X=9811 $Y=20589 $D=636
M1924 vdd 33 1185 vdd hvtpfet l=6e-08 w=8.23e-07 $X=9811 $Y=22440 $D=636
M1925 vdd 33 1186 vdd hvtpfet l=6e-08 w=8.23e-07 $X=9811 $Y=27509 $D=636
M1926 b_pxbb_n<3> 146 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=9940 $Y=1941 $D=636
M1927 146 147 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=9940 $Y=5141 $D=636
M1928 147 148 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=9940 $Y=8691 $D=636
M1929 149 148 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=9940 $Y=41842 $D=636
M1930 150 149 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=9940 $Y=44992 $D=636
M1931 t_pxbb_n<3> 150 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=9940 $Y=46622 $D=636
M1932 vdd ab<8> 129 vdd hvtpfet l=6e-08 w=4.11e-07 $X=9986 $Y=14280 $D=636
M1933 1187 33 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=10071 $Y=15520 $D=636
M1934 1188 33 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=10071 $Y=20589 $D=636
M1935 1189 33 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=10071 $Y=22440 $D=636
M1936 1190 33 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=10071 $Y=27509 $D=636
M1937 vdd 145 140 vdd hvtpfet l=6e-08 w=4.11e-07 $X=10096 $Y=10156 $D=636
M1938 vdd 145 141 vdd hvtpfet l=6e-08 w=4.11e-07 $X=10096 $Y=40566 $D=636
M1939 dwlb<1> 142 608 vdd hvtpfet l=6e-08 w=1e-06 $X=10199 $Y=29348 $D=636
M1940 24 143 609 vdd hvtpfet l=6e-08 w=1e-06 $X=10199 $Y=35707 $D=636
M1941 vdd 146 b_pxbb_n<3> vdd hvtpfet l=6e-08 w=2.57e-06 $X=10200 $Y=1941 $D=636
M1942 vdd 147 146 vdd hvtpfet l=6e-08 w=1e-06 $X=10200 $Y=5141 $D=636
M1943 vdd 148 147 vdd hvtpfet l=6e-08 w=6e-07 $X=10200 $Y=8691 $D=636
M1944 vdd 148 149 vdd hvtpfet l=6e-08 w=6e-07 $X=10200 $Y=41842 $D=636
M1945 vdd 149 150 vdd hvtpfet l=6e-08 w=1e-06 $X=10200 $Y=44992 $D=636
M1946 vdd 150 t_pxbb_n<3> vdd hvtpfet l=6e-08 w=2.57e-06 $X=10200 $Y=46622 $D=636
M1947 160 129 vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=10246 $Y=14280 $D=636
M1948 168 132 1187 vdd hvtpfet l=6e-08 w=4.11e-07 $X=10341 $Y=15932 $D=636
M1949 169 133 1188 vdd hvtpfet l=6e-08 w=4.11e-07 $X=10341 $Y=20589 $D=636
M1950 170 132 1189 vdd hvtpfet l=6e-08 w=4.11e-07 $X=10341 $Y=22852 $D=636
M1951 171 133 1190 vdd hvtpfet l=6e-08 w=4.11e-07 $X=10341 $Y=27509 $D=636
M1952 140 dwlb<1> vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=10356 $Y=10156 $D=636
M1953 141 dwlb<0> vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=10356 $Y=40566 $D=636
M1954 vdd 153 124 vdd hvtpfet l=6e-08 w=8e-07 $X=10406 $Y=33493 $D=636
M1955 608 142 dwlb<1> vdd hvtpfet l=6e-08 w=1e-06 $X=10459 $Y=29348 $D=636
M1956 609 143 24 vdd hvtpfet l=6e-08 w=1e-06 $X=10459 $Y=35707 $D=636
M1957 b_pxbb_n<4> 156 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=10710 $Y=1941 $D=636
M1958 156 157 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=10710 $Y=5141 $D=636
M1959 157 105 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=10710 $Y=8691 $D=636
M1960 158 105 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=10710 $Y=41842 $D=636
M1961 159 158 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=10710 $Y=44992 $D=636
M1962 t_pxbb_n<4> 159 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=10710 $Y=46622 $D=636
M1963 vdd 132 133 vdd hvtpfet l=6e-08 w=4.11e-07 $X=10846 $Y=14280 $D=636
M1964 1191 33 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=10851 $Y=15520 $D=636
M1965 1192 33 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=10851 $Y=20589 $D=636
M1966 1193 33 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=10851 $Y=22440 $D=636
M1967 1194 33 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=10851 $Y=27509 $D=636
M1968 vdd dwlb<1> 162 vdd hvtpfet l=6e-08 w=4.11e-07 $X=10866 $Y=10156 $D=636
M1969 vdd dwlb<0> 163 vdd hvtpfet l=6e-08 w=4.11e-07 $X=10866 $Y=40566 $D=636
M1970 608 153 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=10969 $Y=29348 $D=636
M1971 609 153 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=10969 $Y=35707 $D=636
M1972 vdd 156 b_pxbb_n<4> vdd hvtpfet l=6e-08 w=2.57e-06 $X=10970 $Y=1941 $D=636
M1973 vdd 157 156 vdd hvtpfet l=6e-08 w=1e-06 $X=10970 $Y=5141 $D=636
M1974 vdd 105 157 vdd hvtpfet l=6e-08 w=6e-07 $X=10970 $Y=8691 $D=636
M1975 vdd 105 158 vdd hvtpfet l=6e-08 w=6e-07 $X=10970 $Y=41842 $D=636
M1976 vdd 158 159 vdd hvtpfet l=6e-08 w=1e-06 $X=10970 $Y=44992 $D=636
M1977 vdd 159 t_pxbb_n<4> vdd hvtpfet l=6e-08 w=2.57e-06 $X=10970 $Y=46622 $D=636
M1978 132 ab<7> vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=11106 $Y=14280 $D=636
M1979 153 154 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=11106 $Y=33493 $D=636
M1980 168 160 1191 vdd hvtpfet l=6e-08 w=4.11e-07 $X=11121 $Y=15932 $D=636
M1981 169 160 1192 vdd hvtpfet l=6e-08 w=4.11e-07 $X=11121 $Y=20589 $D=636
M1982 170 160 1193 vdd hvtpfet l=6e-08 w=4.11e-07 $X=11121 $Y=22852 $D=636
M1983 171 160 1194 vdd hvtpfet l=6e-08 w=4.11e-07 $X=11121 $Y=27509 $D=636
M1984 162 155 vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=11126 $Y=10156 $D=636
M1985 163 155 vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=11126 $Y=40566 $D=636
M1986 vdd 153 608 vdd hvtpfet l=6e-08 w=1e-06 $X=11229 $Y=29348 $D=636
M1987 vdd 153 609 vdd hvtpfet l=6e-08 w=1e-06 $X=11229 $Y=35707 $D=636
M1988 1195 121 168 vdd hvtpfet l=6e-08 w=4.11e-07 $X=11381 $Y=15932 $D=636
M1989 1196 121 169 vdd hvtpfet l=6e-08 w=4.11e-07 $X=11381 $Y=20589 $D=636
M1990 1197 122 170 vdd hvtpfet l=6e-08 w=4.11e-07 $X=11381 $Y=22852 $D=636
M1991 1198 122 171 vdd hvtpfet l=6e-08 w=4.11e-07 $X=11381 $Y=27509 $D=636
M1992 b_pxbb_n<5> 164 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=11480 $Y=1941 $D=636
M1993 164 165 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=11480 $Y=5141 $D=636
M1994 165 106 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=11480 $Y=8691 $D=636
M1995 166 106 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=11480 $Y=41842 $D=636
M1996 167 166 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=11480 $Y=44992 $D=636
M1997 t_pxbb_n<5> 167 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=11480 $Y=46622 $D=636
M1998 47 162 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=11636 $Y=10167 $D=636
M1999 50 163 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=11636 $Y=40566 $D=636
M2000 vdd 33 1195 vdd hvtpfet l=6e-08 w=8.23e-07 $X=11651 $Y=15520 $D=636
M2001 vdd 33 1196 vdd hvtpfet l=6e-08 w=8.23e-07 $X=11651 $Y=20589 $D=636
M2002 vdd 33 1197 vdd hvtpfet l=6e-08 w=8.23e-07 $X=11651 $Y=22440 $D=636
M2003 vdd 33 1198 vdd hvtpfet l=6e-08 w=8.23e-07 $X=11651 $Y=27509 $D=636
M2004 172 142 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=11739 $Y=29948 $D=636
M2005 vdd 164 b_pxbb_n<5> vdd hvtpfet l=6e-08 w=2.57e-06 $X=11740 $Y=1941 $D=636
M2006 vdd 165 164 vdd hvtpfet l=6e-08 w=1e-06 $X=11740 $Y=5141 $D=636
M2007 vdd 106 165 vdd hvtpfet l=6e-08 w=6e-07 $X=11740 $Y=8691 $D=636
M2008 vdd 106 166 vdd hvtpfet l=6e-08 w=6e-07 $X=11740 $Y=41842 $D=636
M2009 vdd 166 167 vdd hvtpfet l=6e-08 w=1e-06 $X=11740 $Y=44992 $D=636
M2010 vdd 167 t_pxbb_n<5> vdd hvtpfet l=6e-08 w=2.57e-06 $X=11740 $Y=46622 $D=636
M2011 vdd tm<0> dbl_pd_n<0> vdd hvtpfet l=6e-08 w=4.28e-07 $X=11746 $Y=14263 $D=636
M2012 616 172 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=11933 $Y=35707 $D=636
M2013 dbl_pd_n<0> tm<0> vdd vdd hvtpfet l=6e-08 w=4.28e-07 $X=12006 $Y=14263 $D=636
M2014 179 173 vdd vdd hvtpfet l=6e-08 w=3e-07 $X=12086 $Y=33468 $D=636
M2015 vdd 174 2 vdd hvtpfet l=6e-08 w=4e-07 $X=12146 $Y=10167 $D=636
M2016 vdd 175 6 vdd hvtpfet l=6e-08 w=4e-07 $X=12146 $Y=40566 $D=636
M2017 177 168 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=12161 $Y=15321 $D=636
M2018 1199 43 168 vdd hvtpfet l=6e-08 w=2.74e-07 $X=12161 $Y=16069 $D=636
M2019 1200 43 169 vdd hvtpfet l=6e-08 w=2.74e-07 $X=12161 $Y=20589 $D=636
M2020 178 169 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=12161 $Y=21405 $D=636
M2021 137 170 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=12161 $Y=22241 $D=636
M2022 1201 43 170 vdd hvtpfet l=6e-08 w=2.74e-07 $X=12161 $Y=22989 $D=636
M2023 1202 43 171 vdd hvtpfet l=6e-08 w=2.74e-07 $X=12161 $Y=27509 $D=636
M2024 148 171 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=12161 $Y=28325 $D=636
M2025 vdd 172 616 vdd hvtpfet l=6e-08 w=1e-06 $X=12193 $Y=35707 $D=636
M2026 b_pxbb_n<6> 180 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=12250 $Y=1941 $D=636
M2027 180 181 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=12250 $Y=5141 $D=636
M2028 181 177 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=12250 $Y=8691 $D=636
M2029 182 177 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=12250 $Y=41842 $D=636
M2030 183 182 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=12250 $Y=44992 $D=636
M2031 t_pxbb_n<6> 183 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=12250 $Y=46622 $D=636
M2032 vdd tm<0> dbl_pd_n<0> vdd hvtpfet l=6e-08 w=4.28e-07 $X=12266 $Y=14263 $D=636
M2033 vdd 142 184 vdd hvtpfet l=6e-08 w=5e-07 $X=12339 $Y=29813 $D=636
M2034 vdd 168 177 vdd hvtpfet l=6e-08 w=2.06e-07 $X=12421 $Y=15321 $D=636
M2035 vdd 177 1199 vdd hvtpfet l=6e-08 w=2.74e-07 $X=12421 $Y=16069 $D=636
M2036 vdd 178 1200 vdd hvtpfet l=6e-08 w=2.74e-07 $X=12421 $Y=20589 $D=636
M2037 vdd 169 178 vdd hvtpfet l=6e-08 w=2.06e-07 $X=12421 $Y=21405 $D=636
M2038 vdd 170 137 vdd hvtpfet l=6e-08 w=2.06e-07 $X=12421 $Y=22241 $D=636
M2039 vdd 137 1201 vdd hvtpfet l=6e-08 w=2.74e-07 $X=12421 $Y=22989 $D=636
M2040 vdd 148 1202 vdd hvtpfet l=6e-08 w=2.74e-07 $X=12421 $Y=27509 $D=636
M2041 vdd 171 148 vdd hvtpfet l=6e-08 w=2.06e-07 $X=12421 $Y=28325 $D=636
M2042 616 172 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=12453 $Y=35707 $D=636
M2043 vdd 180 b_pxbb_n<6> vdd hvtpfet l=6e-08 w=2.57e-06 $X=12510 $Y=1941 $D=636
M2044 vdd 181 180 vdd hvtpfet l=6e-08 w=1e-06 $X=12510 $Y=5141 $D=636
M2045 vdd 177 181 vdd hvtpfet l=6e-08 w=6e-07 $X=12510 $Y=8691 $D=636
M2046 vdd 177 182 vdd hvtpfet l=6e-08 w=6e-07 $X=12510 $Y=41842 $D=636
M2047 vdd 182 183 vdd hvtpfet l=6e-08 w=1e-06 $X=12510 $Y=44992 $D=636
M2048 vdd 183 t_pxbb_n<6> vdd hvtpfet l=6e-08 w=2.57e-06 $X=12510 $Y=46622 $D=636
M2049 615 179 186 vdd hvtpfet l=6e-08 w=6e-07 $X=12596 $Y=33468 $D=636
M2050 191 184 vdd vdd hvtpfet l=2.5e-07 w=5e-07 $X=12599 $Y=29813 $D=636
M2051 vdd 185 174 vdd hvtpfet l=6e-08 w=4.11e-07 $X=12656 $Y=10156 $D=636
M2052 vdd 185 175 vdd hvtpfet l=6e-08 w=4.11e-07 $X=12656 $Y=40566 $D=636
M2053 620 186 616 vdd hvtpfet l=6e-08 w=1e-06 $X=12713 $Y=35707 $D=636
M2054 vdd 131 dbl_pd_n<2> vdd hvtpfet l=6e-08 w=4.28e-07 $X=12776 $Y=14263 $D=636
M2055 vdd 191 615 vdd hvtpfet l=6e-08 w=6e-07 $X=12856 $Y=33468 $D=636
M2056 174 dwlb<1> vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=12916 $Y=10156 $D=636
M2057 175 dwlb<0> vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=12916 $Y=40566 $D=636
M2058 187 192 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=12931 $Y=15321 $D=636
M2059 1203 187 vdd vdd hvtpfet l=6e-08 w=2.74e-07 $X=12931 $Y=16069 $D=636
M2060 1204 188 vdd vdd hvtpfet l=6e-08 w=2.74e-07 $X=12931 $Y=20589 $D=636
M2061 188 193 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=12931 $Y=21405 $D=636
M2062 189 194 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=12931 $Y=22241 $D=636
M2063 1205 189 vdd vdd hvtpfet l=6e-08 w=2.74e-07 $X=12931 $Y=22989 $D=636
M2064 1206 190 vdd vdd hvtpfet l=6e-08 w=2.74e-07 $X=12931 $Y=27509 $D=636
M2065 190 195 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=12931 $Y=28325 $D=636
M2066 616 186 620 vdd hvtpfet l=6e-08 w=1e-06 $X=12973 $Y=35707 $D=636
M2067 b_pxbb_n<7> 196 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=13020 $Y=1941 $D=636
M2068 196 197 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=13020 $Y=5141 $D=636
M2069 197 178 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=13020 $Y=8691 $D=636
M2070 198 178 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=13020 $Y=41842 $D=636
M2071 199 198 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=13020 $Y=44992 $D=636
M2072 t_pxbb_n<7> 199 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=13020 $Y=46622 $D=636
M2073 dbl_pd_n<2> 131 vdd vdd hvtpfet l=6e-08 w=4.28e-07 $X=13036 $Y=14263 $D=636
M2074 vdd 192 187 vdd hvtpfet l=6e-08 w=2.06e-07 $X=13191 $Y=15321 $D=636
M2075 192 43 1203 vdd hvtpfet l=6e-08 w=2.74e-07 $X=13191 $Y=16069 $D=636
M2076 193 43 1204 vdd hvtpfet l=6e-08 w=2.74e-07 $X=13191 $Y=20589 $D=636
M2077 vdd 193 188 vdd hvtpfet l=6e-08 w=2.06e-07 $X=13191 $Y=21405 $D=636
M2078 vdd 194 189 vdd hvtpfet l=6e-08 w=2.06e-07 $X=13191 $Y=22241 $D=636
M2079 194 43 1205 vdd hvtpfet l=6e-08 w=2.74e-07 $X=13191 $Y=22989 $D=636
M2080 195 43 1206 vdd hvtpfet l=6e-08 w=2.74e-07 $X=13191 $Y=27509 $D=636
M2081 vdd 195 190 vdd hvtpfet l=6e-08 w=2.06e-07 $X=13191 $Y=28325 $D=636
M2082 620 186 616 vdd hvtpfet l=6e-08 w=1e-06 $X=13233 $Y=35707 $D=636
M2083 vdd 196 b_pxbb_n<7> vdd hvtpfet l=6e-08 w=2.57e-06 $X=13280 $Y=1941 $D=636
M2084 vdd 197 196 vdd hvtpfet l=6e-08 w=1e-06 $X=13280 $Y=5141 $D=636
M2085 vdd 178 197 vdd hvtpfet l=6e-08 w=6e-07 $X=13280 $Y=8691 $D=636
M2086 vdd 178 198 vdd hvtpfet l=6e-08 w=6e-07 $X=13280 $Y=41842 $D=636
M2087 vdd 198 199 vdd hvtpfet l=6e-08 w=1e-06 $X=13280 $Y=44992 $D=636
M2088 vdd 199 t_pxbb_n<7> vdd hvtpfet l=6e-08 w=2.57e-06 $X=13280 $Y=46622 $D=636
M2089 vdd 131 dbl_pd_n<2> vdd hvtpfet l=6e-08 w=4.28e-07 $X=13296 $Y=14263 $D=636
M2090 vdd tm<7> 203 vdd hvtpfet l=6e-08 w=3e-07 $X=13432 $Y=33468 $D=636
M2091 vdd 191 202 vdd hvtpfet l=6e-08 w=5e-07 $X=13459 $Y=29813 $D=636
M2092 143 200 620 vdd hvtpfet l=6e-08 w=1e-06 $X=13493 $Y=35707 $D=636
M2093 1207 33 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=13701 $Y=15520 $D=636
M2094 1208 33 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=13701 $Y=20589 $D=636
M2095 1209 33 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=13701 $Y=22440 $D=636
M2096 1210 33 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=13701 $Y=27509 $D=636
M2097 211 202 vdd vdd hvtpfet l=2.5e-07 w=5e-07 $X=13719 $Y=29813 $D=636
M2098 620 200 143 vdd hvtpfet l=6e-08 w=1e-06 $X=13753 $Y=35707 $D=636
M2099 b_pxcb_n<0> 206 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=13790 $Y=1941 $D=636
M2100 206 207 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=13790 $Y=5141 $D=636
M2101 207 189 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=13790 $Y=8691 $D=636
M2102 208 189 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=13790 $Y=41842 $D=636
M2103 209 208 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=13790 $Y=44992 $D=636
M2104 t_pxcb_n<0> 209 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=13790 $Y=46622 $D=636
M2105 vdd 205 204 vdd hvtpfet l=6e-08 w=4.11e-07 $X=13936 $Y=14280 $D=636
M2106 623 203 200 vdd hvtpfet l=6e-08 w=6e-07 $X=13942 $Y=33468 $D=636
M2107 192 204 1207 vdd hvtpfet l=6e-08 w=4.11e-07 $X=13971 $Y=15932 $D=636
M2108 193 204 1208 vdd hvtpfet l=6e-08 w=4.11e-07 $X=13971 $Y=20589 $D=636
M2109 194 205 1209 vdd hvtpfet l=6e-08 w=4.11e-07 $X=13971 $Y=22852 $D=636
M2110 195 205 1210 vdd hvtpfet l=6e-08 w=4.11e-07 $X=13971 $Y=27509 $D=636
M2111 143 200 620 vdd hvtpfet l=6e-08 w=1e-06 $X=14013 $Y=35707 $D=636
M2112 vdd 206 b_pxcb_n<0> vdd hvtpfet l=6e-08 w=2.57e-06 $X=14050 $Y=1941 $D=636
M2113 vdd 207 206 vdd hvtpfet l=6e-08 w=1e-06 $X=14050 $Y=5141 $D=636
M2114 vdd 189 207 vdd hvtpfet l=6e-08 w=6e-07 $X=14050 $Y=8691 $D=636
M2115 vdd 189 208 vdd hvtpfet l=6e-08 w=6e-07 $X=14050 $Y=41842 $D=636
M2116 vdd 208 209 vdd hvtpfet l=6e-08 w=1e-06 $X=14050 $Y=44992 $D=636
M2117 vdd 209 t_pxcb_n<0> vdd hvtpfet l=6e-08 w=2.57e-06 $X=14050 $Y=46622 $D=636
M2118 vdd 211 623 vdd hvtpfet l=6e-08 w=6e-07 $X=14202 $Y=33468 $D=636
M2119 vdd dwlb<1> 216 vdd hvtpfet l=6e-08 w=4.11e-07 $X=14216 $Y=10156 $D=636
M2120 vdd dwlb<0> 217 vdd hvtpfet l=6e-08 w=4.11e-07 $X=14216 $Y=40566 $D=636
M2121 1211 210 192 vdd hvtpfet l=6e-08 w=4.11e-07 $X=14231 $Y=15932 $D=636
M2122 1212 210 193 vdd hvtpfet l=6e-08 w=4.11e-07 $X=14231 $Y=20589 $D=636
M2123 1213 210 194 vdd hvtpfet l=6e-08 w=4.11e-07 $X=14231 $Y=22852 $D=636
M2124 1214 210 195 vdd hvtpfet l=6e-08 w=4.11e-07 $X=14231 $Y=27509 $D=636
M2125 205 ab<12> vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=14446 $Y=14280 $D=636
M2126 216 212 vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=14476 $Y=10156 $D=636
M2127 217 212 vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=14476 $Y=40566 $D=636
M2128 vdd 33 1211 vdd hvtpfet l=6e-08 w=8.23e-07 $X=14501 $Y=15520 $D=636
M2129 vdd 33 1212 vdd hvtpfet l=6e-08 w=8.23e-07 $X=14501 $Y=20589 $D=636
M2130 vdd 33 1213 vdd hvtpfet l=6e-08 w=8.23e-07 $X=14501 $Y=22440 $D=636
M2131 vdd 33 1214 vdd hvtpfet l=6e-08 w=8.23e-07 $X=14501 $Y=27509 $D=636
M2132 b_pxcb_n<1> 218 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=14560 $Y=1941 $D=636
M2133 218 219 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=14560 $Y=5141 $D=636
M2134 219 190 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=14560 $Y=8691 $D=636
M2135 220 190 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=14560 $Y=41842 $D=636
M2136 221 220 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=14560 $Y=44992 $D=636
M2137 t_pxcb_n<1> 221 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=14560 $Y=46622 $D=636
M2138 vdd 123 624 vdd hvtpfet l=6e-08 w=1.2e-06 $X=14796 $Y=29148 $D=636
M2139 vdd 218 b_pxcb_n<1> vdd hvtpfet l=6e-08 w=2.57e-06 $X=14820 $Y=1941 $D=636
M2140 vdd 219 218 vdd hvtpfet l=6e-08 w=1e-06 $X=14820 $Y=5141 $D=636
M2141 vdd 190 219 vdd hvtpfet l=6e-08 w=6e-07 $X=14820 $Y=8691 $D=636
M2142 vdd 190 220 vdd hvtpfet l=6e-08 w=6e-07 $X=14820 $Y=41842 $D=636
M2143 vdd 220 221 vdd hvtpfet l=6e-08 w=1e-06 $X=14820 $Y=44992 $D=636
M2144 vdd 221 t_pxcb_n<1> vdd hvtpfet l=6e-08 w=2.57e-06 $X=14820 $Y=46622 $D=636
M2145 vdd 72 58 vdd hvtpfet l=6e-08 w=4e-07 $X=14872 $Y=35682 $D=636
M2146 48 216 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=14986 $Y=10167 $D=636
M2147 49 217 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=14986 $Y=40566 $D=636
M2148 1215 213 192 vdd hvtpfet l=6e-08 w=4.11e-07 $X=15011 $Y=15932 $D=636
M2149 1216 214 193 vdd hvtpfet l=6e-08 w=4.11e-07 $X=15011 $Y=20589 $D=636
M2150 1217 213 194 vdd hvtpfet l=6e-08 w=4.11e-07 $X=15011 $Y=22852 $D=636
M2151 1218 214 195 vdd hvtpfet l=6e-08 w=4.11e-07 $X=15011 $Y=27509 $D=636
M2152 33 43 vdd vdd hvtpfet l=6e-08 w=7e-07 $X=15056 $Y=29648 $D=636
M2153 vdd 33 1215 vdd hvtpfet l=6e-08 w=8.23e-07 $X=15281 $Y=15520 $D=636
M2154 vdd 33 1216 vdd hvtpfet l=6e-08 w=8.23e-07 $X=15281 $Y=20589 $D=636
M2155 vdd 33 1217 vdd hvtpfet l=6e-08 w=8.23e-07 $X=15281 $Y=22440 $D=636
M2156 vdd 33 1218 vdd hvtpfet l=6e-08 w=8.23e-07 $X=15281 $Y=27509 $D=636
M2157 vdd 43 33 vdd hvtpfet l=6e-08 w=7e-07 $X=15316 $Y=29648 $D=636
M2158 b_pxcb_n<2> 223 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=15330 $Y=1941 $D=636
M2159 223 224 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=15330 $Y=5141 $D=636
M2160 224 225 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=15330 $Y=8691 $D=636
M2161 226 225 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=15330 $Y=41842 $D=636
M2162 227 226 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=15330 $Y=44992 $D=636
M2163 t_pxcb_n<2> 227 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=15330 $Y=46622 $D=636
M2164 vdd 229 72 vdd hvtpfet l=6e-08 w=4e-07 $X=15382 $Y=35682 $D=636
M2165 vdd ab<11> 210 vdd hvtpfet l=6e-08 w=4.11e-07 $X=15456 $Y=14280 $D=636
M2166 1219 33 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=15541 $Y=15520 $D=636
M2167 1220 33 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=15541 $Y=20589 $D=636
M2168 1221 33 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=15541 $Y=22440 $D=636
M2169 1222 33 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=15541 $Y=27509 $D=636
M2170 33 43 vdd vdd hvtpfet l=6e-08 w=7e-07 $X=15576 $Y=29648 $D=636
M2171 vdd 223 b_pxcb_n<2> vdd hvtpfet l=6e-08 w=2.57e-06 $X=15590 $Y=1941 $D=636
M2172 vdd 224 223 vdd hvtpfet l=6e-08 w=1e-06 $X=15590 $Y=5141 $D=636
M2173 vdd 225 224 vdd hvtpfet l=6e-08 w=6e-07 $X=15590 $Y=8691 $D=636
M2174 vdd 225 226 vdd hvtpfet l=6e-08 w=6e-07 $X=15590 $Y=41842 $D=636
M2175 vdd 226 227 vdd hvtpfet l=6e-08 w=1e-06 $X=15590 $Y=44992 $D=636
M2176 vdd 227 t_pxcb_n<2> vdd hvtpfet l=6e-08 w=2.57e-06 $X=15590 $Y=46622 $D=636
M2177 vdd 228 231 vdd hvtpfet l=6e-08 w=3.2e-07 $X=15621 $Y=33942 $D=636
M2178 72 172 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=15642 $Y=35682 $D=636
M2179 240 210 vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=15716 $Y=14280 $D=636
M2180 249 213 1219 vdd hvtpfet l=6e-08 w=4.11e-07 $X=15811 $Y=15932 $D=636
M2181 250 214 1220 vdd hvtpfet l=6e-08 w=4.11e-07 $X=15811 $Y=20589 $D=636
M2182 251 213 1221 vdd hvtpfet l=6e-08 w=4.11e-07 $X=15811 $Y=22852 $D=636
M2183 252 214 1222 vdd hvtpfet l=6e-08 w=4.11e-07 $X=15811 $Y=27509 $D=636
M2184 vdd 43 33 vdd hvtpfet l=6e-08 w=7e-07 $X=15836 $Y=29648 $D=636
M2185 631 tm<0> vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=15880 $Y=40177 $D=636
M2186 632 123 vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=15881 $Y=33942 $D=636
M2187 vdd tm<3> 242 vdd hvtpfet l=7e-08 w=4.8e-07 $X=16057 $Y=10476 $D=636
M2188 b_pxcb_n<3> 235 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=16100 $Y=1941 $D=636
M2189 235 236 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=16100 $Y=5141 $D=636
M2190 236 237 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=16100 $Y=8691 $D=636
M2191 238 237 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=16100 $Y=41842 $D=636
M2192 239 238 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=16100 $Y=44992 $D=636
M2193 t_pxcb_n<3> 239 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=16100 $Y=46622 $D=636
M2194 228 231 632 vdd hvtpfet l=6e-08 w=3.2e-07 $X=16141 $Y=33942 $D=636
M2195 vdd 213 214 vdd hvtpfet l=6e-08 w=4.11e-07 $X=16316 $Y=14280 $D=636
M2196 1225 33 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=16321 $Y=15520 $D=636
M2197 1226 33 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=16321 $Y=20589 $D=636
M2198 1227 33 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=16321 $Y=22440 $D=636
M2199 1228 33 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=16321 $Y=27509 $D=636
M2200 1223 232 vdd vdd hvtpfet l=6e-08 w=4.8e-07 $X=16322 $Y=35753 $D=636
M2201 243 tm<4> vdd vdd hvtpfet l=7e-08 w=4.8e-07 $X=16327 $Y=10476 $D=636
M2202 642 123 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=16346 $Y=29274 $D=636
M2203 vdd 235 b_pxcb_n<3> vdd hvtpfet l=6e-08 w=2.57e-06 $X=16360 $Y=1941 $D=636
M2204 vdd 236 235 vdd hvtpfet l=6e-08 w=1e-06 $X=16360 $Y=5141 $D=636
M2205 vdd 237 236 vdd hvtpfet l=6e-08 w=6e-07 $X=16360 $Y=8691 $D=636
M2206 vdd 237 238 vdd hvtpfet l=6e-08 w=6e-07 $X=16360 $Y=41842 $D=636
M2207 vdd 238 239 vdd hvtpfet l=6e-08 w=1e-06 $X=16360 $Y=44992 $D=636
M2208 vdd 239 t_pxcb_n<3> vdd hvtpfet l=6e-08 w=2.57e-06 $X=16360 $Y=46622 $D=636
M2209 1224 131 228 vdd hvtpfet l=6e-08 w=4.8e-07 $X=16401 $Y=33942 $D=636
M2210 213 ab<10> vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=16576 $Y=14280 $D=636
M2211 229 172 1223 vdd hvtpfet l=6e-08 w=4.8e-07 $X=16582 $Y=35753 $D=636
M2212 249 240 1225 vdd hvtpfet l=6e-08 w=4.11e-07 $X=16591 $Y=15932 $D=636
M2213 250 240 1226 vdd hvtpfet l=6e-08 w=4.11e-07 $X=16591 $Y=20589 $D=636
M2214 251 240 1227 vdd hvtpfet l=6e-08 w=4.11e-07 $X=16591 $Y=22852 $D=636
M2215 252 240 1228 vdd hvtpfet l=6e-08 w=4.11e-07 $X=16591 $Y=27509 $D=636
M2216 vdd 123 642 vdd hvtpfet l=6e-08 w=6e-07 $X=16606 $Y=29274 $D=636
M2217 vdd 123 1224 vdd hvtpfet l=6e-08 w=4.8e-07 $X=16661 $Y=33942 $D=636
M2218 637 tm<6> vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=16680 $Y=40177 $D=636
M2219 639 244 229 vdd hvtpfet l=6e-08 w=3.2e-07 $X=16842 $Y=35913 $D=636
M2220 1229 243 643 vdd hvtpfet l=6e-08 w=4.8e-07 $X=16847 $Y=10476 $D=636
M2221 1230 204 249 vdd hvtpfet l=6e-08 w=4.11e-07 $X=16851 $Y=15932 $D=636
M2222 1231 204 250 vdd hvtpfet l=6e-08 w=4.11e-07 $X=16851 $Y=20589 $D=636
M2223 1232 205 251 vdd hvtpfet l=6e-08 w=4.11e-07 $X=16851 $Y=22852 $D=636
M2224 1233 205 252 vdd hvtpfet l=6e-08 w=4.11e-07 $X=16851 $Y=27509 $D=636
M2225 642 123 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=16866 $Y=29274 $D=636
M2226 b_pxcb_n<4> 245 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=16870 $Y=1941 $D=636
M2227 245 246 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=16870 $Y=5141 $D=636
M2228 246 187 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=16870 $Y=8691 $D=636
M2229 247 187 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=16870 $Y=41842 $D=636
M2230 248 247 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=16870 $Y=44992 $D=636
M2231 t_pxcb_n<4> 248 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=16870 $Y=46622 $D=636
M2232 vdd 142 639 vdd hvtpfet l=6e-08 w=3.2e-07 $X=17102 $Y=35913 $D=636
M2233 vdd 242 1229 vdd hvtpfet l=6e-08 w=4.8e-07 $X=17107 $Y=10476 $D=636
M2234 vdd 33 1230 vdd hvtpfet l=6e-08 w=8.23e-07 $X=17121 $Y=15520 $D=636
M2235 vdd 33 1231 vdd hvtpfet l=6e-08 w=8.23e-07 $X=17121 $Y=20589 $D=636
M2236 vdd 33 1232 vdd hvtpfet l=6e-08 w=8.23e-07 $X=17121 $Y=22440 $D=636
M2237 vdd 33 1233 vdd hvtpfet l=6e-08 w=8.23e-07 $X=17121 $Y=27509 $D=636
M2238 vdd 123 642 vdd hvtpfet l=6e-08 w=6e-07 $X=17126 $Y=29274 $D=636
M2239 vdd 245 b_pxcb_n<4> vdd hvtpfet l=6e-08 w=2.57e-06 $X=17130 $Y=1941 $D=636
M2240 vdd 246 245 vdd hvtpfet l=6e-08 w=1e-06 $X=17130 $Y=5141 $D=636
M2241 vdd 187 246 vdd hvtpfet l=6e-08 w=6e-07 $X=17130 $Y=8691 $D=636
M2242 vdd 187 247 vdd hvtpfet l=6e-08 w=6e-07 $X=17130 $Y=41842 $D=636
M2243 vdd 247 248 vdd hvtpfet l=6e-08 w=1e-06 $X=17130 $Y=44992 $D=636
M2244 vdd 248 t_pxcb_n<4> vdd hvtpfet l=6e-08 w=2.57e-06 $X=17130 $Y=46622 $D=636
M2245 244 229 vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=17362 $Y=35913 $D=636
M2246 1234 242 vdd vdd hvtpfet l=6e-08 w=4.8e-07 $X=17617 $Y=10476 $D=636
M2247 253 249 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=17631 $Y=15321 $D=636
M2248 1235 43 249 vdd hvtpfet l=6e-08 w=2.74e-07 $X=17631 $Y=16069 $D=636
M2249 1236 43 250 vdd hvtpfet l=6e-08 w=2.74e-07 $X=17631 $Y=20589 $D=636
M2250 254 250 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=17631 $Y=21405 $D=636
M2251 225 251 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=17631 $Y=22241 $D=636
M2252 1237 43 251 vdd hvtpfet l=6e-08 w=2.74e-07 $X=17631 $Y=22989 $D=636
M2253 1238 43 252 vdd hvtpfet l=6e-08 w=2.74e-07 $X=17631 $Y=27509 $D=636
M2254 237 252 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=17631 $Y=28325 $D=636
M2255 b_pxcb_n<5> 255 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=17640 $Y=1941 $D=636
M2256 255 256 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=17640 $Y=5141 $D=636
M2257 256 188 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=17640 $Y=8691 $D=636
M2258 257 188 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=17640 $Y=41842 $D=636
M2259 258 257 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=17640 $Y=44992 $D=636
M2260 t_pxcb_n<5> 258 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=17640 $Y=46622 $D=636
M2261 23 clkb vdd vdd hvtpfet l=6e-08 w=9e-07 $X=17646 $Y=29274 $D=636
M2262 647 tm<4> 1234 vdd hvtpfet l=6e-08 w=4.8e-07 $X=17877 $Y=10476 $D=636
M2263 vdd 249 253 vdd hvtpfet l=6e-08 w=2.06e-07 $X=17891 $Y=15321 $D=636
M2264 vdd 253 1235 vdd hvtpfet l=6e-08 w=2.74e-07 $X=17891 $Y=16069 $D=636
M2265 vdd 254 1236 vdd hvtpfet l=6e-08 w=2.74e-07 $X=17891 $Y=20589 $D=636
M2266 vdd 250 254 vdd hvtpfet l=6e-08 w=2.06e-07 $X=17891 $Y=21405 $D=636
M2267 vdd 251 225 vdd hvtpfet l=6e-08 w=2.06e-07 $X=17891 $Y=22241 $D=636
M2268 vdd 225 1237 vdd hvtpfet l=6e-08 w=2.74e-07 $X=17891 $Y=22989 $D=636
M2269 vdd 237 1238 vdd hvtpfet l=6e-08 w=2.74e-07 $X=17891 $Y=27509 $D=636
M2270 vdd 252 237 vdd hvtpfet l=6e-08 w=2.06e-07 $X=17891 $Y=28325 $D=636
M2271 vdd 255 b_pxcb_n<5> vdd hvtpfet l=6e-08 w=2.57e-06 $X=17900 $Y=1941 $D=636
M2272 vdd 256 255 vdd hvtpfet l=6e-08 w=1e-06 $X=17900 $Y=5141 $D=636
M2273 vdd 188 256 vdd hvtpfet l=6e-08 w=6e-07 $X=17900 $Y=8691 $D=636
M2274 vdd 188 257 vdd hvtpfet l=6e-08 w=6e-07 $X=17900 $Y=41842 $D=636
M2275 vdd 257 258 vdd hvtpfet l=6e-08 w=1e-06 $X=17900 $Y=44992 $D=636
M2276 vdd 258 t_pxcb_n<5> vdd hvtpfet l=6e-08 w=2.57e-06 $X=17900 $Y=46622 $D=636
M2277 vdd 260 273 vdd hvtpfet l=6e-08 w=4.11e-07 $X=18106 $Y=14280 $D=636
M2278 1239 wenb 232 vdd hvtpfet l=6e-08 w=8e-07 $X=18366 $Y=35907 $D=636
M2279 1240 tm<4> 648 vdd hvtpfet l=6e-08 w=4.8e-07 $X=18387 $Y=10476 $D=636
M2280 b_pxcb_n<6> 265 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=18410 $Y=1941 $D=636
M2281 265 266 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=18410 $Y=5141 $D=636
M2282 266 253 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=18410 $Y=8691 $D=636
M2283 267 253 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=18410 $Y=41842 $D=636
M2284 268 267 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=18410 $Y=44992 $D=636
M2285 t_pxcb_n<6> 268 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=18410 $Y=46622 $D=636
M2286 1241 ab<4> vdd vdd hvtpfet l=6e-08 w=4.8e-07 $X=18460 $Y=29394 $D=636
M2287 1242 wenb vdd vdd hvtpfet l=6e-08 w=4.8e-07 $X=18460 $Y=33942 $D=636
M2288 vdd tm<2> 173 vdd hvtpfet l=6e-08 w=4.11e-07 $X=18510 $Y=40177 $D=636
M2289 260 ab<1> vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=18616 $Y=14280 $D=636
M2290 vdd 264 1239 vdd hvtpfet l=6e-08 w=8e-07 $X=18626 $Y=35907 $D=636
M2291 1243 33 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=18641 $Y=15520 $D=636
M2292 1244 33 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=18641 $Y=20589 $D=636
M2293 1245 33 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=18641 $Y=22440 $D=636
M2294 1246 33 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=18641 $Y=27509 $D=636
M2295 vdd tm<3> 1240 vdd hvtpfet l=6e-08 w=4.8e-07 $X=18647 $Y=10476 $D=636
M2296 vdd 265 b_pxcb_n<6> vdd hvtpfet l=6e-08 w=2.57e-06 $X=18670 $Y=1941 $D=636
M2297 vdd 266 265 vdd hvtpfet l=6e-08 w=1e-06 $X=18670 $Y=5141 $D=636
M2298 vdd 253 266 vdd hvtpfet l=6e-08 w=6e-07 $X=18670 $Y=8691 $D=636
M2299 vdd 253 267 vdd hvtpfet l=6e-08 w=6e-07 $X=18670 $Y=41842 $D=636
M2300 vdd 267 268 vdd hvtpfet l=6e-08 w=1e-06 $X=18670 $Y=44992 $D=636
M2301 vdd 268 t_pxcb_n<6> vdd hvtpfet l=6e-08 w=2.57e-06 $X=18670 $Y=46622 $D=636
M2302 154 clkb 1241 vdd hvtpfet l=6e-08 w=4.8e-07 $X=18720 $Y=29394 $D=636
M2303 274 clkb 1242 vdd hvtpfet l=6e-08 w=4.8e-07 $X=18720 $Y=33942 $D=636
M2304 280 269 1243 vdd hvtpfet l=6e-08 w=4.11e-07 $X=18911 $Y=15932 $D=636
M2305 281 270 1244 vdd hvtpfet l=6e-08 w=4.11e-07 $X=18911 $Y=20589 $D=636
M2306 282 269 1245 vdd hvtpfet l=6e-08 w=4.11e-07 $X=18911 $Y=22852 $D=636
M2307 283 270 1246 vdd hvtpfet l=6e-08 w=4.11e-07 $X=18911 $Y=27509 $D=636
M2308 655 271 154 vdd hvtpfet l=6e-08 w=3.2e-07 $X=18980 $Y=29554 $D=636
M2309 656 272 274 vdd hvtpfet l=6e-08 w=3.2e-07 $X=18980 $Y=33942 $D=636
M2310 vdd 270 269 vdd hvtpfet l=6e-08 w=4.11e-07 $X=19126 $Y=14280 $D=636
M2311 1247 tm<3> vdd vdd hvtpfet l=6e-08 w=4.8e-07 $X=19157 $Y=10476 $D=636
M2312 1248 273 280 vdd hvtpfet l=6e-08 w=4.11e-07 $X=19171 $Y=15932 $D=636
M2313 1249 273 281 vdd hvtpfet l=6e-08 w=4.11e-07 $X=19171 $Y=20589 $D=636
M2314 1250 260 282 vdd hvtpfet l=6e-08 w=4.11e-07 $X=19171 $Y=22852 $D=636
M2315 1251 260 283 vdd hvtpfet l=6e-08 w=4.11e-07 $X=19171 $Y=27509 $D=636
M2316 b_pxcb_n<7> 275 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=19180 $Y=1941 $D=636
M2317 275 276 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=19180 $Y=5141 $D=636
M2318 276 254 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=19180 $Y=8691 $D=636
M2319 277 254 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=19180 $Y=41842 $D=636
M2320 278 277 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=19180 $Y=44992 $D=636
M2321 t_pxcb_n<7> 278 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=19180 $Y=46622 $D=636
M2322 vdd 23 655 vdd hvtpfet l=6e-08 w=3.2e-07 $X=19240 $Y=29554 $D=636
M2323 vdd 23 656 vdd hvtpfet l=6e-08 w=3.2e-07 $X=19240 $Y=33942 $D=636
M2324 659 243 1247 vdd hvtpfet l=6e-08 w=4.8e-07 $X=19417 $Y=10476 $D=636
M2325 vdd 275 b_pxcb_n<7> vdd hvtpfet l=6e-08 w=2.57e-06 $X=19440 $Y=1941 $D=636
M2326 vdd 276 275 vdd hvtpfet l=6e-08 w=1e-06 $X=19440 $Y=5141 $D=636
M2327 vdd 254 276 vdd hvtpfet l=6e-08 w=6e-07 $X=19440 $Y=8691 $D=636
M2328 vdd 254 277 vdd hvtpfet l=6e-08 w=6e-07 $X=19440 $Y=41842 $D=636
M2329 vdd 277 278 vdd hvtpfet l=6e-08 w=1e-06 $X=19440 $Y=44992 $D=636
M2330 vdd 278 t_pxcb_n<7> vdd hvtpfet l=6e-08 w=2.57e-06 $X=19440 $Y=46622 $D=636
M2331 vdd 33 1248 vdd hvtpfet l=6e-08 w=8.23e-07 $X=19441 $Y=15520 $D=636
M2332 vdd 33 1249 vdd hvtpfet l=6e-08 w=8.23e-07 $X=19441 $Y=20589 $D=636
M2333 vdd 33 1250 vdd hvtpfet l=6e-08 w=8.23e-07 $X=19441 $Y=22440 $D=636
M2334 vdd 33 1251 vdd hvtpfet l=6e-08 w=8.23e-07 $X=19441 $Y=27509 $D=636
M2335 271 154 vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=19500 $Y=29554 $D=636
M2336 272 274 vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=19500 $Y=33942 $D=636
M2337 270 ab<0> vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=19636 $Y=14280 $D=636
M2338 vdd 15 r_saeb_n vdd hvtpfet l=6e-08 w=1.43e-06 $X=19675 $Y=35277 $D=636
M2339 r_saeb_n 15 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=19935 $Y=35277 $D=636
M2340 212 280 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=19951 $Y=15321 $D=636
M2341 1252 43 280 vdd hvtpfet l=6e-08 w=2.74e-07 $X=19951 $Y=16069 $D=636
M2342 1253 43 281 vdd hvtpfet l=6e-08 w=2.74e-07 $X=19951 $Y=20589 $D=636
M2343 185 281 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=19951 $Y=21405 $D=636
M2344 155 282 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=19951 $Y=22241 $D=636
M2345 1254 43 282 vdd hvtpfet l=6e-08 w=2.74e-07 $X=19951 $Y=22989 $D=636
M2346 1255 43 283 vdd hvtpfet l=6e-08 w=2.74e-07 $X=19951 $Y=27509 $D=636
M2347 145 283 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=19951 $Y=28325 $D=636
M2348 vdd 11 rb_cb<0> vdd hvtpfet l=6e-08 w=1.43e-06 $X=20195 $Y=1506 $D=636
M2349 vdd 12 rb_cb<2> vdd hvtpfet l=6e-08 w=1.43e-06 $X=20195 $Y=3566 $D=636
M2350 vdd 13 rb_mb<0> vdd hvtpfet l=6e-08 w=1.43e-06 $X=20195 $Y=7966 $D=636
M2351 vdd 14 rb_mb<2> vdd hvtpfet l=6e-08 w=1.43e-06 $X=20195 $Y=10026 $D=636
M2352 vdd 15 r_saeb_n vdd hvtpfet l=6e-08 w=1.43e-06 $X=20195 $Y=35277 $D=636
M2353 vdd 16 rt_mb<2> vdd hvtpfet l=6e-08 w=1.43e-06 $X=20195 $Y=39677 $D=636
M2354 vdd 17 rt_mb<0> vdd hvtpfet l=6e-08 w=1.43e-06 $X=20195 $Y=41737 $D=636
M2355 vdd 18 rt_cb<2> vdd hvtpfet l=6e-08 w=1.43e-06 $X=20195 $Y=46137 $D=636
M2356 vdd 19 rt_cb<0> vdd hvtpfet l=6e-08 w=1.43e-06 $X=20195 $Y=48197 $D=636
M2357 vdd 280 212 vdd hvtpfet l=6e-08 w=2.06e-07 $X=20211 $Y=15321 $D=636
M2358 vdd 212 1252 vdd hvtpfet l=6e-08 w=2.74e-07 $X=20211 $Y=16069 $D=636
M2359 vdd 185 1253 vdd hvtpfet l=6e-08 w=2.74e-07 $X=20211 $Y=20589 $D=636
M2360 vdd 281 185 vdd hvtpfet l=6e-08 w=2.06e-07 $X=20211 $Y=21405 $D=636
M2361 vdd 282 155 vdd hvtpfet l=6e-08 w=2.06e-07 $X=20211 $Y=22241 $D=636
M2362 vdd 155 1254 vdd hvtpfet l=6e-08 w=2.74e-07 $X=20211 $Y=22989 $D=636
M2363 vdd 145 1255 vdd hvtpfet l=6e-08 w=2.74e-07 $X=20211 $Y=27509 $D=636
M2364 vdd 283 145 vdd hvtpfet l=6e-08 w=2.06e-07 $X=20211 $Y=28325 $D=636
M2365 rb_cb<0> 11 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=20455 $Y=1506 $D=636
M2366 rb_cb<2> 12 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=20455 $Y=3566 $D=636
M2367 rb_mb<0> 13 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=20455 $Y=7966 $D=636
M2368 rb_mb<2> 14 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=20455 $Y=10026 $D=636
M2369 r_saeb_n 15 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=20455 $Y=35277 $D=636
M2370 rt_mb<2> 16 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=20455 $Y=39677 $D=636
M2371 rt_mb<0> 17 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=20455 $Y=41737 $D=636
M2372 rt_cb<2> 18 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=20455 $Y=46137 $D=636
M2373 rt_cb<0> 19 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=20455 $Y=48197 $D=636
M2374 vdd 11 rb_cb<0> vdd hvtpfet l=6e-08 w=1.43e-06 $X=20715 $Y=1506 $D=636
M2375 vdd 12 rb_cb<2> vdd hvtpfet l=6e-08 w=1.43e-06 $X=20715 $Y=3566 $D=636
M2376 vdd 13 rb_mb<0> vdd hvtpfet l=6e-08 w=1.43e-06 $X=20715 $Y=7966 $D=636
M2377 vdd 14 rb_mb<2> vdd hvtpfet l=6e-08 w=1.43e-06 $X=20715 $Y=10026 $D=636
M2378 vdd 15 r_saeb_n vdd hvtpfet l=6e-08 w=1.43e-06 $X=20715 $Y=35277 $D=636
M2379 vdd 16 rt_mb<2> vdd hvtpfet l=6e-08 w=1.43e-06 $X=20715 $Y=39677 $D=636
M2380 vdd 17 rt_mb<0> vdd hvtpfet l=6e-08 w=1.43e-06 $X=20715 $Y=41737 $D=636
M2381 vdd 18 rt_cb<2> vdd hvtpfet l=6e-08 w=1.43e-06 $X=20715 $Y=46137 $D=636
M2382 vdd 19 rt_cb<0> vdd hvtpfet l=6e-08 w=1.43e-06 $X=20715 $Y=48197 $D=636
M2383 10 274 vdd vdd hvtpfet l=6e-08 w=1.2e-06 $X=20725 $Y=32684 $D=636
M2384 rb_cb<1> 34 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=20975 $Y=1506 $D=636
M2385 rb_cb<3> 35 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=20975 $Y=3566 $D=636
M2386 rb_mb<1> 36 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=20975 $Y=7966 $D=636
M2387 rb_mb<3> 37 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=20975 $Y=10026 $D=636
M2388 r_clk_dqb 8 vdd vdd hvtpfet l=6e-08 w=2.1e-06 $X=20975 $Y=23696 $D=636
M2389 r_clk_dqb_n 9 vdd vdd hvtpfet l=6e-08 w=2.1e-06 $X=20975 $Y=26512 $D=636
M2390 r_sa_preb_n 51 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=20975 $Y=35277 $D=636
M2391 rt_mb<3> 39 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=20975 $Y=39677 $D=636
M2392 rt_mb<1> 40 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=20975 $Y=41737 $D=636
M2393 rt_cb<3> 41 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=20975 $Y=46137 $D=636
M2394 rt_cb<1> 42 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=20975 $Y=48197 $D=636
M2395 vdd 34 rb_cb<1> vdd hvtpfet l=6e-08 w=1.43e-06 $X=21235 $Y=1506 $D=636
M2396 vdd 35 rb_cb<3> vdd hvtpfet l=6e-08 w=1.43e-06 $X=21235 $Y=3566 $D=636
M2397 vdd 36 rb_mb<1> vdd hvtpfet l=6e-08 w=1.43e-06 $X=21235 $Y=7966 $D=636
M2398 vdd 37 rb_mb<3> vdd hvtpfet l=6e-08 w=1.43e-06 $X=21235 $Y=10026 $D=636
M2399 rb_tm_preb_n 20 vdd vdd hvtpfet l=6e-08 w=2.145e-06 $X=21235 $Y=14887 $D=636
M2400 rt_tm_preb_n 21 vdd vdd hvtpfet l=6e-08 w=2.145e-06 $X=21235 $Y=17659 $D=636
M2401 vdd 8 r_clk_dqb vdd hvtpfet l=6e-08 w=2.1e-06 $X=21235 $Y=23696 $D=636
M2402 vdd 9 r_clk_dqb_n vdd hvtpfet l=6e-08 w=2.1e-06 $X=21235 $Y=26512 $D=636
M2403 r_lweb 10 vdd vdd hvtpfet l=6e-08 w=2.145e-06 $X=21235 $Y=32504 $D=636
M2404 vdd 51 r_sa_preb_n vdd hvtpfet l=6e-08 w=1.43e-06 $X=21235 $Y=35277 $D=636
M2405 vdd 39 rt_mb<3> vdd hvtpfet l=6e-08 w=1.43e-06 $X=21235 $Y=39677 $D=636
M2406 vdd 40 rt_mb<1> vdd hvtpfet l=6e-08 w=1.43e-06 $X=21235 $Y=41737 $D=636
M2407 vdd 41 rt_cb<3> vdd hvtpfet l=6e-08 w=1.43e-06 $X=21235 $Y=46137 $D=636
M2408 vdd 42 rt_cb<1> vdd hvtpfet l=6e-08 w=1.43e-06 $X=21235 $Y=48197 $D=636
M2409 rb_cb<1> 34 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=21495 $Y=1506 $D=636
M2410 rb_cb<3> 35 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=21495 $Y=3566 $D=636
M2411 rb_mb<1> 36 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=21495 $Y=7966 $D=636
M2412 rb_mb<3> 37 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=21495 $Y=10026 $D=636
M2413 vdd 20 rb_tm_preb_n vdd hvtpfet l=6e-08 w=2.145e-06 $X=21495 $Y=14887 $D=636
M2414 vdd 21 rt_tm_preb_n vdd hvtpfet l=6e-08 w=2.145e-06 $X=21495 $Y=17659 $D=636
M2415 r_clk_dqb 8 vdd vdd hvtpfet l=6e-08 w=2.1e-06 $X=21495 $Y=23696 $D=636
M2416 r_clk_dqb_n 9 vdd vdd hvtpfet l=6e-08 w=2.1e-06 $X=21495 $Y=26512 $D=636
M2417 vdd 10 r_lweb vdd hvtpfet l=6e-08 w=2.145e-06 $X=21495 $Y=32504 $D=636
M2418 r_sa_preb_n 51 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=21495 $Y=35277 $D=636
M2419 rt_mb<3> 39 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=21495 $Y=39677 $D=636
M2420 rt_mb<1> 40 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=21495 $Y=41737 $D=636
M2421 rt_cb<3> 41 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=21495 $Y=46137 $D=636
M2422 rt_cb<1> 42 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=21495 $Y=48197 $D=636
M2423 vdd 289 lb_ca<1> vdd hvtpfet l=6e-08 w=1.43e-06 $X=22005 $Y=1506 $D=636
M2424 vdd 290 lb_ca<3> vdd hvtpfet l=6e-08 w=1.43e-06 $X=22005 $Y=3566 $D=636
M2425 vdd 291 lb_ma<1> vdd hvtpfet l=6e-08 w=1.43e-06 $X=22005 $Y=7966 $D=636
M2426 vdd 292 lb_ma<3> vdd hvtpfet l=6e-08 w=1.43e-06 $X=22005 $Y=10026 $D=636
M2427 lb_tm_prea_n 285 vdd vdd hvtpfet l=6e-08 w=2.145e-06 $X=22005 $Y=14887 $D=636
M2428 lt_tm_prea_n 286 vdd vdd hvtpfet l=6e-08 w=2.145e-06 $X=22005 $Y=17659 $D=636
M2429 vdd 287 l_clk_dqa vdd hvtpfet l=6e-08 w=2.1e-06 $X=22005 $Y=23696 $D=636
M2430 vdd 288 l_clk_dqa_n vdd hvtpfet l=6e-08 w=2.1e-06 $X=22005 $Y=26512 $D=636
M2431 l_lwea 284 vdd vdd hvtpfet l=6e-08 w=2.145e-06 $X=22005 $Y=32504 $D=636
M2432 vdd 293 l_sa_prea_n vdd hvtpfet l=6e-08 w=1.43e-06 $X=22005 $Y=35277 $D=636
M2433 vdd 294 lt_ma<3> vdd hvtpfet l=6e-08 w=1.43e-06 $X=22005 $Y=39677 $D=636
M2434 vdd 295 lt_ma<1> vdd hvtpfet l=6e-08 w=1.43e-06 $X=22005 $Y=41737 $D=636
M2435 vdd 296 lt_ca<3> vdd hvtpfet l=6e-08 w=1.43e-06 $X=22005 $Y=46137 $D=636
M2436 vdd 297 lt_ca<1> vdd hvtpfet l=6e-08 w=1.43e-06 $X=22005 $Y=48197 $D=636
M2437 lb_ca<1> 289 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=22265 $Y=1506 $D=636
M2438 lb_ca<3> 290 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=22265 $Y=3566 $D=636
M2439 lb_ma<1> 291 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=22265 $Y=7966 $D=636
M2440 lb_ma<3> 292 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=22265 $Y=10026 $D=636
M2441 vdd 285 lb_tm_prea_n vdd hvtpfet l=6e-08 w=2.145e-06 $X=22265 $Y=14887 $D=636
M2442 vdd 286 lt_tm_prea_n vdd hvtpfet l=6e-08 w=2.145e-06 $X=22265 $Y=17659 $D=636
M2443 l_clk_dqa 287 vdd vdd hvtpfet l=6e-08 w=2.1e-06 $X=22265 $Y=23696 $D=636
M2444 l_clk_dqa_n 288 vdd vdd hvtpfet l=6e-08 w=2.1e-06 $X=22265 $Y=26512 $D=636
M2445 vdd 284 l_lwea vdd hvtpfet l=6e-08 w=2.145e-06 $X=22265 $Y=32504 $D=636
M2446 l_sa_prea_n 293 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=22265 $Y=35277 $D=636
M2447 lt_ma<3> 294 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=22265 $Y=39677 $D=636
M2448 lt_ma<1> 295 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=22265 $Y=41737 $D=636
M2449 lt_ca<3> 296 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=22265 $Y=46137 $D=636
M2450 lt_ca<1> 297 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=22265 $Y=48197 $D=636
M2451 vdd 289 lb_ca<1> vdd hvtpfet l=6e-08 w=1.43e-06 $X=22525 $Y=1506 $D=636
M2452 vdd 290 lb_ca<3> vdd hvtpfet l=6e-08 w=1.43e-06 $X=22525 $Y=3566 $D=636
M2453 vdd 291 lb_ma<1> vdd hvtpfet l=6e-08 w=1.43e-06 $X=22525 $Y=7966 $D=636
M2454 vdd 292 lb_ma<3> vdd hvtpfet l=6e-08 w=1.43e-06 $X=22525 $Y=10026 $D=636
M2455 vdd 287 l_clk_dqa vdd hvtpfet l=6e-08 w=2.1e-06 $X=22525 $Y=23696 $D=636
M2456 vdd 288 l_clk_dqa_n vdd hvtpfet l=6e-08 w=2.1e-06 $X=22525 $Y=26512 $D=636
M2457 vdd 293 l_sa_prea_n vdd hvtpfet l=6e-08 w=1.43e-06 $X=22525 $Y=35277 $D=636
M2458 vdd 294 lt_ma<3> vdd hvtpfet l=6e-08 w=1.43e-06 $X=22525 $Y=39677 $D=636
M2459 vdd 295 lt_ma<1> vdd hvtpfet l=6e-08 w=1.43e-06 $X=22525 $Y=41737 $D=636
M2460 vdd 296 lt_ca<3> vdd hvtpfet l=6e-08 w=1.43e-06 $X=22525 $Y=46137 $D=636
M2461 vdd 297 lt_ca<1> vdd hvtpfet l=6e-08 w=1.43e-06 $X=22525 $Y=48197 $D=636
M2462 vdd 298 284 vdd hvtpfet l=6e-08 w=1.2e-06 $X=22775 $Y=32684 $D=636
M2463 lb_ca<0> 299 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=22785 $Y=1506 $D=636
M2464 lb_ca<2> 300 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=22785 $Y=3566 $D=636
M2465 lb_ma<0> 301 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=22785 $Y=7966 $D=636
M2466 lb_ma<2> 302 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=22785 $Y=10026 $D=636
M2467 l_saea_n 303 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=22785 $Y=35277 $D=636
M2468 lt_ma<2> 304 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=22785 $Y=39677 $D=636
M2469 lt_ma<0> 305 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=22785 $Y=41737 $D=636
M2470 lt_ca<2> 306 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=22785 $Y=46137 $D=636
M2471 lt_ca<0> 307 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=22785 $Y=48197 $D=636
M2472 vdd 299 lb_ca<0> vdd hvtpfet l=6e-08 w=1.43e-06 $X=23045 $Y=1506 $D=636
M2473 vdd 300 lb_ca<2> vdd hvtpfet l=6e-08 w=1.43e-06 $X=23045 $Y=3566 $D=636
M2474 vdd 301 lb_ma<0> vdd hvtpfet l=6e-08 w=1.43e-06 $X=23045 $Y=7966 $D=636
M2475 vdd 302 lb_ma<2> vdd hvtpfet l=6e-08 w=1.43e-06 $X=23045 $Y=10026 $D=636
M2476 vdd 303 l_saea_n vdd hvtpfet l=6e-08 w=1.43e-06 $X=23045 $Y=35277 $D=636
M2477 vdd 304 lt_ma<2> vdd hvtpfet l=6e-08 w=1.43e-06 $X=23045 $Y=39677 $D=636
M2478 vdd 305 lt_ma<0> vdd hvtpfet l=6e-08 w=1.43e-06 $X=23045 $Y=41737 $D=636
M2479 vdd 306 lt_ca<2> vdd hvtpfet l=6e-08 w=1.43e-06 $X=23045 $Y=46137 $D=636
M2480 vdd 307 lt_ca<0> vdd hvtpfet l=6e-08 w=1.43e-06 $X=23045 $Y=48197 $D=636
M2481 308 312 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=23289 $Y=15321 $D=636
M2482 1256 308 vdd vdd hvtpfet l=6e-08 w=2.74e-07 $X=23289 $Y=16069 $D=636
M2483 1257 309 vdd vdd hvtpfet l=6e-08 w=2.74e-07 $X=23289 $Y=20589 $D=636
M2484 309 313 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=23289 $Y=21405 $D=636
M2485 310 314 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=23289 $Y=22241 $D=636
M2486 1258 310 vdd vdd hvtpfet l=6e-08 w=2.74e-07 $X=23289 $Y=22989 $D=636
M2487 1259 311 vdd vdd hvtpfet l=6e-08 w=2.74e-07 $X=23289 $Y=27509 $D=636
M2488 311 315 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=23289 $Y=28325 $D=636
M2489 lb_ca<0> 299 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=23305 $Y=1506 $D=636
M2490 lb_ca<2> 300 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=23305 $Y=3566 $D=636
M2491 lb_ma<0> 301 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=23305 $Y=7966 $D=636
M2492 lb_ma<2> 302 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=23305 $Y=10026 $D=636
M2493 l_saea_n 303 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=23305 $Y=35277 $D=636
M2494 lt_ma<2> 304 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=23305 $Y=39677 $D=636
M2495 lt_ma<0> 305 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=23305 $Y=41737 $D=636
M2496 lt_ca<2> 306 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=23305 $Y=46137 $D=636
M2497 lt_ca<0> 307 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=23305 $Y=48197 $D=636
M2498 vdd 312 308 vdd hvtpfet l=6e-08 w=2.06e-07 $X=23549 $Y=15321 $D=636
M2499 312 323 1256 vdd hvtpfet l=6e-08 w=2.74e-07 $X=23549 $Y=16069 $D=636
M2500 313 323 1257 vdd hvtpfet l=6e-08 w=2.74e-07 $X=23549 $Y=20589 $D=636
M2501 vdd 313 309 vdd hvtpfet l=6e-08 w=2.06e-07 $X=23549 $Y=21405 $D=636
M2502 vdd 314 310 vdd hvtpfet l=6e-08 w=2.06e-07 $X=23549 $Y=22241 $D=636
M2503 314 323 1258 vdd hvtpfet l=6e-08 w=2.74e-07 $X=23549 $Y=22989 $D=636
M2504 315 323 1259 vdd hvtpfet l=6e-08 w=2.74e-07 $X=23549 $Y=27509 $D=636
M2505 vdd 315 311 vdd hvtpfet l=6e-08 w=2.06e-07 $X=23549 $Y=28325 $D=636
M2506 vdd 303 l_saea_n vdd hvtpfet l=6e-08 w=1.43e-06 $X=23565 $Y=35277 $D=636
M2507 l_saea_n 303 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=23825 $Y=35277 $D=636
M2508 vdd aa<0> 327 vdd hvtpfet l=6e-08 w=4.11e-07 $X=23864 $Y=14280 $D=636
M2509 vdd 324 331 vdd hvtpfet l=6e-08 w=3.2e-07 $X=24000 $Y=29554 $D=636
M2510 vdd 298 332 vdd hvtpfet l=6e-08 w=3.2e-07 $X=24000 $Y=33942 $D=636
M2511 1261 317 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=24059 $Y=15520 $D=636
M2512 1262 317 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=24059 $Y=20589 $D=636
M2513 1263 317 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=24059 $Y=22440 $D=636
M2514 1264 317 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=24059 $Y=27509 $D=636
M2515 b_pxca_n<7> 318 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=24060 $Y=1941 $D=636
M2516 318 319 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=24060 $Y=5141 $D=636
M2517 319 320 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=24060 $Y=8691 $D=636
M2518 321 320 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=24060 $Y=41842 $D=636
M2519 322 321 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=24060 $Y=44992 $D=636
M2520 t_pxca_n<7> 322 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=24060 $Y=46622 $D=636
M2521 1260 325 709 vdd hvtpfet l=6e-08 w=4.8e-07 $X=24083 $Y=10476 $D=636
M2522 712 340 vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=24260 $Y=29554 $D=636
M2523 713 340 vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=24260 $Y=33942 $D=636
M2524 vdd 318 b_pxca_n<7> vdd hvtpfet l=6e-08 w=2.57e-06 $X=24320 $Y=1941 $D=636
M2525 vdd 319 318 vdd hvtpfet l=6e-08 w=1e-06 $X=24320 $Y=5141 $D=636
M2526 vdd 320 319 vdd hvtpfet l=6e-08 w=6e-07 $X=24320 $Y=8691 $D=636
M2527 vdd 320 321 vdd hvtpfet l=6e-08 w=6e-07 $X=24320 $Y=41842 $D=636
M2528 vdd 321 322 vdd hvtpfet l=6e-08 w=1e-06 $X=24320 $Y=44992 $D=636
M2529 vdd 322 t_pxca_n<7> vdd hvtpfet l=6e-08 w=2.57e-06 $X=24320 $Y=46622 $D=636
M2530 312 328 1261 vdd hvtpfet l=6e-08 w=4.11e-07 $X=24329 $Y=15932 $D=636
M2531 313 328 1262 vdd hvtpfet l=6e-08 w=4.11e-07 $X=24329 $Y=20589 $D=636
M2532 314 329 1263 vdd hvtpfet l=6e-08 w=4.11e-07 $X=24329 $Y=22852 $D=636
M2533 315 329 1264 vdd hvtpfet l=6e-08 w=4.11e-07 $X=24329 $Y=27509 $D=636
M2534 vdd tm<8> 1260 vdd hvtpfet l=6e-08 w=4.8e-07 $X=24343 $Y=10476 $D=636
M2535 334 327 vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=24374 $Y=14280 $D=636
M2536 vdd tm<5> 264 vdd hvtpfet l=6e-08 w=4.11e-07 $X=24518 $Y=40177 $D=636
M2537 324 331 712 vdd hvtpfet l=6e-08 w=3.2e-07 $X=24520 $Y=29554 $D=636
M2538 298 332 713 vdd hvtpfet l=6e-08 w=3.2e-07 $X=24520 $Y=33942 $D=636
M2539 1265 334 312 vdd hvtpfet l=6e-08 w=4.11e-07 $X=24589 $Y=15932 $D=636
M2540 1266 327 313 vdd hvtpfet l=6e-08 w=4.11e-07 $X=24589 $Y=20589 $D=636
M2541 1267 334 314 vdd hvtpfet l=6e-08 w=4.11e-07 $X=24589 $Y=22852 $D=636
M2542 1268 327 315 vdd hvtpfet l=6e-08 w=4.11e-07 $X=24589 $Y=27509 $D=636
M2543 1269 clka 324 vdd hvtpfet l=6e-08 w=4.8e-07 $X=24780 $Y=29394 $D=636
M2544 1270 clka 298 vdd hvtpfet l=6e-08 w=4.8e-07 $X=24780 $Y=33942 $D=636
M2545 b_pxca_n<6> 335 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=24830 $Y=1941 $D=636
M2546 335 336 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=24830 $Y=5141 $D=636
M2547 336 337 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=24830 $Y=8691 $D=636
M2548 338 337 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=24830 $Y=41842 $D=636
M2549 339 338 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=24830 $Y=44992 $D=636
M2550 t_pxca_n<6> 339 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=24830 $Y=46622 $D=636
M2551 1271 tm<8> vdd vdd hvtpfet l=6e-08 w=4.8e-07 $X=24853 $Y=10476 $D=636
M2552 vdd 317 1265 vdd hvtpfet l=6e-08 w=8.23e-07 $X=24859 $Y=15520 $D=636
M2553 vdd 317 1266 vdd hvtpfet l=6e-08 w=8.23e-07 $X=24859 $Y=20589 $D=636
M2554 vdd 317 1267 vdd hvtpfet l=6e-08 w=8.23e-07 $X=24859 $Y=22440 $D=636
M2555 vdd 317 1268 vdd hvtpfet l=6e-08 w=8.23e-07 $X=24859 $Y=27509 $D=636
M2556 1272 264 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=24874 $Y=35907 $D=636
M2557 vdd aa<1> 329 vdd hvtpfet l=6e-08 w=4.11e-07 $X=24884 $Y=14280 $D=636
M2558 vdd aa<4> 1269 vdd hvtpfet l=6e-08 w=4.8e-07 $X=25040 $Y=29394 $D=636
M2559 vdd wena 1270 vdd hvtpfet l=6e-08 w=4.8e-07 $X=25040 $Y=33942 $D=636
M2560 vdd 335 b_pxca_n<6> vdd hvtpfet l=6e-08 w=2.57e-06 $X=25090 $Y=1941 $D=636
M2561 vdd 336 335 vdd hvtpfet l=6e-08 w=1e-06 $X=25090 $Y=5141 $D=636
M2562 vdd 337 336 vdd hvtpfet l=6e-08 w=6e-07 $X=25090 $Y=8691 $D=636
M2563 vdd 337 338 vdd hvtpfet l=6e-08 w=6e-07 $X=25090 $Y=41842 $D=636
M2564 vdd 338 339 vdd hvtpfet l=6e-08 w=1e-06 $X=25090 $Y=44992 $D=636
M2565 vdd 339 t_pxca_n<6> vdd hvtpfet l=6e-08 w=2.57e-06 $X=25090 $Y=46622 $D=636
M2566 718 tm<9> 1271 vdd hvtpfet l=6e-08 w=4.8e-07 $X=25113 $Y=10476 $D=636
M2567 376 wena 1272 vdd hvtpfet l=6e-08 w=8e-07 $X=25134 $Y=35907 $D=636
M2568 328 329 vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=25394 $Y=14280 $D=636
M2569 b_pxca_n<5> 345 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=25600 $Y=1941 $D=636
M2570 345 346 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=25600 $Y=5141 $D=636
M2571 346 347 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=25600 $Y=8691 $D=636
M2572 348 347 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=25600 $Y=41842 $D=636
M2573 349 348 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=25600 $Y=44992 $D=636
M2574 t_pxca_n<5> 349 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=25600 $Y=46622 $D=636
M2575 337 352 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=25609 $Y=15321 $D=636
M2576 1273 337 vdd vdd hvtpfet l=6e-08 w=2.74e-07 $X=25609 $Y=16069 $D=636
M2577 1274 320 vdd vdd hvtpfet l=6e-08 w=2.74e-07 $X=25609 $Y=20589 $D=636
M2578 320 353 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=25609 $Y=21405 $D=636
M2579 350 354 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=25609 $Y=22241 $D=636
M2580 1275 350 vdd vdd hvtpfet l=6e-08 w=2.74e-07 $X=25609 $Y=22989 $D=636
M2581 1276 351 vdd vdd hvtpfet l=6e-08 w=2.74e-07 $X=25609 $Y=27509 $D=636
M2582 351 355 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=25609 $Y=28325 $D=636
M2583 1277 tm<9> 721 vdd hvtpfet l=6e-08 w=4.8e-07 $X=25623 $Y=10476 $D=636
M2584 vdd clka 340 vdd hvtpfet l=6e-08 w=9e-07 $X=25854 $Y=29274 $D=636
M2585 vdd 345 b_pxca_n<5> vdd hvtpfet l=6e-08 w=2.57e-06 $X=25860 $Y=1941 $D=636
M2586 vdd 346 345 vdd hvtpfet l=6e-08 w=1e-06 $X=25860 $Y=5141 $D=636
M2587 vdd 347 346 vdd hvtpfet l=6e-08 w=6e-07 $X=25860 $Y=8691 $D=636
M2588 vdd 347 348 vdd hvtpfet l=6e-08 w=6e-07 $X=25860 $Y=41842 $D=636
M2589 vdd 348 349 vdd hvtpfet l=6e-08 w=1e-06 $X=25860 $Y=44992 $D=636
M2590 vdd 349 t_pxca_n<5> vdd hvtpfet l=6e-08 w=2.57e-06 $X=25860 $Y=46622 $D=636
M2591 vdd 352 337 vdd hvtpfet l=6e-08 w=2.06e-07 $X=25869 $Y=15321 $D=636
M2592 352 323 1273 vdd hvtpfet l=6e-08 w=2.74e-07 $X=25869 $Y=16069 $D=636
M2593 353 323 1274 vdd hvtpfet l=6e-08 w=2.74e-07 $X=25869 $Y=20589 $D=636
M2594 vdd 353 320 vdd hvtpfet l=6e-08 w=2.06e-07 $X=25869 $Y=21405 $D=636
M2595 vdd 354 350 vdd hvtpfet l=6e-08 w=2.06e-07 $X=25869 $Y=22241 $D=636
M2596 354 323 1275 vdd hvtpfet l=6e-08 w=2.74e-07 $X=25869 $Y=22989 $D=636
M2597 355 323 1276 vdd hvtpfet l=6e-08 w=2.74e-07 $X=25869 $Y=27509 $D=636
M2598 vdd 355 351 vdd hvtpfet l=6e-08 w=2.06e-07 $X=25869 $Y=28325 $D=636
M2599 vdd 366 1277 vdd hvtpfet l=6e-08 w=4.8e-07 $X=25883 $Y=10476 $D=636
M2600 vdd 356 363 vdd hvtpfet l=6e-08 w=3.2e-07 $X=26138 $Y=35913 $D=636
M2601 b_pxca_n<4> 357 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=26370 $Y=1941 $D=636
M2602 357 358 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=26370 $Y=5141 $D=636
M2603 358 359 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=26370 $Y=8691 $D=636
M2604 360 359 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=26370 $Y=41842 $D=636
M2605 361 360 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=26370 $Y=44992 $D=636
M2606 t_pxca_n<4> 361 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=26370 $Y=46622 $D=636
M2607 729 123 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=26374 $Y=29274 $D=636
M2608 1279 317 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=26379 $Y=15520 $D=636
M2609 1280 317 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=26379 $Y=20589 $D=636
M2610 1281 317 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=26379 $Y=22440 $D=636
M2611 1282 317 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=26379 $Y=27509 $D=636
M2612 1278 366 vdd vdd hvtpfet l=6e-08 w=4.8e-07 $X=26393 $Y=10476 $D=636
M2613 725 368 vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=26398 $Y=35913 $D=636
M2614 vdd 357 b_pxca_n<4> vdd hvtpfet l=6e-08 w=2.57e-06 $X=26630 $Y=1941 $D=636
M2615 vdd 358 357 vdd hvtpfet l=6e-08 w=1e-06 $X=26630 $Y=5141 $D=636
M2616 vdd 359 358 vdd hvtpfet l=6e-08 w=6e-07 $X=26630 $Y=8691 $D=636
M2617 vdd 359 360 vdd hvtpfet l=6e-08 w=6e-07 $X=26630 $Y=41842 $D=636
M2618 vdd 360 361 vdd hvtpfet l=6e-08 w=1e-06 $X=26630 $Y=44992 $D=636
M2619 vdd 361 t_pxca_n<4> vdd hvtpfet l=6e-08 w=2.57e-06 $X=26630 $Y=46622 $D=636
M2620 vdd 123 729 vdd hvtpfet l=6e-08 w=6e-07 $X=26634 $Y=29274 $D=636
M2621 352 364 1279 vdd hvtpfet l=6e-08 w=4.11e-07 $X=26649 $Y=15932 $D=636
M2622 353 364 1280 vdd hvtpfet l=6e-08 w=4.11e-07 $X=26649 $Y=20589 $D=636
M2623 354 365 1281 vdd hvtpfet l=6e-08 w=4.11e-07 $X=26649 $Y=22852 $D=636
M2624 355 365 1282 vdd hvtpfet l=6e-08 w=4.11e-07 $X=26649 $Y=27509 $D=636
M2625 727 325 1278 vdd hvtpfet l=6e-08 w=4.8e-07 $X=26653 $Y=10476 $D=636
M2626 356 363 725 vdd hvtpfet l=6e-08 w=3.2e-07 $X=26658 $Y=35913 $D=636
M2627 vdd tm<7> 726 vdd hvtpfet l=6e-08 w=4.11e-07 $X=26820 $Y=40177 $D=636
M2628 1283 123 vdd vdd hvtpfet l=6e-08 w=4.8e-07 $X=26839 $Y=33942 $D=636
M2629 729 123 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=26894 $Y=29274 $D=636
M2630 1285 369 352 vdd hvtpfet l=6e-08 w=4.11e-07 $X=26909 $Y=15932 $D=636
M2631 1286 369 353 vdd hvtpfet l=6e-08 w=4.11e-07 $X=26909 $Y=20589 $D=636
M2632 1287 369 354 vdd hvtpfet l=6e-08 w=4.11e-07 $X=26909 $Y=22852 $D=636
M2633 1288 369 355 vdd hvtpfet l=6e-08 w=4.11e-07 $X=26909 $Y=27509 $D=636
M2634 1284 362 356 vdd hvtpfet l=6e-08 w=4.8e-07 $X=26918 $Y=35753 $D=636
M2635 vdd aa<10> 374 vdd hvtpfet l=6e-08 w=4.11e-07 $X=26924 $Y=14280 $D=636
M2636 379 131 1283 vdd hvtpfet l=6e-08 w=4.8e-07 $X=27099 $Y=33942 $D=636
M2637 b_pxca_n<3> 370 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=27140 $Y=1941 $D=636
M2638 370 371 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=27140 $Y=5141 $D=636
M2639 371 351 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=27140 $Y=8691 $D=636
M2640 372 351 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=27140 $Y=41842 $D=636
M2641 373 372 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=27140 $Y=44992 $D=636
M2642 t_pxca_n<3> 373 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=27140 $Y=46622 $D=636
M2643 vdd 123 729 vdd hvtpfet l=6e-08 w=6e-07 $X=27154 $Y=29274 $D=636
M2644 vdd tm<9> 325 vdd hvtpfet l=7e-08 w=4.8e-07 $X=27163 $Y=10476 $D=636
M2645 vdd 376 1284 vdd hvtpfet l=6e-08 w=4.8e-07 $X=27178 $Y=35753 $D=636
M2646 vdd 317 1285 vdd hvtpfet l=6e-08 w=8.23e-07 $X=27179 $Y=15520 $D=636
M2647 vdd 317 1286 vdd hvtpfet l=6e-08 w=8.23e-07 $X=27179 $Y=20589 $D=636
M2648 vdd 317 1287 vdd hvtpfet l=6e-08 w=8.23e-07 $X=27179 $Y=22440 $D=636
M2649 vdd 317 1288 vdd hvtpfet l=6e-08 w=8.23e-07 $X=27179 $Y=27509 $D=636
M2650 375 374 vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=27184 $Y=14280 $D=636
M2651 736 377 379 vdd hvtpfet l=6e-08 w=3.2e-07 $X=27359 $Y=33942 $D=636
M2652 vdd 370 b_pxca_n<3> vdd hvtpfet l=6e-08 w=2.57e-06 $X=27400 $Y=1941 $D=636
M2653 vdd 371 370 vdd hvtpfet l=6e-08 w=1e-06 $X=27400 $Y=5141 $D=636
M2654 vdd 351 371 vdd hvtpfet l=6e-08 w=6e-07 $X=27400 $Y=8691 $D=636
M2655 vdd 351 372 vdd hvtpfet l=6e-08 w=6e-07 $X=27400 $Y=41842 $D=636
M2656 vdd 372 373 vdd hvtpfet l=6e-08 w=1e-06 $X=27400 $Y=44992 $D=636
M2657 vdd 373 t_pxca_n<3> vdd hvtpfet l=6e-08 w=2.57e-06 $X=27400 $Y=46622 $D=636
M2658 366 tm<8> vdd vdd hvtpfet l=7e-08 w=4.8e-07 $X=27433 $Y=10476 $D=636
M2659 vdd 123 736 vdd hvtpfet l=6e-08 w=3.2e-07 $X=27619 $Y=33942 $D=636
M2660 vdd tm<1> 735 vdd hvtpfet l=6e-08 w=4.11e-07 $X=27620 $Y=40177 $D=636
M2661 317 323 vdd vdd hvtpfet l=6e-08 w=7e-07 $X=27664 $Y=29648 $D=636
M2662 1289 374 352 vdd hvtpfet l=6e-08 w=4.11e-07 $X=27689 $Y=15932 $D=636
M2663 1290 375 353 vdd hvtpfet l=6e-08 w=4.11e-07 $X=27689 $Y=20589 $D=636
M2664 1291 374 354 vdd hvtpfet l=6e-08 w=4.11e-07 $X=27689 $Y=22852 $D=636
M2665 1292 375 355 vdd hvtpfet l=6e-08 w=4.11e-07 $X=27689 $Y=27509 $D=636
M2666 vdd 380 369 vdd hvtpfet l=6e-08 w=4.11e-07 $X=27784 $Y=14280 $D=636
M2667 vdd 362 386 vdd hvtpfet l=6e-08 w=4e-07 $X=27858 $Y=35682 $D=636
M2668 377 379 vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=27879 $Y=33942 $D=636
M2669 b_pxca_n<2> 381 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=27910 $Y=1941 $D=636
M2670 381 382 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=27910 $Y=5141 $D=636
M2671 382 350 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=27910 $Y=8691 $D=636
M2672 383 350 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=27910 $Y=41842 $D=636
M2673 384 383 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=27910 $Y=44992 $D=636
M2674 t_pxca_n<2> 384 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=27910 $Y=46622 $D=636
M2675 vdd 323 317 vdd hvtpfet l=6e-08 w=7e-07 $X=27924 $Y=29648 $D=636
M2676 vdd 317 1289 vdd hvtpfet l=6e-08 w=8.23e-07 $X=27959 $Y=15520 $D=636
M2677 vdd 317 1290 vdd hvtpfet l=6e-08 w=8.23e-07 $X=27959 $Y=20589 $D=636
M2678 vdd 317 1291 vdd hvtpfet l=6e-08 w=8.23e-07 $X=27959 $Y=22440 $D=636
M2679 vdd 317 1292 vdd hvtpfet l=6e-08 w=8.23e-07 $X=27959 $Y=27509 $D=636
M2680 380 aa<11> vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=28044 $Y=14280 $D=636
M2681 386 356 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=28118 $Y=35682 $D=636
M2682 vdd 381 b_pxca_n<2> vdd hvtpfet l=6e-08 w=2.57e-06 $X=28170 $Y=1941 $D=636
M2683 vdd 382 381 vdd hvtpfet l=6e-08 w=1e-06 $X=28170 $Y=5141 $D=636
M2684 vdd 350 382 vdd hvtpfet l=6e-08 w=6e-07 $X=28170 $Y=8691 $D=636
M2685 vdd 350 383 vdd hvtpfet l=6e-08 w=6e-07 $X=28170 $Y=41842 $D=636
M2686 vdd 383 384 vdd hvtpfet l=6e-08 w=1e-06 $X=28170 $Y=44992 $D=636
M2687 vdd 384 t_pxca_n<2> vdd hvtpfet l=6e-08 w=2.57e-06 $X=28170 $Y=46622 $D=636
M2688 317 323 vdd vdd hvtpfet l=6e-08 w=7e-07 $X=28184 $Y=29648 $D=636
M2689 1293 317 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=28219 $Y=15520 $D=636
M2690 1294 317 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=28219 $Y=20589 $D=636
M2691 1295 317 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=28219 $Y=22440 $D=636
M2692 1296 317 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=28219 $Y=27509 $D=636
M2693 vdd 323 317 vdd hvtpfet l=6e-08 w=7e-07 $X=28444 $Y=29648 $D=636
M2694 407 374 1293 vdd hvtpfet l=6e-08 w=4.11e-07 $X=28489 $Y=15932 $D=636
M2695 408 375 1294 vdd hvtpfet l=6e-08 w=4.11e-07 $X=28489 $Y=20589 $D=636
M2696 409 374 1295 vdd hvtpfet l=6e-08 w=4.11e-07 $X=28489 $Y=22852 $D=636
M2697 410 375 1296 vdd hvtpfet l=6e-08 w=4.11e-07 $X=28489 $Y=27509 $D=636
M2698 vdd 392 541 vdd hvtpfet l=6e-08 w=4e-07 $X=28514 $Y=10167 $D=636
M2699 vdd 393 544 vdd hvtpfet l=6e-08 w=4e-07 $X=28514 $Y=40566 $D=636
M2700 494 386 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=28628 $Y=35682 $D=636
M2701 b_pxca_n<1> 387 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=28680 $Y=1941 $D=636
M2702 387 388 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=28680 $Y=5141 $D=636
M2703 388 389 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=28680 $Y=8691 $D=636
M2704 390 389 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=28680 $Y=41842 $D=636
M2705 391 390 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=28680 $Y=44992 $D=636
M2706 t_pxca_n<1> 391 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=28680 $Y=46622 $D=636
M2707 742 123 vdd vdd hvtpfet l=6e-08 w=1.2e-06 $X=28704 $Y=29148 $D=636
M2708 vdd 387 b_pxca_n<1> vdd hvtpfet l=6e-08 w=2.57e-06 $X=28940 $Y=1941 $D=636
M2709 vdd 388 387 vdd hvtpfet l=6e-08 w=1e-06 $X=28940 $Y=5141 $D=636
M2710 vdd 389 388 vdd hvtpfet l=6e-08 w=6e-07 $X=28940 $Y=8691 $D=636
M2711 vdd 389 390 vdd hvtpfet l=6e-08 w=6e-07 $X=28940 $Y=41842 $D=636
M2712 vdd 390 391 vdd hvtpfet l=6e-08 w=1e-06 $X=28940 $Y=44992 $D=636
M2713 vdd 391 t_pxca_n<1> vdd hvtpfet l=6e-08 w=2.57e-06 $X=28940 $Y=46622 $D=636
M2714 1297 317 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=28999 $Y=15520 $D=636
M2715 1298 317 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=28999 $Y=20589 $D=636
M2716 1299 317 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=28999 $Y=22440 $D=636
M2717 1300 317 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=28999 $Y=27509 $D=636
M2718 vdd 308 392 vdd hvtpfet l=6e-08 w=4.11e-07 $X=29024 $Y=10156 $D=636
M2719 vdd 308 393 vdd hvtpfet l=6e-08 w=4.11e-07 $X=29024 $Y=40566 $D=636
M2720 vdd aa<12> 365 vdd hvtpfet l=6e-08 w=4.11e-07 $X=29054 $Y=14280 $D=636
M2721 407 380 1297 vdd hvtpfet l=6e-08 w=4.11e-07 $X=29269 $Y=15932 $D=636
M2722 408 380 1298 vdd hvtpfet l=6e-08 w=4.11e-07 $X=29269 $Y=20589 $D=636
M2723 409 380 1299 vdd hvtpfet l=6e-08 w=4.11e-07 $X=29269 $Y=22852 $D=636
M2724 410 380 1300 vdd hvtpfet l=6e-08 w=4.11e-07 $X=29269 $Y=27509 $D=636
M2725 392 dwla<1> vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=29284 $Y=10156 $D=636
M2726 393 dwla<0> vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=29284 $Y=40566 $D=636
M2727 743 395 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=29298 $Y=33468 $D=636
M2728 b_pxca_n<0> 396 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=29450 $Y=1941 $D=636
M2729 396 397 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=29450 $Y=5141 $D=636
M2730 397 398 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=29450 $Y=8691 $D=636
M2731 399 398 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=29450 $Y=41842 $D=636
M2732 400 399 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=29450 $Y=44992 $D=636
M2733 t_pxca_n<0> 400 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=29450 $Y=46622 $D=636
M2734 748 403 456 vdd hvtpfet l=6e-08 w=1e-06 $X=29487 $Y=35707 $D=636
M2735 1301 364 407 vdd hvtpfet l=6e-08 w=4.11e-07 $X=29529 $Y=15932 $D=636
M2736 1302 364 408 vdd hvtpfet l=6e-08 w=4.11e-07 $X=29529 $Y=20589 $D=636
M2737 1303 365 409 vdd hvtpfet l=6e-08 w=4.11e-07 $X=29529 $Y=22852 $D=636
M2738 1304 365 410 vdd hvtpfet l=6e-08 w=4.11e-07 $X=29529 $Y=27509 $D=636
M2739 403 405 743 vdd hvtpfet l=6e-08 w=6e-07 $X=29558 $Y=33468 $D=636
M2740 364 365 vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=29564 $Y=14280 $D=636
M2741 vdd 404 395 vdd hvtpfet l=2.5e-07 w=5e-07 $X=29591 $Y=29813 $D=636
M2742 vdd 396 b_pxca_n<0> vdd hvtpfet l=6e-08 w=2.57e-06 $X=29710 $Y=1941 $D=636
M2743 vdd 397 396 vdd hvtpfet l=6e-08 w=1e-06 $X=29710 $Y=5141 $D=636
M2744 vdd 398 397 vdd hvtpfet l=6e-08 w=6e-07 $X=29710 $Y=8691 $D=636
M2745 vdd 398 399 vdd hvtpfet l=6e-08 w=6e-07 $X=29710 $Y=41842 $D=636
M2746 vdd 399 400 vdd hvtpfet l=6e-08 w=1e-06 $X=29710 $Y=44992 $D=636
M2747 vdd 400 t_pxca_n<0> vdd hvtpfet l=6e-08 w=2.57e-06 $X=29710 $Y=46622 $D=636
M2748 456 403 748 vdd hvtpfet l=6e-08 w=1e-06 $X=29747 $Y=35707 $D=636
M2749 vdd 317 1301 vdd hvtpfet l=6e-08 w=8.23e-07 $X=29799 $Y=15520 $D=636
M2750 vdd 317 1302 vdd hvtpfet l=6e-08 w=8.23e-07 $X=29799 $Y=20589 $D=636
M2751 vdd 317 1303 vdd hvtpfet l=6e-08 w=8.23e-07 $X=29799 $Y=22440 $D=636
M2752 vdd 317 1304 vdd hvtpfet l=6e-08 w=8.23e-07 $X=29799 $Y=27509 $D=636
M2753 748 403 456 vdd hvtpfet l=6e-08 w=1e-06 $X=30007 $Y=35707 $D=636
M2754 404 406 vdd vdd hvtpfet l=6e-08 w=5e-07 $X=30041 $Y=29813 $D=636
M2755 405 tm<7> vdd vdd hvtpfet l=6e-08 w=3e-07 $X=30068 $Y=33468 $D=636
M2756 dbl_pd_n<3> 131 vdd vdd hvtpfet l=6e-08 w=4.28e-07 $X=30204 $Y=14263 $D=636
M2757 b_pxba_n<7> 411 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=30220 $Y=1941 $D=636
M2758 411 412 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=30220 $Y=5141 $D=636
M2759 412 413 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=30220 $Y=8691 $D=636
M2760 414 413 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=30220 $Y=41842 $D=636
M2761 415 414 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=30220 $Y=44992 $D=636
M2762 t_pxba_n<7> 415 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=30220 $Y=46622 $D=636
M2763 753 416 748 vdd hvtpfet l=6e-08 w=1e-06 $X=30267 $Y=35707 $D=636
M2764 359 407 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=30309 $Y=15321 $D=636
M2765 1305 323 407 vdd hvtpfet l=6e-08 w=2.74e-07 $X=30309 $Y=16069 $D=636
M2766 1306 323 408 vdd hvtpfet l=6e-08 w=2.74e-07 $X=30309 $Y=20589 $D=636
M2767 347 408 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=30309 $Y=21405 $D=636
M2768 398 409 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=30309 $Y=22241 $D=636
M2769 1307 323 409 vdd hvtpfet l=6e-08 w=2.74e-07 $X=30309 $Y=22989 $D=636
M2770 1308 323 410 vdd hvtpfet l=6e-08 w=2.74e-07 $X=30309 $Y=27509 $D=636
M2771 389 410 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=30309 $Y=28325 $D=636
M2772 vdd 131 dbl_pd_n<3> vdd hvtpfet l=6e-08 w=4.28e-07 $X=30464 $Y=14263 $D=636
M2773 vdd 411 b_pxba_n<7> vdd hvtpfet l=6e-08 w=2.57e-06 $X=30480 $Y=1941 $D=636
M2774 vdd 412 411 vdd hvtpfet l=6e-08 w=1e-06 $X=30480 $Y=5141 $D=636
M2775 vdd 413 412 vdd hvtpfet l=6e-08 w=6e-07 $X=30480 $Y=8691 $D=636
M2776 vdd 413 414 vdd hvtpfet l=6e-08 w=6e-07 $X=30480 $Y=41842 $D=636
M2777 vdd 414 415 vdd hvtpfet l=6e-08 w=1e-06 $X=30480 $Y=44992 $D=636
M2778 vdd 415 t_pxba_n<7> vdd hvtpfet l=6e-08 w=2.57e-06 $X=30480 $Y=46622 $D=636
M2779 748 416 753 vdd hvtpfet l=6e-08 w=1e-06 $X=30527 $Y=35707 $D=636
M2780 vdd 407 359 vdd hvtpfet l=6e-08 w=2.06e-07 $X=30569 $Y=15321 $D=636
M2781 vdd 359 1305 vdd hvtpfet l=6e-08 w=2.74e-07 $X=30569 $Y=16069 $D=636
M2782 vdd 347 1306 vdd hvtpfet l=6e-08 w=2.74e-07 $X=30569 $Y=20589 $D=636
M2783 vdd 408 347 vdd hvtpfet l=6e-08 w=2.06e-07 $X=30569 $Y=21405 $D=636
M2784 vdd 409 398 vdd hvtpfet l=6e-08 w=2.06e-07 $X=30569 $Y=22241 $D=636
M2785 vdd 398 1307 vdd hvtpfet l=6e-08 w=2.74e-07 $X=30569 $Y=22989 $D=636
M2786 vdd 389 1308 vdd hvtpfet l=6e-08 w=2.74e-07 $X=30569 $Y=27509 $D=636
M2787 vdd 410 389 vdd hvtpfet l=6e-08 w=2.06e-07 $X=30569 $Y=28325 $D=636
M2788 vdd dwla<1> 426 vdd hvtpfet l=6e-08 w=4.11e-07 $X=30584 $Y=10156 $D=636
M2789 vdd dwla<0> 427 vdd hvtpfet l=6e-08 w=4.11e-07 $X=30584 $Y=40566 $D=636
M2790 749 406 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=30644 $Y=33468 $D=636
M2791 vdd 417 406 vdd hvtpfet l=2.5e-07 w=5e-07 $X=30711 $Y=29813 $D=636
M2792 dbl_pd_n<3> 131 vdd vdd hvtpfet l=6e-08 w=4.28e-07 $X=30724 $Y=14263 $D=636
M2793 753 416 748 vdd hvtpfet l=6e-08 w=1e-06 $X=30787 $Y=35707 $D=636
M2794 426 309 vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=30844 $Y=10156 $D=636
M2795 427 309 vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=30844 $Y=40566 $D=636
M2796 416 423 749 vdd hvtpfet l=6e-08 w=6e-07 $X=30904 $Y=33468 $D=636
M2797 b_pxba_n<6> 418 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=30990 $Y=1941 $D=636
M2798 418 419 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=30990 $Y=5141 $D=636
M2799 419 420 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=30990 $Y=8691 $D=636
M2800 421 420 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=30990 $Y=41842 $D=636
M2801 422 421 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=30990 $Y=44992 $D=636
M2802 t_pxba_n<6> 422 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=30990 $Y=46622 $D=636
M2803 vdd 362 753 vdd hvtpfet l=6e-08 w=1e-06 $X=31047 $Y=35707 $D=636
M2804 420 428 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=31079 $Y=15321 $D=636
M2805 1309 420 vdd vdd hvtpfet l=6e-08 w=2.74e-07 $X=31079 $Y=16069 $D=636
M2806 1310 413 vdd vdd hvtpfet l=6e-08 w=2.74e-07 $X=31079 $Y=20589 $D=636
M2807 413 429 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=31079 $Y=21405 $D=636
M2808 424 430 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=31079 $Y=22241 $D=636
M2809 1311 424 vdd vdd hvtpfet l=6e-08 w=2.74e-07 $X=31079 $Y=22989 $D=636
M2810 1312 425 vdd vdd hvtpfet l=6e-08 w=2.74e-07 $X=31079 $Y=27509 $D=636
M2811 425 431 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=31079 $Y=28325 $D=636
M2812 417 368 vdd vdd hvtpfet l=6e-08 w=5e-07 $X=31161 $Y=29813 $D=636
M2813 dbl_pd_n<1> tm<1> vdd vdd hvtpfet l=6e-08 w=4.28e-07 $X=31234 $Y=14263 $D=636
M2814 vdd 418 b_pxba_n<6> vdd hvtpfet l=6e-08 w=2.57e-06 $X=31250 $Y=1941 $D=636
M2815 vdd 419 418 vdd hvtpfet l=6e-08 w=1e-06 $X=31250 $Y=5141 $D=636
M2816 vdd 420 419 vdd hvtpfet l=6e-08 w=6e-07 $X=31250 $Y=8691 $D=636
M2817 vdd 420 421 vdd hvtpfet l=6e-08 w=6e-07 $X=31250 $Y=41842 $D=636
M2818 vdd 421 422 vdd hvtpfet l=6e-08 w=1e-06 $X=31250 $Y=44992 $D=636
M2819 vdd 422 t_pxba_n<6> vdd hvtpfet l=6e-08 w=2.57e-06 $X=31250 $Y=46622 $D=636
M2820 753 362 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=31307 $Y=35707 $D=636
M2821 vdd 428 420 vdd hvtpfet l=6e-08 w=2.06e-07 $X=31339 $Y=15321 $D=636
M2822 428 323 1309 vdd hvtpfet l=6e-08 w=2.74e-07 $X=31339 $Y=16069 $D=636
M2823 429 323 1310 vdd hvtpfet l=6e-08 w=2.74e-07 $X=31339 $Y=20589 $D=636
M2824 vdd 429 413 vdd hvtpfet l=6e-08 w=2.06e-07 $X=31339 $Y=21405 $D=636
M2825 vdd 430 424 vdd hvtpfet l=6e-08 w=2.06e-07 $X=31339 $Y=22241 $D=636
M2826 430 323 1311 vdd hvtpfet l=6e-08 w=2.74e-07 $X=31339 $Y=22989 $D=636
M2827 431 323 1312 vdd hvtpfet l=6e-08 w=2.74e-07 $X=31339 $Y=27509 $D=636
M2828 vdd 431 425 vdd hvtpfet l=6e-08 w=2.06e-07 $X=31339 $Y=28325 $D=636
M2829 556 426 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=31354 $Y=10167 $D=636
M2830 558 427 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=31354 $Y=40566 $D=636
M2831 vdd 173 423 vdd hvtpfet l=6e-08 w=3e-07 $X=31414 $Y=33468 $D=636
M2832 vdd tm<1> dbl_pd_n<1> vdd hvtpfet l=6e-08 w=4.28e-07 $X=31494 $Y=14263 $D=636
M2833 vdd 362 753 vdd hvtpfet l=6e-08 w=1e-06 $X=31567 $Y=35707 $D=636
M2834 dbl_pd_n<1> tm<1> vdd vdd hvtpfet l=6e-08 w=4.28e-07 $X=31754 $Y=14263 $D=636
M2835 b_pxba_n<5> 432 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=31760 $Y=1941 $D=636
M2836 432 433 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=31760 $Y=5141 $D=636
M2837 433 434 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=31760 $Y=8691 $D=636
M2838 435 434 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=31760 $Y=41842 $D=636
M2839 436 435 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=31760 $Y=44992 $D=636
M2840 t_pxba_n<5> 436 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=31760 $Y=46622 $D=636
M2841 vdd 368 362 vdd hvtpfet l=6e-08 w=4e-07 $X=31761 $Y=29948 $D=636
M2842 1313 317 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=31849 $Y=15520 $D=636
M2843 1314 317 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=31849 $Y=20589 $D=636
M2844 1315 317 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=31849 $Y=22440 $D=636
M2845 1316 317 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=31849 $Y=27509 $D=636
M2846 vdd 437 540 vdd hvtpfet l=6e-08 w=4e-07 $X=31864 $Y=10167 $D=636
M2847 vdd 438 545 vdd hvtpfet l=6e-08 w=4e-07 $X=31864 $Y=40566 $D=636
M2848 vdd 432 b_pxba_n<5> vdd hvtpfet l=6e-08 w=2.57e-06 $X=32020 $Y=1941 $D=636
M2849 vdd 433 432 vdd hvtpfet l=6e-08 w=1e-06 $X=32020 $Y=5141 $D=636
M2850 vdd 434 433 vdd hvtpfet l=6e-08 w=6e-07 $X=32020 $Y=8691 $D=636
M2851 vdd 434 435 vdd hvtpfet l=6e-08 w=6e-07 $X=32020 $Y=41842 $D=636
M2852 vdd 435 436 vdd hvtpfet l=6e-08 w=1e-06 $X=32020 $Y=44992 $D=636
M2853 vdd 436 t_pxba_n<5> vdd hvtpfet l=6e-08 w=2.57e-06 $X=32020 $Y=46622 $D=636
M2854 428 439 1313 vdd hvtpfet l=6e-08 w=4.11e-07 $X=32119 $Y=15932 $D=636
M2855 429 439 1314 vdd hvtpfet l=6e-08 w=4.11e-07 $X=32119 $Y=20589 $D=636
M2856 430 440 1315 vdd hvtpfet l=6e-08 w=4.11e-07 $X=32119 $Y=22852 $D=636
M2857 431 440 1316 vdd hvtpfet l=6e-08 w=4.11e-07 $X=32119 $Y=27509 $D=636
M2858 761 442 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=32271 $Y=29348 $D=636
M2859 762 442 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=32271 $Y=35707 $D=636
M2860 vdd 310 437 vdd hvtpfet l=6e-08 w=4.11e-07 $X=32374 $Y=10156 $D=636
M2861 vdd 310 438 vdd hvtpfet l=6e-08 w=4.11e-07 $X=32374 $Y=40566 $D=636
M2862 1317 443 428 vdd hvtpfet l=6e-08 w=4.11e-07 $X=32379 $Y=15932 $D=636
M2863 1318 443 429 vdd hvtpfet l=6e-08 w=4.11e-07 $X=32379 $Y=20589 $D=636
M2864 1319 443 430 vdd hvtpfet l=6e-08 w=4.11e-07 $X=32379 $Y=22852 $D=636
M2865 1320 443 431 vdd hvtpfet l=6e-08 w=4.11e-07 $X=32379 $Y=27509 $D=636
M2866 vdd aa<7> 449 vdd hvtpfet l=6e-08 w=4.11e-07 $X=32394 $Y=14280 $D=636
M2867 vdd 324 442 vdd hvtpfet l=6e-08 w=1e-06 $X=32394 $Y=33493 $D=636
M2868 b_pxba_n<4> 444 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=32530 $Y=1941 $D=636
M2869 444 445 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=32530 $Y=5141 $D=636
M2870 445 446 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=32530 $Y=8691 $D=636
M2871 447 446 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=32530 $Y=41842 $D=636
M2872 448 447 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=32530 $Y=44992 $D=636
M2873 t_pxba_n<4> 448 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=32530 $Y=46622 $D=636
M2874 vdd 442 761 vdd hvtpfet l=6e-08 w=1e-06 $X=32531 $Y=29348 $D=636
M2875 vdd 442 762 vdd hvtpfet l=6e-08 w=1e-06 $X=32531 $Y=35707 $D=636
M2876 437 dwla<1> vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=32634 $Y=10156 $D=636
M2877 438 dwla<0> vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=32634 $Y=40566 $D=636
M2878 vdd 317 1317 vdd hvtpfet l=6e-08 w=8.23e-07 $X=32649 $Y=15520 $D=636
M2879 vdd 317 1318 vdd hvtpfet l=6e-08 w=8.23e-07 $X=32649 $Y=20589 $D=636
M2880 vdd 317 1319 vdd hvtpfet l=6e-08 w=8.23e-07 $X=32649 $Y=22440 $D=636
M2881 vdd 317 1320 vdd hvtpfet l=6e-08 w=8.23e-07 $X=32649 $Y=27509 $D=636
M2882 450 449 vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=32654 $Y=14280 $D=636
M2883 vdd 444 b_pxba_n<4> vdd hvtpfet l=6e-08 w=2.57e-06 $X=32790 $Y=1941 $D=636
M2884 vdd 445 444 vdd hvtpfet l=6e-08 w=1e-06 $X=32790 $Y=5141 $D=636
M2885 vdd 446 445 vdd hvtpfet l=6e-08 w=6e-07 $X=32790 $Y=8691 $D=636
M2886 vdd 446 447 vdd hvtpfet l=6e-08 w=6e-07 $X=32790 $Y=41842 $D=636
M2887 vdd 447 448 vdd hvtpfet l=6e-08 w=1e-06 $X=32790 $Y=44992 $D=636
M2888 vdd 448 t_pxba_n<4> vdd hvtpfet l=6e-08 w=2.57e-06 $X=32790 $Y=46622 $D=636
M2889 dwla<1> 368 761 vdd hvtpfet l=6e-08 w=1e-06 $X=33041 $Y=29348 $D=636
M2890 497 456 762 vdd hvtpfet l=6e-08 w=1e-06 $X=33041 $Y=35707 $D=636
M2891 465 442 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=33094 $Y=33493 $D=636
M2892 vdd dwla<1> 458 vdd hvtpfet l=6e-08 w=4.11e-07 $X=33144 $Y=10156 $D=636
M2893 vdd dwla<0> 459 vdd hvtpfet l=6e-08 w=4.11e-07 $X=33144 $Y=40566 $D=636
M2894 1321 449 428 vdd hvtpfet l=6e-08 w=4.11e-07 $X=33159 $Y=15932 $D=636
M2895 1322 450 429 vdd hvtpfet l=6e-08 w=4.11e-07 $X=33159 $Y=20589 $D=636
M2896 1323 449 430 vdd hvtpfet l=6e-08 w=4.11e-07 $X=33159 $Y=22852 $D=636
M2897 1324 450 431 vdd hvtpfet l=6e-08 w=4.11e-07 $X=33159 $Y=27509 $D=636
M2898 vdd 455 443 vdd hvtpfet l=6e-08 w=4.11e-07 $X=33254 $Y=14280 $D=636
M2899 b_pxba_n<3> 451 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=33300 $Y=1941 $D=636
M2900 451 452 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=33300 $Y=5141 $D=636
M2901 452 425 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=33300 $Y=8691 $D=636
M2902 453 425 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=33300 $Y=41842 $D=636
M2903 454 453 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=33300 $Y=44992 $D=636
M2904 t_pxba_n<3> 454 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=33300 $Y=46622 $D=636
M2905 761 368 dwla<1> vdd hvtpfet l=6e-08 w=1e-06 $X=33301 $Y=29348 $D=636
M2906 762 456 497 vdd hvtpfet l=6e-08 w=1e-06 $X=33301 $Y=35707 $D=636
M2907 458 311 vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=33404 $Y=10156 $D=636
M2908 459 311 vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=33404 $Y=40566 $D=636
M2909 vdd 317 1321 vdd hvtpfet l=6e-08 w=8.23e-07 $X=33429 $Y=15520 $D=636
M2910 vdd 317 1322 vdd hvtpfet l=6e-08 w=8.23e-07 $X=33429 $Y=20589 $D=636
M2911 vdd 317 1323 vdd hvtpfet l=6e-08 w=8.23e-07 $X=33429 $Y=22440 $D=636
M2912 vdd 317 1324 vdd hvtpfet l=6e-08 w=8.23e-07 $X=33429 $Y=27509 $D=636
M2913 455 aa<8> vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=33514 $Y=14280 $D=636
M2914 vdd 451 b_pxba_n<3> vdd hvtpfet l=6e-08 w=2.57e-06 $X=33560 $Y=1941 $D=636
M2915 vdd 452 451 vdd hvtpfet l=6e-08 w=1e-06 $X=33560 $Y=5141 $D=636
M2916 vdd 425 452 vdd hvtpfet l=6e-08 w=6e-07 $X=33560 $Y=8691 $D=636
M2917 vdd 425 453 vdd hvtpfet l=6e-08 w=6e-07 $X=33560 $Y=41842 $D=636
M2918 vdd 453 454 vdd hvtpfet l=6e-08 w=1e-06 $X=33560 $Y=44992 $D=636
M2919 vdd 454 t_pxba_n<3> vdd hvtpfet l=6e-08 w=2.57e-06 $X=33560 $Y=46622 $D=636
M2920 1325 317 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=33689 $Y=15520 $D=636
M2921 1326 317 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=33689 $Y=20589 $D=636
M2922 1327 317 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=33689 $Y=22440 $D=636
M2923 1328 317 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=33689 $Y=27509 $D=636
M2924 dwla<0> 368 765 vdd hvtpfet l=6e-08 w=1e-06 $X=33811 $Y=29348 $D=636
M2925 498 456 766 vdd hvtpfet l=6e-08 w=1e-06 $X=33811 $Y=35707 $D=636
M2926 555 458 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=33914 $Y=10167 $D=636
M2927 559 459 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=33914 $Y=40566 $D=636
M2928 479 449 1325 vdd hvtpfet l=6e-08 w=4.11e-07 $X=33959 $Y=15932 $D=636
M2929 480 450 1326 vdd hvtpfet l=6e-08 w=4.11e-07 $X=33959 $Y=20589 $D=636
M2930 481 449 1327 vdd hvtpfet l=6e-08 w=4.11e-07 $X=33959 $Y=22852 $D=636
M2931 482 450 1328 vdd hvtpfet l=6e-08 w=4.11e-07 $X=33959 $Y=27509 $D=636
M2932 b_pxba_n<2> 460 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=34070 $Y=1941 $D=636
M2933 460 461 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=34070 $Y=5141 $D=636
M2934 461 424 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=34070 $Y=8691 $D=636
M2935 462 424 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=34070 $Y=41842 $D=636
M2936 463 462 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=34070 $Y=44992 $D=636
M2937 t_pxba_n<2> 463 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=34070 $Y=46622 $D=636
M2938 765 368 dwla<0> vdd hvtpfet l=6e-08 w=1e-06 $X=34071 $Y=29348 $D=636
M2939 766 456 498 vdd hvtpfet l=6e-08 w=1e-06 $X=34071 $Y=35707 $D=636
M2940 vdd 460 b_pxba_n<2> vdd hvtpfet l=6e-08 w=2.57e-06 $X=34330 $Y=1941 $D=636
M2941 vdd 461 460 vdd hvtpfet l=6e-08 w=1e-06 $X=34330 $Y=5141 $D=636
M2942 vdd 424 461 vdd hvtpfet l=6e-08 w=6e-07 $X=34330 $Y=8691 $D=636
M2943 vdd 424 462 vdd hvtpfet l=6e-08 w=6e-07 $X=34330 $Y=41842 $D=636
M2944 vdd 462 463 vdd hvtpfet l=6e-08 w=1e-06 $X=34330 $Y=44992 $D=636
M2945 vdd 463 t_pxba_n<2> vdd hvtpfet l=6e-08 w=2.57e-06 $X=34330 $Y=46622 $D=636
M2946 1329 317 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=34469 $Y=15520 $D=636
M2947 1330 317 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=34469 $Y=20589 $D=636
M2948 1331 317 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=34469 $Y=22440 $D=636
M2949 1332 317 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=34469 $Y=27509 $D=636
M2950 vdd aa<9> 440 vdd hvtpfet l=6e-08 w=4.11e-07 $X=34524 $Y=14280 $D=636
M2951 765 465 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=34581 $Y=29348 $D=636
M2952 766 465 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=34581 $Y=35707 $D=636
M2953 vdd vdd 535 vdd hvtpfet l=6e-08 w=6.4e-07 $X=34621 $Y=33468 $D=636
M2954 479 455 1329 vdd hvtpfet l=6e-08 w=4.11e-07 $X=34739 $Y=15932 $D=636
M2955 480 455 1330 vdd hvtpfet l=6e-08 w=4.11e-07 $X=34739 $Y=20589 $D=636
M2956 481 455 1331 vdd hvtpfet l=6e-08 w=4.11e-07 $X=34739 $Y=22852 $D=636
M2957 482 455 1332 vdd hvtpfet l=6e-08 w=4.11e-07 $X=34739 $Y=27509 $D=636
M2958 b_pxba_n<1> 466 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=34840 $Y=1941 $D=636
M2959 466 467 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=34840 $Y=5141 $D=636
M2960 467 468 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=34840 $Y=8691 $D=636
M2961 469 468 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=34840 $Y=41842 $D=636
M2962 470 469 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=34840 $Y=44992 $D=636
M2963 t_pxba_n<1> 470 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=34840 $Y=46622 $D=636
M2964 vdd 465 765 vdd hvtpfet l=6e-08 w=1e-06 $X=34841 $Y=29348 $D=636
M2965 vdd 465 766 vdd hvtpfet l=6e-08 w=1e-06 $X=34841 $Y=35707 $D=636
M2966 535 471 vdd vdd hvtpfet l=6e-08 w=6.4e-07 $X=34881 $Y=33468 $D=636
M2967 vdd 123 131 vdd hvtpfet l=6e-08 w=2e-07 $X=34906 $Y=10756 $D=636
M2968 1333 439 479 vdd hvtpfet l=6e-08 w=4.11e-07 $X=34999 $Y=15932 $D=636
M2969 1334 439 480 vdd hvtpfet l=6e-08 w=4.11e-07 $X=34999 $Y=20589 $D=636
M2970 1335 440 481 vdd hvtpfet l=6e-08 w=4.11e-07 $X=34999 $Y=22852 $D=636
M2971 1336 440 482 vdd hvtpfet l=6e-08 w=4.11e-07 $X=34999 $Y=27509 $D=636
M2972 439 440 vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=35034 $Y=14280 $D=636
M2973 vdd 466 b_pxba_n<1> vdd hvtpfet l=6e-08 w=2.57e-06 $X=35100 $Y=1941 $D=636
M2974 vdd 467 466 vdd hvtpfet l=6e-08 w=1e-06 $X=35100 $Y=5141 $D=636
M2975 vdd 468 467 vdd hvtpfet l=6e-08 w=6e-07 $X=35100 $Y=8691 $D=636
M2976 vdd 468 469 vdd hvtpfet l=6e-08 w=6e-07 $X=35100 $Y=41842 $D=636
M2977 vdd 469 470 vdd hvtpfet l=6e-08 w=1e-06 $X=35100 $Y=44992 $D=636
M2978 vdd 470 t_pxba_n<1> vdd hvtpfet l=6e-08 w=2.57e-06 $X=35100 $Y=46622 $D=636
M2979 vdd 317 1333 vdd hvtpfet l=6e-08 w=8.23e-07 $X=35269 $Y=15520 $D=636
M2980 vdd 317 1334 vdd hvtpfet l=6e-08 w=8.23e-07 $X=35269 $Y=20589 $D=636
M2981 vdd 317 1335 vdd hvtpfet l=6e-08 w=8.23e-07 $X=35269 $Y=22440 $D=636
M2982 vdd 317 1336 vdd hvtpfet l=6e-08 w=8.23e-07 $X=35269 $Y=27509 $D=636
M2983 vdd 473 484 vdd hvtpfet l=6e-08 w=3e-07 $X=35351 $Y=36377 $D=636
M2984 vdd 472 471 vdd hvtpfet l=2.5e-07 w=5e-07 $X=35416 $Y=33503 $D=636
M2985 b_pxba_n<0> 474 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=35610 $Y=1941 $D=636
M2986 474 475 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=35610 $Y=5141 $D=636
M2987 475 476 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=35610 $Y=8691 $D=636
M2988 477 476 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=35610 $Y=41842 $D=636
M2989 478 477 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=35610 $Y=44992 $D=636
M2990 t_pxba_n<0> 478 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=35610 $Y=46622 $D=636
M2991 446 479 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=35779 $Y=15321 $D=636
M2992 1337 323 479 vdd hvtpfet l=6e-08 w=2.74e-07 $X=35779 $Y=16069 $D=636
M2993 1338 323 480 vdd hvtpfet l=6e-08 w=2.74e-07 $X=35779 $Y=20589 $D=636
M2994 434 480 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=35779 $Y=21405 $D=636
M2995 476 481 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=35779 $Y=22241 $D=636
M2996 1339 323 481 vdd hvtpfet l=6e-08 w=2.74e-07 $X=35779 $Y=22989 $D=636
M2997 1340 323 482 vdd hvtpfet l=6e-08 w=2.74e-07 $X=35779 $Y=27509 $D=636
M2998 468 482 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=35779 $Y=28325 $D=636
M2999 473 484 vdd vdd hvtpfet l=1.2e-07 w=3e-07 $X=35861 $Y=36382 $D=636
M3000 472 483 vdd vdd hvtpfet l=6e-08 w=5e-07 $X=35866 $Y=33503 $D=636
M3001 vdd 474 b_pxba_n<0> vdd hvtpfet l=6e-08 w=2.57e-06 $X=35870 $Y=1941 $D=636
M3002 vdd 475 474 vdd hvtpfet l=6e-08 w=1e-06 $X=35870 $Y=5141 $D=636
M3003 vdd 476 475 vdd hvtpfet l=6e-08 w=6e-07 $X=35870 $Y=8691 $D=636
M3004 vdd 476 477 vdd hvtpfet l=6e-08 w=6e-07 $X=35870 $Y=41842 $D=636
M3005 vdd 477 478 vdd hvtpfet l=6e-08 w=1e-06 $X=35870 $Y=44992 $D=636
M3006 vdd 478 t_pxba_n<0> vdd hvtpfet l=6e-08 w=2.57e-06 $X=35870 $Y=46622 $D=636
M3007 368 495 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=35945 $Y=29548 $D=636
M3008 vdd 479 446 vdd hvtpfet l=6e-08 w=2.06e-07 $X=36039 $Y=15321 $D=636
M3009 vdd 446 1337 vdd hvtpfet l=6e-08 w=2.74e-07 $X=36039 $Y=16069 $D=636
M3010 vdd 434 1338 vdd hvtpfet l=6e-08 w=2.74e-07 $X=36039 $Y=20589 $D=636
M3011 vdd 480 434 vdd hvtpfet l=6e-08 w=2.06e-07 $X=36039 $Y=21405 $D=636
M3012 vdd 481 476 vdd hvtpfet l=6e-08 w=2.06e-07 $X=36039 $Y=22241 $D=636
M3013 vdd 476 1339 vdd hvtpfet l=6e-08 w=2.74e-07 $X=36039 $Y=22989 $D=636
M3014 vdd 468 1340 vdd hvtpfet l=6e-08 w=2.74e-07 $X=36039 $Y=27509 $D=636
M3015 vdd 482 468 vdd hvtpfet l=6e-08 w=2.06e-07 $X=36039 $Y=28325 $D=636
M3016 vdd 495 368 vdd hvtpfet l=6e-08 w=8e-07 $X=36205 $Y=29548 $D=636
M3017 vdd 491 509 vdd hvtpfet l=6e-08 w=4.11e-07 $X=36254 $Y=14280 $D=636
M3018 b_pxaa<3> 485 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=36380 $Y=1941 $D=636
M3019 485 486 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=36380 $Y=5141 $D=636
M3020 486 487 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=36380 $Y=8691 $D=636
M3021 vdd 492 487 vdd hvtpfet l=6e-08 w=4.11e-07 $X=36380 $Y=10156 $D=636
M3022 vdd 492 488 vdd hvtpfet l=6e-08 w=4.11e-07 $X=36380 $Y=40566 $D=636
M3023 489 488 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=36380 $Y=41842 $D=636
M3024 490 489 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=36380 $Y=44992 $D=636
M3025 t_pxaa<3> 490 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=36380 $Y=46622 $D=636
M3026 vdd 493 473 vdd hvtpfet l=6e-08 w=6.4e-07 $X=36431 $Y=35802 $D=636
M3027 vdd 496 483 vdd hvtpfet l=6e-08 w=6.4e-07 $X=36466 $Y=33468 $D=636
M3028 vdd 485 b_pxaa<3> vdd hvtpfet l=6e-08 w=2.57e-06 $X=36640 $Y=1941 $D=636
M3029 vdd 486 485 vdd hvtpfet l=6e-08 w=1e-06 $X=36640 $Y=5141 $D=636
M3030 vdd 487 486 vdd hvtpfet l=6e-08 w=6e-07 $X=36640 $Y=8691 $D=636
M3031 487 497 vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=36640 $Y=10156 $D=636
M3032 488 498 vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=36640 $Y=40566 $D=636
M3033 vdd 488 489 vdd hvtpfet l=6e-08 w=6e-07 $X=36640 $Y=41842 $D=636
M3034 vdd 489 490 vdd hvtpfet l=6e-08 w=1e-06 $X=36640 $Y=44992 $D=636
M3035 vdd 490 t_pxaa<3> vdd hvtpfet l=6e-08 w=2.57e-06 $X=36640 $Y=46622 $D=636
M3036 368 clka vdd vdd hvtpfet l=6e-08 w=8e-07 $X=36715 $Y=29548 $D=636
M3037 491 aa<6> vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=36764 $Y=14280 $D=636
M3038 1341 317 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=36789 $Y=15520 $D=636
M3039 1342 317 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=36789 $Y=20589 $D=636
M3040 1343 317 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=36789 $Y=22440 $D=636
M3041 1344 317 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=36789 $Y=27509 $D=636
M3042 vdd clka 368 vdd hvtpfet l=6e-08 w=8e-07 $X=36975 $Y=29548 $D=636
M3043 vdd 473 496 vdd hvtpfet l=6e-08 w=6.4e-07 $X=36976 $Y=33693 $D=636
M3044 519 501 1341 vdd hvtpfet l=6e-08 w=4.11e-07 $X=37059 $Y=15932 $D=636
M3045 520 502 1342 vdd hvtpfet l=6e-08 w=4.11e-07 $X=37059 $Y=20589 $D=636
M3046 521 501 1343 vdd hvtpfet l=6e-08 w=4.11e-07 $X=37059 $Y=22852 $D=636
M3047 522 502 1344 vdd hvtpfet l=6e-08 w=4.11e-07 $X=37059 $Y=27509 $D=636
M3048 b_pxaa<2> 503 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=37150 $Y=1941 $D=636
M3049 503 504 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=37150 $Y=5141 $D=636
M3050 504 505 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=37150 $Y=8691 $D=636
M3051 vdd 497 505 vdd hvtpfet l=6e-08 w=4.11e-07 $X=37150 $Y=10156 $D=636
M3052 vdd 498 506 vdd hvtpfet l=6e-08 w=4.11e-07 $X=37150 $Y=40566 $D=636
M3053 507 506 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=37150 $Y=41842 $D=636
M3054 508 507 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=37150 $Y=44992 $D=636
M3055 t_pxaa<2> 508 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=37150 $Y=46622 $D=636
M3056 776 ddqa_n vdd vdd hvtpfet l=6e-08 w=6.4e-07 $X=37161 $Y=35802 $D=636
M3057 vdd 502 501 vdd hvtpfet l=6e-08 w=4.11e-07 $X=37274 $Y=14280 $D=636
M3058 1345 509 519 vdd hvtpfet l=6e-08 w=4.11e-07 $X=37319 $Y=15932 $D=636
M3059 1346 509 520 vdd hvtpfet l=6e-08 w=4.11e-07 $X=37319 $Y=20589 $D=636
M3060 1347 491 521 vdd hvtpfet l=6e-08 w=4.11e-07 $X=37319 $Y=22852 $D=636
M3061 1348 491 522 vdd hvtpfet l=6e-08 w=4.11e-07 $X=37319 $Y=27509 $D=636
M3062 vdd 503 b_pxaa<2> vdd hvtpfet l=6e-08 w=2.57e-06 $X=37410 $Y=1941 $D=636
M3063 vdd 504 503 vdd hvtpfet l=6e-08 w=1e-06 $X=37410 $Y=5141 $D=636
M3064 vdd 505 504 vdd hvtpfet l=6e-08 w=6e-07 $X=37410 $Y=8691 $D=636
M3065 505 510 vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=37410 $Y=10156 $D=636
M3066 506 510 vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=37410 $Y=40566 $D=636
M3067 vdd 506 507 vdd hvtpfet l=6e-08 w=6e-07 $X=37410 $Y=41842 $D=636
M3068 vdd 507 508 vdd hvtpfet l=6e-08 w=1e-06 $X=37410 $Y=44992 $D=636
M3069 vdd 508 t_pxaa<2> vdd hvtpfet l=6e-08 w=2.57e-06 $X=37410 $Y=46622 $D=636
M3070 493 ddqa 776 vdd hvtpfet l=6e-08 w=6.4e-07 $X=37421 $Y=35802 $D=636
M3071 vdd clka 524 vdd hvtpfet l=6e-08 w=1.2e-06 $X=37485 $Y=29148 $D=636
M3072 vdd 317 1345 vdd hvtpfet l=6e-08 w=8.23e-07 $X=37589 $Y=15520 $D=636
M3073 vdd 317 1346 vdd hvtpfet l=6e-08 w=8.23e-07 $X=37589 $Y=20589 $D=636
M3074 vdd 317 1347 vdd hvtpfet l=6e-08 w=8.23e-07 $X=37589 $Y=22440 $D=636
M3075 vdd 317 1348 vdd hvtpfet l=6e-08 w=8.23e-07 $X=37589 $Y=27509 $D=636
M3076 vdd 496 557 vdd hvtpfet l=6e-08 w=6.4e-07 $X=37661 $Y=33693 $D=636
M3077 502 aa<5> vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=37784 $Y=14280 $D=636
M3078 b_pxaa<1> 512 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=37920 $Y=1941 $D=636
M3079 512 513 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=37920 $Y=5141 $D=636
M3080 513 514 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=37920 $Y=8691 $D=636
M3081 vdd 523 514 vdd hvtpfet l=6e-08 w=4.11e-07 $X=37920 $Y=10156 $D=636
M3082 vdd 523 515 vdd hvtpfet l=6e-08 w=4.11e-07 $X=37920 $Y=40566 $D=636
M3083 516 515 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=37920 $Y=41842 $D=636
M3084 517 516 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=37920 $Y=44992 $D=636
M3085 t_pxaa<1> 517 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=37920 $Y=46622 $D=636
M3086 557 386 vdd vdd hvtpfet l=6e-08 w=6.4e-07 $X=37921 $Y=33693 $D=636
M3087 492 519 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=38099 $Y=15321 $D=636
M3088 1349 323 519 vdd hvtpfet l=6e-08 w=2.74e-07 $X=38099 $Y=16069 $D=636
M3089 1350 323 520 vdd hvtpfet l=6e-08 w=2.74e-07 $X=38099 $Y=20589 $D=636
M3090 510 520 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=38099 $Y=21405 $D=636
M3091 523 521 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=38099 $Y=22241 $D=636
M3092 1351 323 521 vdd hvtpfet l=6e-08 w=2.74e-07 $X=38099 $Y=22989 $D=636
M3093 1352 323 522 vdd hvtpfet l=6e-08 w=2.74e-07 $X=38099 $Y=27509 $D=636
M3094 525 522 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=38099 $Y=28325 $D=636
M3095 vdd 493 526 vdd hvtpfet l=1.4e-07 w=6.4e-07 $X=38141 $Y=36067 $D=636
M3096 vdd 512 b_pxaa<1> vdd hvtpfet l=6e-08 w=2.57e-06 $X=38180 $Y=1941 $D=636
M3097 vdd 513 512 vdd hvtpfet l=6e-08 w=1e-06 $X=38180 $Y=5141 $D=636
M3098 vdd 514 513 vdd hvtpfet l=6e-08 w=6e-07 $X=38180 $Y=8691 $D=636
M3099 514 497 vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=38180 $Y=10156 $D=636
M3100 515 498 vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=38180 $Y=40566 $D=636
M3101 vdd 515 516 vdd hvtpfet l=6e-08 w=6e-07 $X=38180 $Y=41842 $D=636
M3102 vdd 516 517 vdd hvtpfet l=6e-08 w=1e-06 $X=38180 $Y=44992 $D=636
M3103 vdd 517 t_pxaa<1> vdd hvtpfet l=6e-08 w=2.57e-06 $X=38180 $Y=46622 $D=636
M3104 1353 524 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=38255 $Y=29525 $D=636
M3105 vdd 519 492 vdd hvtpfet l=6e-08 w=2.06e-07 $X=38359 $Y=15321 $D=636
M3106 vdd 492 1349 vdd hvtpfet l=6e-08 w=2.74e-07 $X=38359 $Y=16069 $D=636
M3107 vdd 510 1350 vdd hvtpfet l=6e-08 w=2.74e-07 $X=38359 $Y=20589 $D=636
M3108 vdd 520 510 vdd hvtpfet l=6e-08 w=2.06e-07 $X=38359 $Y=21405 $D=636
M3109 vdd 521 523 vdd hvtpfet l=6e-08 w=2.06e-07 $X=38359 $Y=22241 $D=636
M3110 vdd 523 1351 vdd hvtpfet l=6e-08 w=2.74e-07 $X=38359 $Y=22989 $D=636
M3111 vdd 525 1352 vdd hvtpfet l=6e-08 w=2.74e-07 $X=38359 $Y=27509 $D=636
M3112 vdd 522 525 vdd hvtpfet l=6e-08 w=2.06e-07 $X=38359 $Y=28325 $D=636
M3113 779 494 vdd vdd hvtpfet l=6e-08 w=6.4e-07 $X=38431 $Y=33468 $D=636
M3114 780 526 vdd vdd hvtpfet l=1.4e-07 w=6.4e-07 $X=38481 $Y=36067 $D=636
M3115 534 495 1353 vdd hvtpfet l=6e-08 w=8.23e-07 $X=38515 $Y=29525 $D=636
M3116 vdd 533 546 vdd hvtpfet l=6e-08 w=4.11e-07 $X=38574 $Y=14280 $D=636
M3117 b_pxaa<0> 527 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=38690 $Y=1941 $D=636
M3118 527 528 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=38690 $Y=5141 $D=636
M3119 528 529 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=38690 $Y=8691 $D=636
M3120 vdd 497 529 vdd hvtpfet l=6e-08 w=4.11e-07 $X=38690 $Y=10156 $D=636
M3121 vdd 498 530 vdd hvtpfet l=6e-08 w=4.11e-07 $X=38690 $Y=40566 $D=636
M3122 531 530 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=38690 $Y=41842 $D=636
M3123 532 531 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=38690 $Y=44992 $D=636
M3124 t_pxaa<0> 532 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=38690 $Y=46622 $D=636
M3125 vdd 527 b_pxaa<0> vdd hvtpfet l=6e-08 w=2.57e-06 $X=38950 $Y=1941 $D=636
M3126 vdd 528 527 vdd hvtpfet l=6e-08 w=1e-06 $X=38950 $Y=5141 $D=636
M3127 vdd 529 528 vdd hvtpfet l=6e-08 w=6e-07 $X=38950 $Y=8691 $D=636
M3128 529 525 vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=38950 $Y=10156 $D=636
M3129 530 525 vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=38950 $Y=40566 $D=636
M3130 vdd 530 531 vdd hvtpfet l=6e-08 w=6e-07 $X=38950 $Y=41842 $D=636
M3131 vdd 531 532 vdd hvtpfet l=6e-08 w=1e-06 $X=38950 $Y=44992 $D=636
M3132 vdd 532 t_pxaa<0> vdd hvtpfet l=6e-08 w=2.57e-06 $X=38950 $Y=46622 $D=636
M3133 1354 534 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=39025 $Y=29525 $D=636
M3134 533 aa<3> vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=39084 $Y=14280 $D=636
M3135 1355 317 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=39109 $Y=15520 $D=636
M3136 1356 317 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=39109 $Y=20589 $D=636
M3137 1357 317 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=39109 $Y=22440 $D=636
M3138 1358 317 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=39109 $Y=27509 $D=636
M3139 vdd clka 323 vdd hvtpfet l=6e-08 w=6e-07 $X=39174 $Y=33747 $D=636
M3140 293 535 vdd vdd hvtpfet l=6e-08 w=1.2e-06 $X=39185 $Y=35277 $D=636
M3141 495 539 1354 vdd hvtpfet l=6e-08 w=8.23e-07 $X=39285 $Y=29525 $D=636
M3142 549 537 1355 vdd hvtpfet l=6e-08 w=4.11e-07 $X=39379 $Y=15932 $D=636
M3143 550 538 1356 vdd hvtpfet l=6e-08 w=4.11e-07 $X=39379 $Y=20589 $D=636
M3144 551 537 1357 vdd hvtpfet l=6e-08 w=4.11e-07 $X=39379 $Y=22852 $D=636
M3145 552 538 1358 vdd hvtpfet l=6e-08 w=4.11e-07 $X=39379 $Y=27509 $D=636
M3146 323 clka vdd vdd hvtpfet l=6e-08 w=6e-07 $X=39434 $Y=33747 $D=636
M3147 vdd 538 537 vdd hvtpfet l=6e-08 w=4.11e-07 $X=39594 $Y=14280 $D=636
M3148 1359 546 549 vdd hvtpfet l=6e-08 w=4.11e-07 $X=39639 $Y=15932 $D=636
M3149 1360 546 550 vdd hvtpfet l=6e-08 w=4.11e-07 $X=39639 $Y=20589 $D=636
M3150 1361 533 551 vdd hvtpfet l=6e-08 w=4.11e-07 $X=39639 $Y=22852 $D=636
M3151 1362 533 552 vdd hvtpfet l=6e-08 w=4.11e-07 $X=39639 $Y=27509 $D=636
M3152 vdd clka 323 vdd hvtpfet l=6e-08 w=6e-07 $X=39694 $Y=33747 $D=636
M3153 r_sa_prea_n 293 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=39695 $Y=35277 $D=636
M3154 289 540 vdd vdd hvtpfet l=6e-08 w=1.2e-06 $X=39705 $Y=1736 $D=636
M3155 290 541 vdd vdd hvtpfet l=6e-08 w=1.2e-06 $X=39705 $Y=3566 $D=636
M3156 291 542 vdd vdd hvtpfet l=6e-08 w=1.2e-06 $X=39705 $Y=8196 $D=636
M3157 292 543 vdd vdd hvtpfet l=6e-08 w=1.2e-06 $X=39705 $Y=10026 $D=636
M3158 294 543 vdd vdd hvtpfet l=6e-08 w=1.2e-06 $X=39705 $Y=39907 $D=636
M3159 295 542 vdd vdd hvtpfet l=6e-08 w=1.2e-06 $X=39705 $Y=41737 $D=636
M3160 296 544 vdd vdd hvtpfet l=6e-08 w=1.2e-06 $X=39705 $Y=46367 $D=636
M3161 297 545 vdd vdd hvtpfet l=6e-08 w=1.2e-06 $X=39705 $Y=48197 $D=636
M3162 vdd stclka 539 vdd hvtpfet l=6e-08 w=4.11e-07 $X=39795 $Y=29937 $D=636
M3163 vdd 317 1359 vdd hvtpfet l=6e-08 w=8.23e-07 $X=39909 $Y=15520 $D=636
M3164 vdd 317 1360 vdd hvtpfet l=6e-08 w=8.23e-07 $X=39909 $Y=20589 $D=636
M3165 vdd 317 1361 vdd hvtpfet l=6e-08 w=8.23e-07 $X=39909 $Y=22440 $D=636
M3166 vdd 317 1362 vdd hvtpfet l=6e-08 w=8.23e-07 $X=39909 $Y=27509 $D=636
M3167 323 clka vdd vdd hvtpfet l=6e-08 w=6e-07 $X=39954 $Y=33747 $D=636
M3168 vdd 293 r_sa_prea_n vdd hvtpfet l=6e-08 w=1.43e-06 $X=39955 $Y=35277 $D=636
M3169 538 aa<2> vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=40104 $Y=14280 $D=636
M3170 rb_ca<1> 289 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=40215 $Y=1506 $D=636
M3171 rb_ca<3> 290 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=40215 $Y=3566 $D=636
M3172 rb_ma<1> 291 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=40215 $Y=7966 $D=636
M3173 rb_ma<3> 292 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=40215 $Y=10026 $D=636
M3174 r_sa_prea_n 293 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=40215 $Y=35277 $D=636
M3175 rt_ma<3> 294 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=40215 $Y=39677 $D=636
M3176 rt_ma<1> 295 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=40215 $Y=41737 $D=636
M3177 rt_ca<3> 296 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=40215 $Y=46137 $D=636
M3178 rt_ca<1> 297 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=40215 $Y=48197 $D=636
M3179 543 549 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=40419 $Y=15321 $D=636
M3180 1363 323 549 vdd hvtpfet l=6e-08 w=2.74e-07 $X=40419 $Y=16069 $D=636
M3181 1364 323 550 vdd hvtpfet l=6e-08 w=2.74e-07 $X=40419 $Y=20589 $D=636
M3182 553 550 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=40419 $Y=21405 $D=636
M3183 542 551 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=40419 $Y=22241 $D=636
M3184 1365 323 551 vdd hvtpfet l=6e-08 w=2.74e-07 $X=40419 $Y=22989 $D=636
M3185 1366 323 552 vdd hvtpfet l=6e-08 w=2.74e-07 $X=40419 $Y=27509 $D=636
M3186 554 552 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=40419 $Y=28325 $D=636
M3187 vdd 289 rb_ca<1> vdd hvtpfet l=6e-08 w=1.43e-06 $X=40475 $Y=1506 $D=636
M3188 vdd 290 rb_ca<3> vdd hvtpfet l=6e-08 w=1.43e-06 $X=40475 $Y=3566 $D=636
M3189 vdd 291 rb_ma<1> vdd hvtpfet l=6e-08 w=1.43e-06 $X=40475 $Y=7966 $D=636
M3190 vdd 292 rb_ma<3> vdd hvtpfet l=6e-08 w=1.43e-06 $X=40475 $Y=10026 $D=636
M3191 vdd 294 rt_ma<3> vdd hvtpfet l=6e-08 w=1.43e-06 $X=40475 $Y=39677 $D=636
M3192 vdd 295 rt_ma<1> vdd hvtpfet l=6e-08 w=1.43e-06 $X=40475 $Y=41737 $D=636
M3193 vdd 296 rt_ca<3> vdd hvtpfet l=6e-08 w=1.43e-06 $X=40475 $Y=46137 $D=636
M3194 vdd 297 rt_ca<1> vdd hvtpfet l=6e-08 w=1.43e-06 $X=40475 $Y=48197 $D=636
M3195 vdd 549 543 vdd hvtpfet l=6e-08 w=2.06e-07 $X=40679 $Y=15321 $D=636
M3196 vdd 543 1363 vdd hvtpfet l=6e-08 w=2.74e-07 $X=40679 $Y=16069 $D=636
M3197 vdd 553 1364 vdd hvtpfet l=6e-08 w=2.74e-07 $X=40679 $Y=20589 $D=636
M3198 vdd 550 553 vdd hvtpfet l=6e-08 w=2.06e-07 $X=40679 $Y=21405 $D=636
M3199 vdd 551 542 vdd hvtpfet l=6e-08 w=2.06e-07 $X=40679 $Y=22241 $D=636
M3200 vdd 542 1365 vdd hvtpfet l=6e-08 w=2.74e-07 $X=40679 $Y=22989 $D=636
M3201 vdd 554 1366 vdd hvtpfet l=6e-08 w=2.74e-07 $X=40679 $Y=27509 $D=636
M3202 vdd 552 554 vdd hvtpfet l=6e-08 w=2.06e-07 $X=40679 $Y=28325 $D=636
M3203 vdd 303 r_saea_n vdd hvtpfet l=6e-08 w=1.43e-06 $X=40725 $Y=35277 $D=636
M3204 rb_ca<1> 289 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=40735 $Y=1506 $D=636
M3205 rb_ca<3> 290 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=40735 $Y=3566 $D=636
M3206 rb_ma<1> 291 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=40735 $Y=7966 $D=636
M3207 rb_ma<3> 292 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=40735 $Y=10026 $D=636
M3208 rt_ma<3> 294 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=40735 $Y=39677 $D=636
M3209 rt_ma<1> 295 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=40735 $Y=41737 $D=636
M3210 rt_ca<3> 296 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=40735 $Y=46137 $D=636
M3211 rt_ca<1> 297 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=40735 $Y=48197 $D=636
M3212 r_saea_n 303 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=40985 $Y=35277 $D=636
M3213 vdd 299 rb_ca<0> vdd hvtpfet l=6e-08 w=1.43e-06 $X=41245 $Y=1506 $D=636
M3214 vdd 300 rb_ca<2> vdd hvtpfet l=6e-08 w=1.43e-06 $X=41245 $Y=3566 $D=636
M3215 vdd 301 rb_ma<0> vdd hvtpfet l=6e-08 w=1.43e-06 $X=41245 $Y=7966 $D=636
M3216 vdd 302 rb_ma<2> vdd hvtpfet l=6e-08 w=1.43e-06 $X=41245 $Y=10026 $D=636
M3217 vdd 303 r_saea_n vdd hvtpfet l=6e-08 w=1.43e-06 $X=41245 $Y=35277 $D=636
M3218 vdd 304 rt_ma<2> vdd hvtpfet l=6e-08 w=1.43e-06 $X=41245 $Y=39677 $D=636
M3219 vdd 305 rt_ma<0> vdd hvtpfet l=6e-08 w=1.43e-06 $X=41245 $Y=41737 $D=636
M3220 vdd 306 rt_ca<2> vdd hvtpfet l=6e-08 w=1.43e-06 $X=41245 $Y=46137 $D=636
M3221 vdd 307 rt_ca<0> vdd hvtpfet l=6e-08 w=1.43e-06 $X=41245 $Y=48197 $D=636
M3222 vdd clka 287 vdd hvtpfet l=6e-08 w=2.1e-06 $X=41495 $Y=23621 $D=636
M3223 vdd 340 288 vdd hvtpfet l=6e-08 w=2.1e-06 $X=41495 $Y=26587 $D=636
M3224 rb_ca<0> 299 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=41505 $Y=1506 $D=636
M3225 rb_ca<2> 300 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=41505 $Y=3566 $D=636
M3226 rb_ma<0> 301 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=41505 $Y=7966 $D=636
M3227 rb_ma<2> 302 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=41505 $Y=10026 $D=636
M3228 285 497 vdd vdd hvtpfet l=6e-08 w=1.2e-06 $X=41505 $Y=15067 $D=636
M3229 286 498 vdd vdd hvtpfet l=6e-08 w=1.2e-06 $X=41505 $Y=18424 $D=636
M3230 r_saea_n 303 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=41505 $Y=35277 $D=636
M3231 rt_ma<2> 304 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=41505 $Y=39677 $D=636
M3232 rt_ma<0> 305 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=41505 $Y=41737 $D=636
M3233 rt_ca<2> 306 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=41505 $Y=46137 $D=636
M3234 rt_ca<0> 307 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=41505 $Y=48197 $D=636
M3235 r_clk_dqa 287 vdd vdd hvtpfet l=6e-08 w=2.1e-06 $X=41755 $Y=23621 $D=636
M3236 r_clk_dqa_n 288 vdd vdd hvtpfet l=6e-08 w=2.1e-06 $X=41755 $Y=26587 $D=636
M3237 vdd 299 rb_ca<0> vdd hvtpfet l=6e-08 w=1.43e-06 $X=41765 $Y=1506 $D=636
M3238 vdd 300 rb_ca<2> vdd hvtpfet l=6e-08 w=1.43e-06 $X=41765 $Y=3566 $D=636
M3239 vdd 301 rb_ma<0> vdd hvtpfet l=6e-08 w=1.43e-06 $X=41765 $Y=7966 $D=636
M3240 vdd 302 rb_ma<2> vdd hvtpfet l=6e-08 w=1.43e-06 $X=41765 $Y=10026 $D=636
M3241 vdd 303 r_saea_n vdd hvtpfet l=6e-08 w=1.43e-06 $X=41765 $Y=35277 $D=636
M3242 vdd 304 rt_ma<2> vdd hvtpfet l=6e-08 w=1.43e-06 $X=41765 $Y=39677 $D=636
M3243 vdd 305 rt_ma<0> vdd hvtpfet l=6e-08 w=1.43e-06 $X=41765 $Y=41737 $D=636
M3244 vdd 306 rt_ca<2> vdd hvtpfet l=6e-08 w=1.43e-06 $X=41765 $Y=46137 $D=636
M3245 vdd 307 rt_ca<0> vdd hvtpfet l=6e-08 w=1.43e-06 $X=41765 $Y=48197 $D=636
M3246 rb_tm_prea_n 285 vdd vdd hvtpfet l=6e-08 w=2.145e-06 $X=42015 $Y=14887 $D=636
M3247 rt_tm_prea_n 286 vdd vdd hvtpfet l=6e-08 w=2.145e-06 $X=42015 $Y=17659 $D=636
M3248 vdd 287 r_clk_dqa vdd hvtpfet l=6e-08 w=2.1e-06 $X=42015 $Y=23621 $D=636
M3249 vdd 288 r_clk_dqa_n vdd hvtpfet l=6e-08 w=2.1e-06 $X=42015 $Y=26587 $D=636
M3250 r_lwea 284 vdd vdd hvtpfet l=6e-08 w=2.145e-06 $X=42015 $Y=32504 $D=636
M3251 vdd 555 299 vdd hvtpfet l=6e-08 w=1.2e-06 $X=42275 $Y=1736 $D=636
M3252 vdd 556 300 vdd hvtpfet l=6e-08 w=1.2e-06 $X=42275 $Y=3566 $D=636
M3253 vdd 554 301 vdd hvtpfet l=6e-08 w=1.2e-06 $X=42275 $Y=8196 $D=636
M3254 vdd 553 302 vdd hvtpfet l=6e-08 w=1.2e-06 $X=42275 $Y=10026 $D=636
M3255 vdd 285 rb_tm_prea_n vdd hvtpfet l=6e-08 w=2.145e-06 $X=42275 $Y=14887 $D=636
M3256 vdd 286 rt_tm_prea_n vdd hvtpfet l=6e-08 w=2.145e-06 $X=42275 $Y=17659 $D=636
M3257 r_clk_dqa 287 vdd vdd hvtpfet l=6e-08 w=2.1e-06 $X=42275 $Y=23621 $D=636
M3258 r_clk_dqa_n 288 vdd vdd hvtpfet l=6e-08 w=2.1e-06 $X=42275 $Y=26587 $D=636
M3259 vdd 284 r_lwea vdd hvtpfet l=6e-08 w=2.145e-06 $X=42275 $Y=32504 $D=636
M3260 vdd 557 303 vdd hvtpfet l=6e-08 w=1.2e-06 $X=42275 $Y=35277 $D=636
M3261 vdd 553 304 vdd hvtpfet l=6e-08 w=1.2e-06 $X=42275 $Y=39907 $D=636
M3262 vdd 554 305 vdd hvtpfet l=6e-08 w=1.2e-06 $X=42275 $Y=41737 $D=636
M3263 vdd 558 306 vdd hvtpfet l=6e-08 w=1.2e-06 $X=42275 $Y=46367 $D=636
M3264 vdd 559 307 vdd hvtpfet l=6e-08 w=1.2e-06 $X=42275 $Y=48197 $D=636
M3265 303 557 vdd vdd hvtpfet l=6e-08 w=1.2e-06 $X=42535 $Y=35277 $D=636
.ends

************************************************************************
* Library Name: XMC55_DPS
* Cell Name:    xmc55_dps_localc16io_bw
************************************************************************
.SUBCKT xmc55_dps_localc16io_bw b_bla<15> b_bla<14> b_bla<13> b_bla<12> 
+ b_bla<11> b_bla<10> b_bla<9> b_bla<8> b_bla<7> b_bla<6> b_bla<5> b_bla<4> 
+ b_bla<3> b_bla<2> b_bla<1> b_bla<0> b_bla_n<15> b_bla_n<14> b_bla_n<13> 
+ b_bla_n<12> b_bla_n<11> b_bla_n<10> b_bla_n<9> b_bla_n<8> b_bla_n<7> 
+ b_bla_n<6> b_bla_n<5> b_bla_n<4> b_bla_n<3> b_bla_n<2> b_bla_n<1> b_bla_n<0> 
+ b_blb<15> b_blb<14> b_blb<13> b_blb<12> b_blb<11> b_blb<10> b_blb<9> 
+ b_blb<8> b_blb<7> b_blb<6> b_blb<5> b_blb<4> b_blb<3> b_blb<2> b_blb<1> 
+ b_blb<0> b_blb_n<15> b_blb_n<14> b_blb_n<13> b_blb_n<12> b_blb_n<11> 
+ b_blb_n<10> b_blb_n<9> b_blb_n<8> b_blb_n<7> b_blb_n<6> b_blb_n<5> 
+ b_blb_n<4> b_blb_n<3> b_blb_n<2> b_blb_n<1> b_blb_n<0> b_ca<3> b_ca<2> 
+ b_ca<1> b_ca<0> b_cb<3> b_cb<2> b_cb<1> b_cb<0> b_ma<3> b_ma<2> b_ma<1> 
+ b_ma<0> b_mb<3> b_mb<2> b_mb<1> b_mb<0> b_tm_prea_n b_tm_preb_n bwena bwenb 
+ clk_dqa clk_dqa_n clk_dqb clk_dqb_n da db ddqa ddqa_n ddqb ddqb_n lwea lweb 
+ qa qb sa_prea_n sa_preb_n saea_n saeb_n t_bla<15> t_bla<14> t_bla<13> 
+ t_bla<12> t_bla<11> t_bla<10> t_bla<9> t_bla<8> t_bla<7> t_bla<6> t_bla<5> 
+ t_bla<4> t_bla<3> t_bla<2> t_bla<1> t_bla<0> t_bla_n<15> t_bla_n<14> 
+ t_bla_n<13> t_bla_n<12> t_bla_n<11> t_bla_n<10> t_bla_n<9> t_bla_n<8> 
+ t_bla_n<7> t_bla_n<6> t_bla_n<5> t_bla_n<4> t_bla_n<3> t_bla_n<2> t_bla_n<1> 
+ t_bla_n<0> t_blb<15> t_blb<14> t_blb<13> t_blb<12> t_blb<11> t_blb<10> 
+ t_blb<9> t_blb<8> t_blb<7> t_blb<6> t_blb<5> t_blb<4> t_blb<3> t_blb<2> 
+ t_blb<1> t_blb<0> t_blb_n<15> t_blb_n<14> t_blb_n<13> t_blb_n<12> 
+ t_blb_n<11> t_blb_n<10> t_blb_n<9> t_blb_n<8> t_blb_n<7> t_blb_n<6> 
+ t_blb_n<5> t_blb_n<4> t_blb_n<3> t_blb_n<2> t_blb_n<1> t_blb_n<0> t_ca<3> 
+ t_ca<2> t_ca<1> t_ca<0> t_cb<3> t_cb<2> t_cb<1> t_cb<0> t_ma<3> t_ma<2> 
+ t_ma<1> t_ma<0> t_mb<3> t_mb<2> t_mb<1> t_mb<0> t_tm_prea_n t_tm_preb_n vdd 
+ vss
** N=20544 EP=186 IP=0 FDC=2568
M0 299 8 b_blb<15> vss hvtnfet l=6e-08 w=6e-07 $X=210 $Y=2941 $D=616
M1 299 8 b_blb<15> vss hvtnfet l=6e-08 w=6e-07 $X=210 $Y=3201 $D=616
M2 308 16 b_bla_n<15> vss hvtnfet l=6e-08 w=6e-07 $X=210 $Y=3881 $D=616
M3 308 16 b_bla_n<15> vss hvtnfet l=6e-08 w=6e-07 $X=210 $Y=4141 $D=616
M4 t_bla_n<15> 17 308 vss hvtnfet l=6e-08 w=6e-07 $X=210 $Y=46932 $D=616
M5 308 17 t_bla_n<15> vss hvtnfet l=6e-08 w=6e-07 $X=210 $Y=47192 $D=616
M6 t_blb<15> 9 299 vss hvtnfet l=6e-08 w=6e-07 $X=210 $Y=47872 $D=616
M7 299 9 t_blb<15> vss hvtnfet l=6e-08 w=6e-07 $X=210 $Y=48132 $D=616
M8 8 5 vss vss hvtnfet l=6e-08 w=4e-07 $X=535 $Y=4836 $D=616
M9 1025 b_cb<3> 5 vss hvtnfet l=6e-08 w=4e-07 $X=535 $Y=11331 $D=616
M10 1026 5 2 vss hvtnfet l=6e-08 w=4e-07 $X=535 $Y=12191 $D=616
M11 1027 6 3 vss hvtnfet l=6e-08 w=4e-07 $X=535 $Y=38542 $D=616
M12 1028 t_cb<3> 6 vss hvtnfet l=6e-08 w=4e-07 $X=535 $Y=39402 $D=616
M13 9 6 vss vss hvtnfet l=6e-08 w=4e-07 $X=535 $Y=45897 $D=616
M14 319 vdd vss vss hvtnfet l=6e-08 w=2.5e-07 $X=540 $Y=17720 $D=616
M15 vss vss vss vss hvtnfet l=7e-08 w=3.2e-07 $X=610 $Y=33798 $D=616
M16 vss vss vss vss hvtnfet l=1.4e-07 w=7.5e-07 $X=650 $Y=34593 $D=616
M17 vss 11 8 vss hvtnfet l=6e-08 w=4e-07 $X=795 $Y=4836 $D=616
M18 vss b_mb<3> 1025 vss hvtnfet l=6e-08 w=4e-07 $X=795 $Y=11331 $D=616
M19 vss 13 1026 vss hvtnfet l=6e-08 w=4e-07 $X=795 $Y=12191 $D=616
M20 vss 14 1027 vss hvtnfet l=6e-08 w=4e-07 $X=795 $Y=38542 $D=616
M21 vss t_mb<3> 1028 vss hvtnfet l=6e-08 w=4e-07 $X=795 $Y=39402 $D=616
M22 vss 11 9 vss hvtnfet l=6e-08 w=4e-07 $X=795 $Y=45897 $D=616
M23 vss vdd 319 vss hvtnfet l=6e-08 w=2.5e-07 $X=800 $Y=17720 $D=616
M24 vss vss vss vss hvtnfet l=6e-08 w=3e-07 $X=867 $Y=31223 $D=616
M25 vss vss vss vss hvtnfet l=8e-08 w=3.75e-07 $X=890 $Y=33798 $D=616
M26 302 vdd vss vss hvtnfet l=6e-08 w=2e-07 $X=975 $Y=21427 $D=616
M27 303 vdd vss vss hvtnfet l=6e-08 w=2e-07 $X=975 $Y=23694 $D=616
M28 304 vdd vss vss hvtnfet l=6e-08 w=2e-07 $X=975 $Y=24394 $D=616
M29 305 vdd vss vss hvtnfet l=6e-08 w=2e-07 $X=975 $Y=24904 $D=616
M30 vss vss vss vss hvtnfet l=1.4e-07 w=7.5e-07 $X=990 $Y=34593 $D=616
M31 318 vdd vss vss hvtnfet l=6e-08 w=6e-07 $X=1007 $Y=26159 $D=616
M32 16 20 vss vss hvtnfet l=6e-08 w=4e-07 $X=1055 $Y=4836 $D=616
M33 1029 b_ma<3> vss vss hvtnfet l=6e-08 w=4e-07 $X=1055 $Y=11331 $D=616
M34 1030 22 vss vss hvtnfet l=6e-08 w=4e-07 $X=1055 $Y=12191 $D=616
M35 1031 23 vss vss hvtnfet l=6e-08 w=4e-07 $X=1055 $Y=38542 $D=616
M36 1032 t_ma<3> vss vss hvtnfet l=6e-08 w=4e-07 $X=1055 $Y=39402 $D=616
M37 17 20 vss vss hvtnfet l=6e-08 w=4e-07 $X=1055 $Y=45897 $D=616
M38 319 vdd vss vss hvtnfet l=6e-08 w=2.5e-07 $X=1060 $Y=17720 $D=616
M39 317 8 b_blb_n<15> vss hvtnfet l=6e-08 w=6e-07 $X=1100 $Y=2941 $D=616
M40 317 8 b_blb_n<15> vss hvtnfet l=6e-08 w=6e-07 $X=1100 $Y=3201 $D=616
M41 b_bla<15> 16 328 vss hvtnfet l=6e-08 w=6e-07 $X=1100 $Y=3881 $D=616
M42 b_bla<15> 16 328 vss hvtnfet l=6e-08 w=6e-07 $X=1100 $Y=4141 $D=616
M43 328 17 t_bla<15> vss hvtnfet l=6e-08 w=6e-07 $X=1100 $Y=46932 $D=616
M44 t_bla<15> 17 328 vss hvtnfet l=6e-08 w=6e-07 $X=1100 $Y=47192 $D=616
M45 t_blb_n<15> 9 317 vss hvtnfet l=6e-08 w=6e-07 $X=1100 $Y=47872 $D=616
M46 317 9 t_blb_n<15> vss hvtnfet l=6e-08 w=6e-07 $X=1100 $Y=48132 $D=616
M47 vss vss vss vss hvtnfet l=6e-08 w=3e-07 $X=1127 $Y=31223 $D=616
M48 vss vss vss vss hvtnfet l=8e-08 w=3.75e-07 $X=1170 $Y=33798 $D=616
M49 vss vdd 318 vss hvtnfet l=6e-08 w=6e-07 $X=1267 $Y=26159 $D=616
M50 vss 18 16 vss hvtnfet l=6e-08 w=4e-07 $X=1315 $Y=4836 $D=616
M51 18 b_ca<3> 1029 vss hvtnfet l=6e-08 w=4e-07 $X=1315 $Y=11331 $D=616
M52 25 18 1030 vss hvtnfet l=6e-08 w=4e-07 $X=1315 $Y=12191 $D=616
M53 26 19 1031 vss hvtnfet l=6e-08 w=4e-07 $X=1315 $Y=38542 $D=616
M54 19 t_ca<3> 1032 vss hvtnfet l=6e-08 w=4e-07 $X=1315 $Y=39402 $D=616
M55 vss 19 17 vss hvtnfet l=6e-08 w=4e-07 $X=1315 $Y=45897 $D=616
M56 vss vdd 319 vss hvtnfet l=6e-08 w=2.5e-07 $X=1320 $Y=17720 $D=616
M57 vss vss vss vss hvtnfet l=1.4e-07 w=7.5e-07 $X=1330 $Y=34593 $D=616
M58 vss vss vss vss hvtnfet l=8e-08 w=3.75e-07 $X=1450 $Y=33798 $D=616
M59 vss vss vss vss hvtnfet l=1.4e-07 w=7.5e-07 $X=1670 $Y=34593 $D=616
M60 vss vss vss vss hvtnfet l=8e-08 w=3.75e-07 $X=1730 $Y=33798 $D=616
M61 343 vdd 346 vss hvtnfet l=6e-08 w=8e-07 $X=1787 $Y=26159 $D=616
M62 337 vdd vss vss hvtnfet l=1.4e-07 w=2.1e-07 $X=1805 $Y=14550 $D=616
M63 338 vdd vss vss hvtnfet l=1.4e-07 w=2.1e-07 $X=1805 $Y=16760 $D=616
M64 353 vdd vss vss hvtnfet l=6e-08 w=3e-07 $X=1830 $Y=17670 $D=616
M65 vss vss vss vss hvtnfet l=6e-08 w=3.2e-07 $X=1920 $Y=19812 $D=616
M66 vss vss vss vss hvtnfet l=6e-08 w=3.2e-07 $X=1920 $Y=20072 $D=616
M67 vss vss vss vss hvtnfet l=6e-08 w=3.2e-07 $X=1920 $Y=21162 $D=616
M68 vss vss vss vss hvtnfet l=6e-08 w=3.2e-07 $X=1920 $Y=21422 $D=616
M69 vss vss vss vss hvtnfet l=6e-08 w=3.2e-07 $X=1920 $Y=21682 $D=616
M70 vss vss vss vss hvtnfet l=6e-08 w=3.2e-07 $X=1920 $Y=21942 $D=616
M71 vss vss vss vss hvtnfet l=6e-08 w=3.2e-07 $X=1920 $Y=22762 $D=616
M72 vss vss vss vss hvtnfet l=6e-08 w=3.2e-07 $X=1920 $Y=23879 $D=616
M73 vss vss vss vss hvtnfet l=6e-08 w=3.2e-07 $X=1920 $Y=24139 $D=616
M74 vss vss vss vss hvtnfet l=6e-08 w=3.2e-07 $X=1920 $Y=24399 $D=616
M75 vss vss vss vss hvtnfet l=6e-08 w=3.2e-07 $X=1920 $Y=24659 $D=616
M76 vss vss vss vss hvtnfet l=8e-08 w=3.75e-07 $X=2010 $Y=33798 $D=616
M77 vss vss vss vss hvtnfet l=1.4e-07 w=7.5e-07 $X=2010 $Y=34593 $D=616
M78 vss vss vss vss hvtnfet l=6e-08 w=3e-07 $X=2037 $Y=31223 $D=616
M79 346 vdd 343 vss hvtnfet l=6e-08 w=8e-07 $X=2047 $Y=26159 $D=616
M80 vss vdd 353 vss hvtnfet l=6e-08 w=3e-07 $X=2090 $Y=17670 $D=616
M81 317 39 b_blb_n<14> vss hvtnfet l=6e-08 w=6e-07 $X=2120 $Y=2941 $D=616
M82 317 39 b_blb_n<14> vss hvtnfet l=6e-08 w=6e-07 $X=2120 $Y=3201 $D=616
M83 b_bla<14> 35 328 vss hvtnfet l=6e-08 w=6e-07 $X=2120 $Y=3881 $D=616
M84 b_bla<14> 35 328 vss hvtnfet l=6e-08 w=6e-07 $X=2120 $Y=4141 $D=616
M85 328 36 t_bla<14> vss hvtnfet l=6e-08 w=6e-07 $X=2120 $Y=46932 $D=616
M86 t_bla<14> 36 328 vss hvtnfet l=6e-08 w=6e-07 $X=2120 $Y=47192 $D=616
M87 t_blb_n<14> 40 317 vss hvtnfet l=6e-08 w=6e-07 $X=2120 $Y=47872 $D=616
M88 317 40 t_blb_n<14> vss hvtnfet l=6e-08 w=6e-07 $X=2120 $Y=48132 $D=616
M89 vss vdd 337 vss hvtnfet l=1.4e-07 w=2.1e-07 $X=2145 $Y=14550 $D=616
M90 vss vdd 338 vss hvtnfet l=1.4e-07 w=2.1e-07 $X=2145 $Y=16760 $D=616
M91 vss vss vss vss hvtnfet l=8e-08 w=3.75e-07 $X=2290 $Y=33798 $D=616
M92 vss vss vss vss hvtnfet l=6e-08 w=3e-07 $X=2297 $Y=31223 $D=616
M93 vss vdd 346 vss hvtnfet l=6e-08 w=8e-07 $X=2307 $Y=26159 $D=616
M94 353 vdd vss vss hvtnfet l=6e-08 w=3e-07 $X=2350 $Y=17670 $D=616
M95 vss vss vss vss hvtnfet l=1.4e-07 w=7.5e-07 $X=2350 $Y=34593 $D=616
M96 35 30 vss vss hvtnfet l=6e-08 w=4e-07 $X=2445 $Y=4836 $D=616
M97 1033 b_ca<2> 30 vss hvtnfet l=6e-08 w=4e-07 $X=2445 $Y=11331 $D=616
M98 1034 30 33 vss hvtnfet l=6e-08 w=4e-07 $X=2445 $Y=12191 $D=616
M99 1035 31 34 vss hvtnfet l=6e-08 w=4e-07 $X=2445 $Y=38542 $D=616
M100 1036 t_ca<2> 31 vss hvtnfet l=6e-08 w=4e-07 $X=2445 $Y=39402 $D=616
M101 36 31 vss vss hvtnfet l=6e-08 w=4e-07 $X=2445 $Y=45897 $D=616
M102 vss vss vss vss hvtnfet l=6e-08 w=3e-07 $X=2557 $Y=31223 $D=616
M103 346 vdd vss vss hvtnfet l=6e-08 w=8e-07 $X=2567 $Y=26159 $D=616
M104 vss vss vss vss hvtnfet l=8e-08 w=3.75e-07 $X=2570 $Y=33798 $D=616
M105 vss vdd 353 vss hvtnfet l=6e-08 w=3e-07 $X=2610 $Y=17670 $D=616
M106 vss vss vss vss hvtnfet l=1.4e-07 w=7.5e-07 $X=2690 $Y=34593 $D=616
M107 vss 20 35 vss hvtnfet l=6e-08 w=4e-07 $X=2705 $Y=4836 $D=616
M108 vss b_ma<3> 1033 vss hvtnfet l=6e-08 w=4e-07 $X=2705 $Y=11331 $D=616
M109 vss 22 1034 vss hvtnfet l=6e-08 w=4e-07 $X=2705 $Y=12191 $D=616
M110 vss 23 1035 vss hvtnfet l=6e-08 w=4e-07 $X=2705 $Y=38542 $D=616
M111 vss t_ma<3> 1036 vss hvtnfet l=6e-08 w=4e-07 $X=2705 $Y=39402 $D=616
M112 vss 20 36 vss hvtnfet l=6e-08 w=4e-07 $X=2705 $Y=45897 $D=616
M113 351 vdd vss vss hvtnfet l=1.4e-07 w=2.1e-07 $X=2735 $Y=14550 $D=616
M114 352 vdd vss vss hvtnfet l=1.4e-07 w=2.1e-07 $X=2735 $Y=16760 $D=616
M115 vss vss vss vss hvtnfet l=6e-08 w=3e-07 $X=2817 $Y=31223 $D=616
M116 vss vss vss vss hvtnfet l=8e-08 w=3.75e-07 $X=2850 $Y=33798 $D=616
M117 353 vdd vss vss hvtnfet l=6e-08 w=3e-07 $X=2870 $Y=17670 $D=616
M118 39 11 vss vss hvtnfet l=6e-08 w=4e-07 $X=2965 $Y=4836 $D=616
M119 1037 b_mb<3> vss vss hvtnfet l=6e-08 w=4e-07 $X=2965 $Y=11331 $D=616
M120 1038 13 vss vss hvtnfet l=6e-08 w=4e-07 $X=2965 $Y=12191 $D=616
M121 1039 14 vss vss hvtnfet l=6e-08 w=4e-07 $X=2965 $Y=38542 $D=616
M122 1040 t_mb<3> vss vss hvtnfet l=6e-08 w=4e-07 $X=2965 $Y=39402 $D=616
M123 40 11 vss vss hvtnfet l=6e-08 w=4e-07 $X=2965 $Y=45897 $D=616
M124 299 39 b_blb<14> vss hvtnfet l=6e-08 w=6e-07 $X=3010 $Y=2941 $D=616
M125 299 39 b_blb<14> vss hvtnfet l=6e-08 w=6e-07 $X=3010 $Y=3201 $D=616
M126 308 35 b_bla_n<14> vss hvtnfet l=6e-08 w=6e-07 $X=3010 $Y=3881 $D=616
M127 308 35 b_bla_n<14> vss hvtnfet l=6e-08 w=6e-07 $X=3010 $Y=4141 $D=616
M128 t_bla_n<14> 36 308 vss hvtnfet l=6e-08 w=6e-07 $X=3010 $Y=46932 $D=616
M129 308 36 t_bla_n<14> vss hvtnfet l=6e-08 w=6e-07 $X=3010 $Y=47192 $D=616
M130 t_blb<14> 40 299 vss hvtnfet l=6e-08 w=6e-07 $X=3010 $Y=47872 $D=616
M131 299 40 t_blb<14> vss hvtnfet l=6e-08 w=6e-07 $X=3010 $Y=48132 $D=616
M132 vss vss vss vss hvtnfet l=1.4e-07 w=7.5e-07 $X=3030 $Y=34593 $D=616
M133 vss vdd 351 vss hvtnfet l=1.4e-07 w=2.1e-07 $X=3075 $Y=14550 $D=616
M134 vss vdd 352 vss hvtnfet l=1.4e-07 w=2.1e-07 $X=3075 $Y=16760 $D=616
M135 360 vdd vss vss hvtnfet l=6e-08 w=6e-07 $X=3077 $Y=26159 $D=616
M136 vss vdd 353 vss hvtnfet l=6e-08 w=3e-07 $X=3130 $Y=17670 $D=616
M137 vss vss vss vss hvtnfet l=7e-08 w=3.2e-07 $X=3140 $Y=33798 $D=616
M138 vss 37 39 vss hvtnfet l=6e-08 w=4e-07 $X=3225 $Y=4836 $D=616
M139 37 b_cb<2> 1037 vss hvtnfet l=6e-08 w=4e-07 $X=3225 $Y=11331 $D=616
M140 41 37 1038 vss hvtnfet l=6e-08 w=4e-07 $X=3225 $Y=12191 $D=616
M141 42 38 1039 vss hvtnfet l=6e-08 w=4e-07 $X=3225 $Y=38542 $D=616
M142 38 t_cb<2> 1040 vss hvtnfet l=6e-08 w=4e-07 $X=3225 $Y=39402 $D=616
M143 vss 38 40 vss hvtnfet l=6e-08 w=4e-07 $X=3225 $Y=45897 $D=616
M144 vss vdd 360 vss hvtnfet l=6e-08 w=6e-07 $X=3337 $Y=26159 $D=616
M145 299 51 b_blb<13> vss hvtnfet l=6e-08 w=6e-07 $X=4030 $Y=2941 $D=616
M146 299 51 b_blb<13> vss hvtnfet l=6e-08 w=6e-07 $X=4030 $Y=3201 $D=616
M147 308 53 b_bla_n<13> vss hvtnfet l=6e-08 w=6e-07 $X=4030 $Y=3881 $D=616
M148 308 53 b_bla_n<13> vss hvtnfet l=6e-08 w=6e-07 $X=4030 $Y=4141 $D=616
M149 t_bla_n<13> 54 308 vss hvtnfet l=6e-08 w=6e-07 $X=4030 $Y=46932 $D=616
M150 308 54 t_bla_n<13> vss hvtnfet l=6e-08 w=6e-07 $X=4030 $Y=47192 $D=616
M151 t_blb<13> 52 299 vss hvtnfet l=6e-08 w=6e-07 $X=4030 $Y=47872 $D=616
M152 299 52 t_blb<13> vss hvtnfet l=6e-08 w=6e-07 $X=4030 $Y=48132 $D=616
M153 373 vdd vss vss hvtnfet l=6e-08 w=6e-07 $X=4243 $Y=26159 $D=616
M154 51 48 vss vss hvtnfet l=6e-08 w=4e-07 $X=4355 $Y=4836 $D=616
M155 1041 b_cb<1> 48 vss hvtnfet l=6e-08 w=4e-07 $X=4355 $Y=11331 $D=616
M156 1042 48 45 vss hvtnfet l=6e-08 w=4e-07 $X=4355 $Y=12191 $D=616
M157 1043 49 46 vss hvtnfet l=6e-08 w=4e-07 $X=4355 $Y=38542 $D=616
M158 1044 t_cb<1> 49 vss hvtnfet l=6e-08 w=4e-07 $X=4355 $Y=39402 $D=616
M159 52 49 vss vss hvtnfet l=6e-08 w=4e-07 $X=4355 $Y=45897 $D=616
M160 376 vdd vss vss hvtnfet l=1.4e-07 w=2.1e-07 $X=4425 $Y=14550 $D=616
M161 377 vdd vss vss hvtnfet l=1.4e-07 w=2.1e-07 $X=4425 $Y=16760 $D=616
M162 vss vss vss vss hvtnfet l=7e-08 w=3.2e-07 $X=4430 $Y=33798 $D=616
M163 394 vdd vss vss hvtnfet l=6e-08 w=3e-07 $X=4450 $Y=17670 $D=616
M164 vss vss vss vss hvtnfet l=1.4e-07 w=7.5e-07 $X=4470 $Y=34593 $D=616
M165 vss vdd 373 vss hvtnfet l=6e-08 w=6e-07 $X=4503 $Y=26159 $D=616
M166 vss 11 51 vss hvtnfet l=6e-08 w=4e-07 $X=4615 $Y=4836 $D=616
M167 vss b_mb<3> 1041 vss hvtnfet l=6e-08 w=4e-07 $X=4615 $Y=11331 $D=616
M168 vss 13 1042 vss hvtnfet l=6e-08 w=4e-07 $X=4615 $Y=12191 $D=616
M169 vss 14 1043 vss hvtnfet l=6e-08 w=4e-07 $X=4615 $Y=38542 $D=616
M170 vss t_mb<3> 1044 vss hvtnfet l=6e-08 w=4e-07 $X=4615 $Y=39402 $D=616
M171 vss 11 52 vss hvtnfet l=6e-08 w=4e-07 $X=4615 $Y=45897 $D=616
M172 vss vdd 394 vss hvtnfet l=6e-08 w=3e-07 $X=4710 $Y=17670 $D=616
M173 vss vss vss vss hvtnfet l=8e-08 w=3.75e-07 $X=4710 $Y=33798 $D=616
M174 vss vss vss vss hvtnfet l=6e-08 w=3e-07 $X=4763 $Y=31223 $D=616
M175 vss vdd 376 vss hvtnfet l=1.4e-07 w=2.1e-07 $X=4765 $Y=14550 $D=616
M176 vss vdd 377 vss hvtnfet l=1.4e-07 w=2.1e-07 $X=4765 $Y=16760 $D=616
M177 vss vss vss vss hvtnfet l=1.4e-07 w=7.5e-07 $X=4810 $Y=34593 $D=616
M178 53 20 vss vss hvtnfet l=6e-08 w=4e-07 $X=4875 $Y=4836 $D=616
M179 1045 b_ma<3> vss vss hvtnfet l=6e-08 w=4e-07 $X=4875 $Y=11331 $D=616
M180 1046 22 vss vss hvtnfet l=6e-08 w=4e-07 $X=4875 $Y=12191 $D=616
M181 1047 23 vss vss hvtnfet l=6e-08 w=4e-07 $X=4875 $Y=38542 $D=616
M182 1048 t_ma<3> vss vss hvtnfet l=6e-08 w=4e-07 $X=4875 $Y=39402 $D=616
M183 54 20 vss vss hvtnfet l=6e-08 w=4e-07 $X=4875 $Y=45897 $D=616
M184 317 51 b_blb_n<13> vss hvtnfet l=6e-08 w=6e-07 $X=4920 $Y=2941 $D=616
M185 317 51 b_blb_n<13> vss hvtnfet l=6e-08 w=6e-07 $X=4920 $Y=3201 $D=616
M186 b_bla<13> 53 328 vss hvtnfet l=6e-08 w=6e-07 $X=4920 $Y=3881 $D=616
M187 b_bla<13> 53 328 vss hvtnfet l=6e-08 w=6e-07 $X=4920 $Y=4141 $D=616
M188 328 54 t_bla<13> vss hvtnfet l=6e-08 w=6e-07 $X=4920 $Y=46932 $D=616
M189 t_bla<13> 54 328 vss hvtnfet l=6e-08 w=6e-07 $X=4920 $Y=47192 $D=616
M190 t_blb_n<13> 52 317 vss hvtnfet l=6e-08 w=6e-07 $X=4920 $Y=47872 $D=616
M191 317 52 t_blb_n<13> vss hvtnfet l=6e-08 w=6e-07 $X=4920 $Y=48132 $D=616
M192 394 vdd vss vss hvtnfet l=6e-08 w=3e-07 $X=4970 $Y=17670 $D=616
M193 vss vss vss vss hvtnfet l=8e-08 w=3.75e-07 $X=4990 $Y=33798 $D=616
M194 vss vdd 400 vss hvtnfet l=6e-08 w=8e-07 $X=5013 $Y=26159 $D=616
M195 vss vss vss vss hvtnfet l=6e-08 w=3e-07 $X=5023 $Y=31223 $D=616
M196 vss 55 53 vss hvtnfet l=6e-08 w=4e-07 $X=5135 $Y=4836 $D=616
M197 55 b_ca<1> 1045 vss hvtnfet l=6e-08 w=4e-07 $X=5135 $Y=11331 $D=616
M198 57 55 1046 vss hvtnfet l=6e-08 w=4e-07 $X=5135 $Y=12191 $D=616
M199 58 56 1047 vss hvtnfet l=6e-08 w=4e-07 $X=5135 $Y=38542 $D=616
M200 56 t_ca<1> 1048 vss hvtnfet l=6e-08 w=4e-07 $X=5135 $Y=39402 $D=616
M201 vss 56 54 vss hvtnfet l=6e-08 w=4e-07 $X=5135 $Y=45897 $D=616
M202 vss vss vss vss hvtnfet l=1.4e-07 w=7.5e-07 $X=5150 $Y=34593 $D=616
M203 vss vdd 394 vss hvtnfet l=6e-08 w=3e-07 $X=5230 $Y=17670 $D=616
M204 vss vss vss vss hvtnfet l=8e-08 w=3.75e-07 $X=5270 $Y=33798 $D=616
M205 400 vdd vss vss hvtnfet l=6e-08 w=8e-07 $X=5273 $Y=26159 $D=616
M206 vss vss vss vss hvtnfet l=6e-08 w=3e-07 $X=5283 $Y=31223 $D=616
M207 392 vdd vss vss hvtnfet l=1.4e-07 w=2.1e-07 $X=5355 $Y=14550 $D=616
M208 393 vdd vss vss hvtnfet l=1.4e-07 w=2.1e-07 $X=5355 $Y=16760 $D=616
M209 vss vss vss vss hvtnfet l=6e-08 w=3.2e-07 $X=5400 $Y=19812 $D=616
M210 vss vss vss vss hvtnfet l=6e-08 w=3.2e-07 $X=5400 $Y=20072 $D=616
M211 vss vss vss vss hvtnfet l=6e-08 w=3.2e-07 $X=5400 $Y=21162 $D=616
M212 vss vss vss vss hvtnfet l=6e-08 w=3.2e-07 $X=5400 $Y=21422 $D=616
M213 vss vss vss vss hvtnfet l=6e-08 w=3.2e-07 $X=5400 $Y=21682 $D=616
M214 vss vss vss vss hvtnfet l=6e-08 w=3.2e-07 $X=5400 $Y=21942 $D=616
M215 vss vss vss vss hvtnfet l=6e-08 w=3.2e-07 $X=5400 $Y=22762 $D=616
M216 vss vss vss vss hvtnfet l=6e-08 w=3.2e-07 $X=5400 $Y=23879 $D=616
M217 vss vss vss vss hvtnfet l=6e-08 w=3.2e-07 $X=5400 $Y=24139 $D=616
M218 vss vss vss vss hvtnfet l=6e-08 w=3.2e-07 $X=5400 $Y=24399 $D=616
M219 vss vss vss vss hvtnfet l=6e-08 w=3.2e-07 $X=5400 $Y=24659 $D=616
M220 394 vdd vss vss hvtnfet l=6e-08 w=3e-07 $X=5490 $Y=17670 $D=616
M221 vss vss vss vss hvtnfet l=1.4e-07 w=7.5e-07 $X=5490 $Y=34593 $D=616
M222 395 vdd 400 vss hvtnfet l=6e-08 w=8e-07 $X=5533 $Y=26159 $D=616
M223 vss vss vss vss hvtnfet l=6e-08 w=3e-07 $X=5543 $Y=31223 $D=616
M224 vss vss vss vss hvtnfet l=8e-08 w=3.75e-07 $X=5550 $Y=33798 $D=616
M225 vss vdd 392 vss hvtnfet l=1.4e-07 w=2.1e-07 $X=5695 $Y=14550 $D=616
M226 vss vdd 393 vss hvtnfet l=1.4e-07 w=2.1e-07 $X=5695 $Y=16760 $D=616
M227 vss vdd 394 vss hvtnfet l=6e-08 w=3e-07 $X=5750 $Y=17670 $D=616
M228 400 vdd 395 vss hvtnfet l=6e-08 w=8e-07 $X=5793 $Y=26159 $D=616
M229 vss vss vss vss hvtnfet l=8e-08 w=3.75e-07 $X=5830 $Y=33798 $D=616
M230 vss vss vss vss hvtnfet l=1.4e-07 w=7.5e-07 $X=5830 $Y=34593 $D=616
M231 317 71 b_blb_n<12> vss hvtnfet l=6e-08 w=6e-07 $X=5940 $Y=2941 $D=616
M232 317 71 b_blb_n<12> vss hvtnfet l=6e-08 w=6e-07 $X=5940 $Y=3201 $D=616
M233 b_bla<12> 67 328 vss hvtnfet l=6e-08 w=6e-07 $X=5940 $Y=3881 $D=616
M234 b_bla<12> 67 328 vss hvtnfet l=6e-08 w=6e-07 $X=5940 $Y=4141 $D=616
M235 328 68 t_bla<12> vss hvtnfet l=6e-08 w=6e-07 $X=5940 $Y=46932 $D=616
M236 t_bla<12> 68 328 vss hvtnfet l=6e-08 w=6e-07 $X=5940 $Y=47192 $D=616
M237 t_blb_n<12> 72 317 vss hvtnfet l=6e-08 w=6e-07 $X=5940 $Y=47872 $D=616
M238 317 72 t_blb_n<12> vss hvtnfet l=6e-08 w=6e-07 $X=5940 $Y=48132 $D=616
M239 vss vss vss vss hvtnfet l=8e-08 w=3.75e-07 $X=6110 $Y=33798 $D=616
M240 vss vss vss vss hvtnfet l=1.4e-07 w=7.5e-07 $X=6170 $Y=34593 $D=616
M241 418 vdd vss vss hvtnfet l=6e-08 w=2.5e-07 $X=6260 $Y=17720 $D=616
M242 67 62 vss vss hvtnfet l=6e-08 w=4e-07 $X=6265 $Y=4836 $D=616
M243 1049 b_ca<0> 62 vss hvtnfet l=6e-08 w=4e-07 $X=6265 $Y=11331 $D=616
M244 1050 62 65 vss hvtnfet l=6e-08 w=4e-07 $X=6265 $Y=12191 $D=616
M245 1051 63 66 vss hvtnfet l=6e-08 w=4e-07 $X=6265 $Y=38542 $D=616
M246 1052 t_ca<0> 63 vss hvtnfet l=6e-08 w=4e-07 $X=6265 $Y=39402 $D=616
M247 68 63 vss vss hvtnfet l=6e-08 w=4e-07 $X=6265 $Y=45897 $D=616
M248 407 vdd vss vss hvtnfet l=6e-08 w=6e-07 $X=6313 $Y=26159 $D=616
M249 vss vss vss vss hvtnfet l=8e-08 w=3.75e-07 $X=6390 $Y=33798 $D=616
M250 vss vss vss vss hvtnfet l=6e-08 w=3e-07 $X=6453 $Y=31223 $D=616
M251 408 vdd vss vss hvtnfet l=6e-08 w=2e-07 $X=6465 $Y=21427 $D=616
M252 409 vdd vss vss hvtnfet l=6e-08 w=2e-07 $X=6465 $Y=23694 $D=616
M253 410 vdd vss vss hvtnfet l=6e-08 w=2e-07 $X=6465 $Y=24394 $D=616
M254 411 vdd vss vss hvtnfet l=6e-08 w=2e-07 $X=6465 $Y=24904 $D=616
M255 vss vss vss vss hvtnfet l=1.4e-07 w=7.5e-07 $X=6510 $Y=34593 $D=616
M256 vss vdd 418 vss hvtnfet l=6e-08 w=2.5e-07 $X=6520 $Y=17720 $D=616
M257 vss 20 67 vss hvtnfet l=6e-08 w=4e-07 $X=6525 $Y=4836 $D=616
M258 vss b_ma<3> 1049 vss hvtnfet l=6e-08 w=4e-07 $X=6525 $Y=11331 $D=616
M259 vss 22 1050 vss hvtnfet l=6e-08 w=4e-07 $X=6525 $Y=12191 $D=616
M260 vss 23 1051 vss hvtnfet l=6e-08 w=4e-07 $X=6525 $Y=38542 $D=616
M261 vss t_ma<3> 1052 vss hvtnfet l=6e-08 w=4e-07 $X=6525 $Y=39402 $D=616
M262 vss 20 68 vss hvtnfet l=6e-08 w=4e-07 $X=6525 $Y=45897 $D=616
M263 vss vdd 407 vss hvtnfet l=6e-08 w=6e-07 $X=6573 $Y=26159 $D=616
M264 vss vss vss vss hvtnfet l=8e-08 w=3.75e-07 $X=6670 $Y=33798 $D=616
M265 vss vss vss vss hvtnfet l=6e-08 w=3e-07 $X=6713 $Y=31223 $D=616
M266 418 vdd vss vss hvtnfet l=6e-08 w=2.5e-07 $X=6780 $Y=17720 $D=616
M267 71 11 vss vss hvtnfet l=6e-08 w=4e-07 $X=6785 $Y=4836 $D=616
M268 1053 b_mb<3> vss vss hvtnfet l=6e-08 w=4e-07 $X=6785 $Y=11331 $D=616
M269 1054 13 vss vss hvtnfet l=6e-08 w=4e-07 $X=6785 $Y=12191 $D=616
M270 1055 14 vss vss hvtnfet l=6e-08 w=4e-07 $X=6785 $Y=38542 $D=616
M271 1056 t_mb<3> vss vss hvtnfet l=6e-08 w=4e-07 $X=6785 $Y=39402 $D=616
M272 72 11 vss vss hvtnfet l=6e-08 w=4e-07 $X=6785 $Y=45897 $D=616
M273 299 71 b_blb<12> vss hvtnfet l=6e-08 w=6e-07 $X=6830 $Y=2941 $D=616
M274 299 71 b_blb<12> vss hvtnfet l=6e-08 w=6e-07 $X=6830 $Y=3201 $D=616
M275 308 67 b_bla_n<12> vss hvtnfet l=6e-08 w=6e-07 $X=6830 $Y=3881 $D=616
M276 308 67 b_bla_n<12> vss hvtnfet l=6e-08 w=6e-07 $X=6830 $Y=4141 $D=616
M277 t_bla_n<12> 68 308 vss hvtnfet l=6e-08 w=6e-07 $X=6830 $Y=46932 $D=616
M278 308 68 t_bla_n<12> vss hvtnfet l=6e-08 w=6e-07 $X=6830 $Y=47192 $D=616
M279 t_blb<12> 72 299 vss hvtnfet l=6e-08 w=6e-07 $X=6830 $Y=47872 $D=616
M280 299 72 t_blb<12> vss hvtnfet l=6e-08 w=6e-07 $X=6830 $Y=48132 $D=616
M281 vss vss vss vss hvtnfet l=1.4e-07 w=7.5e-07 $X=6850 $Y=34593 $D=616
M282 vss vss vss vss hvtnfet l=7e-08 w=3.2e-07 $X=6960 $Y=33798 $D=616
M283 vss vdd 418 vss hvtnfet l=6e-08 w=2.5e-07 $X=7040 $Y=17720 $D=616
M284 vss 69 71 vss hvtnfet l=6e-08 w=4e-07 $X=7045 $Y=4836 $D=616
M285 69 b_cb<0> 1053 vss hvtnfet l=6e-08 w=4e-07 $X=7045 $Y=11331 $D=616
M286 73 69 1054 vss hvtnfet l=6e-08 w=4e-07 $X=7045 $Y=12191 $D=616
M287 74 70 1055 vss hvtnfet l=6e-08 w=4e-07 $X=7045 $Y=38542 $D=616
M288 70 t_cb<0> 1056 vss hvtnfet l=6e-08 w=4e-07 $X=7045 $Y=39402 $D=616
M289 vss 70 72 vss hvtnfet l=6e-08 w=4e-07 $X=7045 $Y=45897 $D=616
M290 299 81 b_blb<11> vss hvtnfet l=6e-08 w=6e-07 $X=7850 $Y=2941 $D=616
M291 299 81 b_blb<11> vss hvtnfet l=6e-08 w=6e-07 $X=7850 $Y=3201 $D=616
M292 308 85 b_bla_n<11> vss hvtnfet l=6e-08 w=6e-07 $X=7850 $Y=3881 $D=616
M293 308 85 b_bla_n<11> vss hvtnfet l=6e-08 w=6e-07 $X=7850 $Y=4141 $D=616
M294 t_bla_n<11> 86 308 vss hvtnfet l=6e-08 w=6e-07 $X=7850 $Y=46932 $D=616
M295 308 86 t_bla_n<11> vss hvtnfet l=6e-08 w=6e-07 $X=7850 $Y=47192 $D=616
M296 t_blb<11> 82 299 vss hvtnfet l=6e-08 w=6e-07 $X=7850 $Y=47872 $D=616
M297 299 82 t_blb<11> vss hvtnfet l=6e-08 w=6e-07 $X=7850 $Y=48132 $D=616
M298 81 79 vss vss hvtnfet l=6e-08 w=4e-07 $X=8175 $Y=4836 $D=616
M299 1057 b_cb<3> 79 vss hvtnfet l=6e-08 w=4e-07 $X=8175 $Y=11331 $D=616
M300 1058 79 77 vss hvtnfet l=6e-08 w=4e-07 $X=8175 $Y=12191 $D=616
M301 1059 80 78 vss hvtnfet l=6e-08 w=4e-07 $X=8175 $Y=38542 $D=616
M302 1060 t_cb<3> 80 vss hvtnfet l=6e-08 w=4e-07 $X=8175 $Y=39402 $D=616
M303 82 80 vss vss hvtnfet l=6e-08 w=4e-07 $X=8175 $Y=45897 $D=616
M304 446 vdd vss vss hvtnfet l=6e-08 w=2.5e-07 $X=8180 $Y=17720 $D=616
M305 vss vss vss vss hvtnfet l=7e-08 w=3.2e-07 $X=8250 $Y=33798 $D=616
M306 vss vss vss vss hvtnfet l=1.4e-07 w=7.5e-07 $X=8290 $Y=34593 $D=616
M307 vss 11 81 vss hvtnfet l=6e-08 w=4e-07 $X=8435 $Y=4836 $D=616
M308 vss b_mb<2> 1057 vss hvtnfet l=6e-08 w=4e-07 $X=8435 $Y=11331 $D=616
M309 vss 13 1058 vss hvtnfet l=6e-08 w=4e-07 $X=8435 $Y=12191 $D=616
M310 vss 14 1059 vss hvtnfet l=6e-08 w=4e-07 $X=8435 $Y=38542 $D=616
M311 vss t_mb<2> 1060 vss hvtnfet l=6e-08 w=4e-07 $X=8435 $Y=39402 $D=616
M312 vss 11 82 vss hvtnfet l=6e-08 w=4e-07 $X=8435 $Y=45897 $D=616
M313 vss vdd 446 vss hvtnfet l=6e-08 w=2.5e-07 $X=8440 $Y=17720 $D=616
M314 vss vss vss vss hvtnfet l=6e-08 w=3e-07 $X=8507 $Y=31223 $D=616
M315 vss vss vss vss hvtnfet l=8e-08 w=3.75e-07 $X=8530 $Y=33798 $D=616
M316 431 vdd vss vss hvtnfet l=6e-08 w=2e-07 $X=8615 $Y=21427 $D=616
M317 432 vdd vss vss hvtnfet l=6e-08 w=2e-07 $X=8615 $Y=23694 $D=616
M318 433 vdd vss vss hvtnfet l=6e-08 w=2e-07 $X=8615 $Y=24394 $D=616
M319 434 vdd vss vss hvtnfet l=6e-08 w=2e-07 $X=8615 $Y=24904 $D=616
M320 vss vss vss vss hvtnfet l=1.4e-07 w=7.5e-07 $X=8630 $Y=34593 $D=616
M321 445 vdd vss vss hvtnfet l=6e-08 w=6e-07 $X=8647 $Y=26159 $D=616
M322 85 20 vss vss hvtnfet l=6e-08 w=4e-07 $X=8695 $Y=4836 $D=616
M323 1061 b_ma<2> vss vss hvtnfet l=6e-08 w=4e-07 $X=8695 $Y=11331 $D=616
M324 1062 22 vss vss hvtnfet l=6e-08 w=4e-07 $X=8695 $Y=12191 $D=616
M325 1063 23 vss vss hvtnfet l=6e-08 w=4e-07 $X=8695 $Y=38542 $D=616
M326 1064 t_ma<2> vss vss hvtnfet l=6e-08 w=4e-07 $X=8695 $Y=39402 $D=616
M327 86 20 vss vss hvtnfet l=6e-08 w=4e-07 $X=8695 $Y=45897 $D=616
M328 446 vdd vss vss hvtnfet l=6e-08 w=2.5e-07 $X=8700 $Y=17720 $D=616
M329 317 81 b_blb_n<11> vss hvtnfet l=6e-08 w=6e-07 $X=8740 $Y=2941 $D=616
M330 317 81 b_blb_n<11> vss hvtnfet l=6e-08 w=6e-07 $X=8740 $Y=3201 $D=616
M331 b_bla<11> 85 328 vss hvtnfet l=6e-08 w=6e-07 $X=8740 $Y=3881 $D=616
M332 b_bla<11> 85 328 vss hvtnfet l=6e-08 w=6e-07 $X=8740 $Y=4141 $D=616
M333 328 86 t_bla<11> vss hvtnfet l=6e-08 w=6e-07 $X=8740 $Y=46932 $D=616
M334 t_bla<11> 86 328 vss hvtnfet l=6e-08 w=6e-07 $X=8740 $Y=47192 $D=616
M335 t_blb_n<11> 82 317 vss hvtnfet l=6e-08 w=6e-07 $X=8740 $Y=47872 $D=616
M336 317 82 t_blb_n<11> vss hvtnfet l=6e-08 w=6e-07 $X=8740 $Y=48132 $D=616
M337 vss vss vss vss hvtnfet l=6e-08 w=3e-07 $X=8767 $Y=31223 $D=616
M338 vss vss vss vss hvtnfet l=8e-08 w=3.75e-07 $X=8810 $Y=33798 $D=616
M339 vss vdd 445 vss hvtnfet l=6e-08 w=6e-07 $X=8907 $Y=26159 $D=616
M340 vss 87 85 vss hvtnfet l=6e-08 w=4e-07 $X=8955 $Y=4836 $D=616
M341 87 b_ca<3> 1061 vss hvtnfet l=6e-08 w=4e-07 $X=8955 $Y=11331 $D=616
M342 91 87 1062 vss hvtnfet l=6e-08 w=4e-07 $X=8955 $Y=12191 $D=616
M343 92 88 1063 vss hvtnfet l=6e-08 w=4e-07 $X=8955 $Y=38542 $D=616
M344 88 t_ca<3> 1064 vss hvtnfet l=6e-08 w=4e-07 $X=8955 $Y=39402 $D=616
M345 vss 88 86 vss hvtnfet l=6e-08 w=4e-07 $X=8955 $Y=45897 $D=616
M346 vss vdd 446 vss hvtnfet l=6e-08 w=2.5e-07 $X=8960 $Y=17720 $D=616
M347 vss vss vss vss hvtnfet l=1.4e-07 w=7.5e-07 $X=8970 $Y=34593 $D=616
M348 vss vss vss vss hvtnfet l=8e-08 w=3.75e-07 $X=9090 $Y=33798 $D=616
M349 vss vss vss vss hvtnfet l=1.4e-07 w=7.5e-07 $X=9310 $Y=34593 $D=616
M350 vss vss vss vss hvtnfet l=8e-08 w=3.75e-07 $X=9370 $Y=33798 $D=616
M351 467 vdd 470 vss hvtnfet l=6e-08 w=8e-07 $X=9427 $Y=26159 $D=616
M352 461 vdd vss vss hvtnfet l=1.4e-07 w=2.1e-07 $X=9445 $Y=14550 $D=616
M353 462 vdd vss vss hvtnfet l=1.4e-07 w=2.1e-07 $X=9445 $Y=16760 $D=616
M354 477 vdd vss vss hvtnfet l=6e-08 w=3e-07 $X=9470 $Y=17670 $D=616
M355 vss vss vss vss hvtnfet l=6e-08 w=3.2e-07 $X=9560 $Y=19812 $D=616
M356 vss vss vss vss hvtnfet l=6e-08 w=3.2e-07 $X=9560 $Y=20072 $D=616
M357 vss vss vss vss hvtnfet l=6e-08 w=3.2e-07 $X=9560 $Y=21162 $D=616
M358 vss vss vss vss hvtnfet l=6e-08 w=3.2e-07 $X=9560 $Y=21422 $D=616
M359 vss vss vss vss hvtnfet l=6e-08 w=3.2e-07 $X=9560 $Y=21682 $D=616
M360 vss vss vss vss hvtnfet l=6e-08 w=3.2e-07 $X=9560 $Y=21942 $D=616
M361 vss vss vss vss hvtnfet l=6e-08 w=3.2e-07 $X=9560 $Y=22762 $D=616
M362 vss vss vss vss hvtnfet l=6e-08 w=3.2e-07 $X=9560 $Y=23879 $D=616
M363 vss vss vss vss hvtnfet l=6e-08 w=3.2e-07 $X=9560 $Y=24139 $D=616
M364 vss vss vss vss hvtnfet l=6e-08 w=3.2e-07 $X=9560 $Y=24399 $D=616
M365 vss vss vss vss hvtnfet l=6e-08 w=3.2e-07 $X=9560 $Y=24659 $D=616
M366 vss vss vss vss hvtnfet l=8e-08 w=3.75e-07 $X=9650 $Y=33798 $D=616
M367 vss vss vss vss hvtnfet l=1.4e-07 w=7.5e-07 $X=9650 $Y=34593 $D=616
M368 vss vss vss vss hvtnfet l=6e-08 w=3e-07 $X=9677 $Y=31223 $D=616
M369 470 vdd 467 vss hvtnfet l=6e-08 w=8e-07 $X=9687 $Y=26159 $D=616
M370 vss vdd 477 vss hvtnfet l=6e-08 w=3e-07 $X=9730 $Y=17670 $D=616
M371 317 101 b_blb_n<10> vss hvtnfet l=6e-08 w=6e-07 $X=9760 $Y=2941 $D=616
M372 317 101 b_blb_n<10> vss hvtnfet l=6e-08 w=6e-07 $X=9760 $Y=3201 $D=616
M373 b_bla<10> 97 328 vss hvtnfet l=6e-08 w=6e-07 $X=9760 $Y=3881 $D=616
M374 b_bla<10> 97 328 vss hvtnfet l=6e-08 w=6e-07 $X=9760 $Y=4141 $D=616
M375 328 98 t_bla<10> vss hvtnfet l=6e-08 w=6e-07 $X=9760 $Y=46932 $D=616
M376 t_bla<10> 98 328 vss hvtnfet l=6e-08 w=6e-07 $X=9760 $Y=47192 $D=616
M377 t_blb_n<10> 102 317 vss hvtnfet l=6e-08 w=6e-07 $X=9760 $Y=47872 $D=616
M378 317 102 t_blb_n<10> vss hvtnfet l=6e-08 w=6e-07 $X=9760 $Y=48132 $D=616
M379 vss vdd 461 vss hvtnfet l=1.4e-07 w=2.1e-07 $X=9785 $Y=14550 $D=616
M380 vss vdd 462 vss hvtnfet l=1.4e-07 w=2.1e-07 $X=9785 $Y=16760 $D=616
M381 vss vss vss vss hvtnfet l=8e-08 w=3.75e-07 $X=9930 $Y=33798 $D=616
M382 vss vss vss vss hvtnfet l=6e-08 w=3e-07 $X=9937 $Y=31223 $D=616
M383 vss vdd 470 vss hvtnfet l=6e-08 w=8e-07 $X=9947 $Y=26159 $D=616
M384 477 vdd vss vss hvtnfet l=6e-08 w=3e-07 $X=9990 $Y=17670 $D=616
M385 vss vss vss vss hvtnfet l=1.4e-07 w=7.5e-07 $X=9990 $Y=34593 $D=616
M386 97 93 vss vss hvtnfet l=6e-08 w=4e-07 $X=10085 $Y=4836 $D=616
M387 1065 b_ca<2> 93 vss hvtnfet l=6e-08 w=4e-07 $X=10085 $Y=11331 $D=616
M388 1066 93 95 vss hvtnfet l=6e-08 w=4e-07 $X=10085 $Y=12191 $D=616
M389 1067 94 96 vss hvtnfet l=6e-08 w=4e-07 $X=10085 $Y=38542 $D=616
M390 1068 t_ca<2> 94 vss hvtnfet l=6e-08 w=4e-07 $X=10085 $Y=39402 $D=616
M391 98 94 vss vss hvtnfet l=6e-08 w=4e-07 $X=10085 $Y=45897 $D=616
M392 vss vss vss vss hvtnfet l=6e-08 w=3e-07 $X=10197 $Y=31223 $D=616
M393 470 vdd vss vss hvtnfet l=6e-08 w=8e-07 $X=10207 $Y=26159 $D=616
M394 vss vss vss vss hvtnfet l=8e-08 w=3.75e-07 $X=10210 $Y=33798 $D=616
M395 vss vdd 477 vss hvtnfet l=6e-08 w=3e-07 $X=10250 $Y=17670 $D=616
M396 vss vss vss vss hvtnfet l=1.4e-07 w=7.5e-07 $X=10330 $Y=34593 $D=616
M397 vss 20 97 vss hvtnfet l=6e-08 w=4e-07 $X=10345 $Y=4836 $D=616
M398 vss b_ma<2> 1065 vss hvtnfet l=6e-08 w=4e-07 $X=10345 $Y=11331 $D=616
M399 vss 22 1066 vss hvtnfet l=6e-08 w=4e-07 $X=10345 $Y=12191 $D=616
M400 vss 23 1067 vss hvtnfet l=6e-08 w=4e-07 $X=10345 $Y=38542 $D=616
M401 vss t_ma<2> 1068 vss hvtnfet l=6e-08 w=4e-07 $X=10345 $Y=39402 $D=616
M402 vss 20 98 vss hvtnfet l=6e-08 w=4e-07 $X=10345 $Y=45897 $D=616
M403 475 vdd vss vss hvtnfet l=1.4e-07 w=2.1e-07 $X=10375 $Y=14550 $D=616
M404 476 vdd vss vss hvtnfet l=1.4e-07 w=2.1e-07 $X=10375 $Y=16760 $D=616
M405 vss vss vss vss hvtnfet l=6e-08 w=3e-07 $X=10457 $Y=31223 $D=616
M406 vss vss vss vss hvtnfet l=8e-08 w=3.75e-07 $X=10490 $Y=33798 $D=616
M407 477 vdd vss vss hvtnfet l=6e-08 w=3e-07 $X=10510 $Y=17670 $D=616
M408 101 11 vss vss hvtnfet l=6e-08 w=4e-07 $X=10605 $Y=4836 $D=616
M409 1069 b_mb<2> vss vss hvtnfet l=6e-08 w=4e-07 $X=10605 $Y=11331 $D=616
M410 1070 13 vss vss hvtnfet l=6e-08 w=4e-07 $X=10605 $Y=12191 $D=616
M411 1071 14 vss vss hvtnfet l=6e-08 w=4e-07 $X=10605 $Y=38542 $D=616
M412 1072 t_mb<2> vss vss hvtnfet l=6e-08 w=4e-07 $X=10605 $Y=39402 $D=616
M413 102 11 vss vss hvtnfet l=6e-08 w=4e-07 $X=10605 $Y=45897 $D=616
M414 299 101 b_blb<10> vss hvtnfet l=6e-08 w=6e-07 $X=10650 $Y=2941 $D=616
M415 299 101 b_blb<10> vss hvtnfet l=6e-08 w=6e-07 $X=10650 $Y=3201 $D=616
M416 308 97 b_bla_n<10> vss hvtnfet l=6e-08 w=6e-07 $X=10650 $Y=3881 $D=616
M417 308 97 b_bla_n<10> vss hvtnfet l=6e-08 w=6e-07 $X=10650 $Y=4141 $D=616
M418 t_bla_n<10> 98 308 vss hvtnfet l=6e-08 w=6e-07 $X=10650 $Y=46932 $D=616
M419 308 98 t_bla_n<10> vss hvtnfet l=6e-08 w=6e-07 $X=10650 $Y=47192 $D=616
M420 t_blb<10> 102 299 vss hvtnfet l=6e-08 w=6e-07 $X=10650 $Y=47872 $D=616
M421 299 102 t_blb<10> vss hvtnfet l=6e-08 w=6e-07 $X=10650 $Y=48132 $D=616
M422 vss vss vss vss hvtnfet l=1.4e-07 w=7.5e-07 $X=10670 $Y=34593 $D=616
M423 vss vdd 475 vss hvtnfet l=1.4e-07 w=2.1e-07 $X=10715 $Y=14550 $D=616
M424 vss vdd 476 vss hvtnfet l=1.4e-07 w=2.1e-07 $X=10715 $Y=16760 $D=616
M425 484 vdd vss vss hvtnfet l=6e-08 w=6e-07 $X=10717 $Y=26159 $D=616
M426 vss vdd 477 vss hvtnfet l=6e-08 w=3e-07 $X=10770 $Y=17670 $D=616
M427 vss vss vss vss hvtnfet l=7e-08 w=3.2e-07 $X=10780 $Y=33798 $D=616
M428 vss 99 101 vss hvtnfet l=6e-08 w=4e-07 $X=10865 $Y=4836 $D=616
M429 99 b_cb<2> 1069 vss hvtnfet l=6e-08 w=4e-07 $X=10865 $Y=11331 $D=616
M430 103 99 1070 vss hvtnfet l=6e-08 w=4e-07 $X=10865 $Y=12191 $D=616
M431 104 100 1071 vss hvtnfet l=6e-08 w=4e-07 $X=10865 $Y=38542 $D=616
M432 100 t_cb<2> 1072 vss hvtnfet l=6e-08 w=4e-07 $X=10865 $Y=39402 $D=616
M433 vss 100 102 vss hvtnfet l=6e-08 w=4e-07 $X=10865 $Y=45897 $D=616
M434 vss vdd 484 vss hvtnfet l=6e-08 w=6e-07 $X=10977 $Y=26159 $D=616
M435 299 112 b_blb<9> vss hvtnfet l=6e-08 w=6e-07 $X=11670 $Y=2941 $D=616
M436 299 112 b_blb<9> vss hvtnfet l=6e-08 w=6e-07 $X=11670 $Y=3201 $D=616
M437 308 120 b_bla_n<9> vss hvtnfet l=6e-08 w=6e-07 $X=11670 $Y=3881 $D=616
M438 308 120 b_bla_n<9> vss hvtnfet l=6e-08 w=6e-07 $X=11670 $Y=4141 $D=616
M439 t_bla_n<9> 121 308 vss hvtnfet l=6e-08 w=6e-07 $X=11670 $Y=46932 $D=616
M440 308 121 t_bla_n<9> vss hvtnfet l=6e-08 w=6e-07 $X=11670 $Y=47192 $D=616
M441 t_blb<9> 113 299 vss hvtnfet l=6e-08 w=6e-07 $X=11670 $Y=47872 $D=616
M442 299 113 t_blb<9> vss hvtnfet l=6e-08 w=6e-07 $X=11670 $Y=48132 $D=616
M443 308 119 vss vss hvtnfet l=6e-08 w=6e-07 $X=11883 $Y=26159 $D=616
M444 112 107 vss vss hvtnfet l=6e-08 w=4e-07 $X=11995 $Y=4836 $D=616
M445 1073 b_cb<1> 107 vss hvtnfet l=6e-08 w=4e-07 $X=11995 $Y=11331 $D=616
M446 1074 107 105 vss hvtnfet l=6e-08 w=4e-07 $X=11995 $Y=12191 $D=616
M447 1075 108 106 vss hvtnfet l=6e-08 w=4e-07 $X=11995 $Y=38542 $D=616
M448 1076 t_cb<1> 108 vss hvtnfet l=6e-08 w=4e-07 $X=11995 $Y=39402 $D=616
M449 113 108 vss vss hvtnfet l=6e-08 w=4e-07 $X=11995 $Y=45897 $D=616
M450 vss vdd 498 vss hvtnfet l=6e-08 w=3e-07 $X=12033 $Y=31223 $D=616
M451 vss bwena 122 vss hvtnfet l=1.4e-07 w=2.1e-07 $X=12065 $Y=14555 $D=616
M452 vss 114 134 vss hvtnfet l=1.4e-07 w=2.1e-07 $X=12065 $Y=16755 $D=616
M453 vss 115 ddqa_n vss hvtnfet l=7e-08 w=3.2e-07 $X=12070 $Y=33798 $D=616
M454 516 vdd vss vss hvtnfet l=6e-08 w=3e-07 $X=12090 $Y=17670 $D=616
M455 115 117 538 vss hvtnfet l=1.4e-07 w=7.5e-07 $X=12110 $Y=34593 $D=616
M456 vss 119 308 vss hvtnfet l=6e-08 w=6e-07 $X=12143 $Y=26159 $D=616
M457 vss 11 112 vss hvtnfet l=6e-08 w=4e-07 $X=12255 $Y=4836 $D=616
M458 vss b_mb<2> 1073 vss hvtnfet l=6e-08 w=4e-07 $X=12255 $Y=11331 $D=616
M459 vss 13 1074 vss hvtnfet l=6e-08 w=4e-07 $X=12255 $Y=12191 $D=616
M460 vss 14 1075 vss hvtnfet l=6e-08 w=4e-07 $X=12255 $Y=38542 $D=616
M461 vss t_mb<2> 1076 vss hvtnfet l=6e-08 w=4e-07 $X=12255 $Y=39402 $D=616
M462 vss 11 113 vss hvtnfet l=6e-08 w=4e-07 $X=12255 $Y=45897 $D=616
M463 vss vdd 516 vss hvtnfet l=6e-08 w=3e-07 $X=12350 $Y=17670 $D=616
M464 538 118 vss vss hvtnfet l=8e-08 w=3.75e-07 $X=12350 $Y=33798 $D=616
M465 130 122 vss vss hvtnfet l=1.4e-07 w=2.1e-07 $X=12405 $Y=14555 $D=616
M466 114 133 vss vss hvtnfet l=1.4e-07 w=2.1e-07 $X=12405 $Y=16755 $D=616
M467 538 117 115 vss hvtnfet l=1.4e-07 w=7.5e-07 $X=12450 $Y=34593 $D=616
M468 120 20 vss vss hvtnfet l=6e-08 w=4e-07 $X=12515 $Y=4836 $D=616
M469 1077 b_ma<2> vss vss hvtnfet l=6e-08 w=4e-07 $X=12515 $Y=11331 $D=616
M470 1078 22 vss vss hvtnfet l=6e-08 w=4e-07 $X=12515 $Y=12191 $D=616
M471 1079 23 vss vss hvtnfet l=6e-08 w=4e-07 $X=12515 $Y=38542 $D=616
M472 1080 t_ma<2> vss vss hvtnfet l=6e-08 w=4e-07 $X=12515 $Y=39402 $D=616
M473 121 20 vss vss hvtnfet l=6e-08 w=4e-07 $X=12515 $Y=45897 $D=616
M474 1081 118 vss vss hvtnfet l=6e-08 w=3e-07 $X=12543 $Y=31223 $D=616
M475 317 112 b_blb_n<9> vss hvtnfet l=6e-08 w=6e-07 $X=12560 $Y=2941 $D=616
M476 317 112 b_blb_n<9> vss hvtnfet l=6e-08 w=6e-07 $X=12560 $Y=3201 $D=616
M477 b_bla<9> 120 328 vss hvtnfet l=6e-08 w=6e-07 $X=12560 $Y=3881 $D=616
M478 b_bla<9> 120 328 vss hvtnfet l=6e-08 w=6e-07 $X=12560 $Y=4141 $D=616
M479 328 121 t_bla<9> vss hvtnfet l=6e-08 w=6e-07 $X=12560 $Y=46932 $D=616
M480 t_bla<9> 121 328 vss hvtnfet l=6e-08 w=6e-07 $X=12560 $Y=47192 $D=616
M481 t_blb_n<9> 113 317 vss hvtnfet l=6e-08 w=6e-07 $X=12560 $Y=47872 $D=616
M482 317 113 t_blb_n<9> vss hvtnfet l=6e-08 w=6e-07 $X=12560 $Y=48132 $D=616
M483 516 vdd vss vss hvtnfet l=6e-08 w=3e-07 $X=12610 $Y=17670 $D=616
M484 vss 118 538 vss hvtnfet l=8e-08 w=3.75e-07 $X=12630 $Y=33798 $D=616
M485 vss 126 521 vss hvtnfet l=6e-08 w=8e-07 $X=12653 $Y=26159 $D=616
M486 138 115 1081 vss hvtnfet l=6e-08 w=3e-07 $X=12733 $Y=31223 $D=616
M487 vss 123 120 vss hvtnfet l=6e-08 w=4e-07 $X=12775 $Y=4836 $D=616
M488 123 b_ca<1> 1077 vss hvtnfet l=6e-08 w=4e-07 $X=12775 $Y=11331 $D=616
M489 127 123 1078 vss hvtnfet l=6e-08 w=4e-07 $X=12775 $Y=12191 $D=616
M490 128 124 1079 vss hvtnfet l=6e-08 w=4e-07 $X=12775 $Y=38542 $D=616
M491 124 t_ca<1> 1080 vss hvtnfet l=6e-08 w=4e-07 $X=12775 $Y=39402 $D=616
M492 vss 124 121 vss hvtnfet l=6e-08 w=4e-07 $X=12775 $Y=45897 $D=616
M493 117 115 538 vss hvtnfet l=1.4e-07 w=7.5e-07 $X=12790 $Y=34593 $D=616
M494 vss vdd 516 vss hvtnfet l=6e-08 w=3e-07 $X=12870 $Y=17670 $D=616
M495 538 118 vss vss hvtnfet l=8e-08 w=3.75e-07 $X=12910 $Y=33798 $D=616
M496 521 126 vss vss hvtnfet l=6e-08 w=8e-07 $X=12913 $Y=26159 $D=616
M497 1082 125 138 vss hvtnfet l=6e-08 w=3e-07 $X=12993 $Y=31223 $D=616
M498 vss 130 141 vss hvtnfet l=1.4e-07 w=2.1e-07 $X=12995 $Y=14555 $D=616
M499 vss 136 133 vss hvtnfet l=1.4e-07 w=2.1e-07 $X=12995 $Y=16755 $D=616
M500 qa 125 vss vss hvtnfet l=6e-08 w=4.5e-07 $X=13075 $Y=19812 $D=616
M501 vss 125 qa vss hvtnfet l=6e-08 w=4.5e-07 $X=13075 $Y=20072 $D=616
M502 1083 134 vss vss hvtnfet l=6e-08 w=3.2e-07 $X=13075 $Y=21012 $D=616
M503 1083 129 131 vss hvtnfet l=6e-08 w=3.2e-07 $X=13075 $Y=21202 $D=616
M504 1084 111 131 vss hvtnfet l=6e-08 w=1.4e-07 $X=13075 $Y=21477 $D=616
M505 vss 109 1084 vss hvtnfet l=6e-08 w=1.4e-07 $X=13075 $Y=21667 $D=616
M506 111 131 vss vss hvtnfet l=6e-08 w=2.1e-07 $X=13075 $Y=21942 $D=616
M507 vss 131 119 vss hvtnfet l=6e-08 w=3.2e-07 $X=13075 $Y=22762 $D=616
M508 1085 135 vss vss hvtnfet l=6e-08 w=3.2e-07 $X=13075 $Y=23729 $D=616
M509 1085 129 132 vss hvtnfet l=6e-08 w=3.2e-07 $X=13075 $Y=23919 $D=616
M510 1086 110 132 vss hvtnfet l=6e-08 w=1.4e-07 $X=13075 $Y=24194 $D=616
M511 vss 109 1086 vss hvtnfet l=6e-08 w=1.4e-07 $X=13075 $Y=24384 $D=616
M512 110 132 vss vss hvtnfet l=6e-08 w=2.1e-07 $X=13075 $Y=24659 $D=616
M513 516 vdd vss vss hvtnfet l=6e-08 w=3e-07 $X=13130 $Y=17670 $D=616
M514 538 115 117 vss hvtnfet l=1.4e-07 w=7.5e-07 $X=13130 $Y=34593 $D=616
M515 20 lwea 521 vss hvtnfet l=6e-08 w=8e-07 $X=13173 $Y=26159 $D=616
M516 vss saea_n 1082 vss hvtnfet l=6e-08 w=3e-07 $X=13183 $Y=31223 $D=616
M517 vss 118 538 vss hvtnfet l=8e-08 w=3.75e-07 $X=13190 $Y=33798 $D=616
M518 135 141 vss vss hvtnfet l=1.4e-07 w=2.1e-07 $X=13335 $Y=14555 $D=616
M519 136 da vss vss hvtnfet l=1.4e-07 w=2.1e-07 $X=13335 $Y=16755 $D=616
M520 vss vdd 516 vss hvtnfet l=6e-08 w=3e-07 $X=13390 $Y=17670 $D=616
M521 521 lwea 20 vss hvtnfet l=6e-08 w=8e-07 $X=13433 $Y=26159 $D=616
M522 538 118 vss vss hvtnfet l=8e-08 w=3.75e-07 $X=13470 $Y=33798 $D=616
M523 115 117 538 vss hvtnfet l=1.4e-07 w=7.5e-07 $X=13470 $Y=34593 $D=616
M524 317 155 b_blb_n<8> vss hvtnfet l=6e-08 w=6e-07 $X=13580 $Y=2941 $D=616
M525 317 155 b_blb_n<8> vss hvtnfet l=6e-08 w=6e-07 $X=13580 $Y=3201 $D=616
M526 b_bla<8> 148 328 vss hvtnfet l=6e-08 w=6e-07 $X=13580 $Y=3881 $D=616
M527 b_bla<8> 148 328 vss hvtnfet l=6e-08 w=6e-07 $X=13580 $Y=4141 $D=616
M528 328 149 t_bla<8> vss hvtnfet l=6e-08 w=6e-07 $X=13580 $Y=46932 $D=616
M529 t_bla<8> 149 328 vss hvtnfet l=6e-08 w=6e-07 $X=13580 $Y=47192 $D=616
M530 t_blb_n<8> 156 317 vss hvtnfet l=6e-08 w=6e-07 $X=13580 $Y=47872 $D=616
M531 317 156 t_blb_n<8> vss hvtnfet l=6e-08 w=6e-07 $X=13580 $Y=48132 $D=616
M532 vss 118 538 vss hvtnfet l=8e-08 w=3.75e-07 $X=13750 $Y=33798 $D=616
M533 538 117 115 vss hvtnfet l=1.4e-07 w=7.5e-07 $X=13810 $Y=34593 $D=616
M534 22 b_tm_prea_n vss vss hvtnfet l=6e-08 w=2.5e-07 $X=13900 $Y=17720 $D=616
M535 148 143 vss vss hvtnfet l=6e-08 w=4e-07 $X=13905 $Y=4836 $D=616
M536 1087 b_ca<0> 143 vss hvtnfet l=6e-08 w=4e-07 $X=13905 $Y=11331 $D=616
M537 1088 143 145 vss hvtnfet l=6e-08 w=4e-07 $X=13905 $Y=12191 $D=616
M538 1089 144 146 vss hvtnfet l=6e-08 w=4e-07 $X=13905 $Y=38542 $D=616
M539 1090 t_ca<0> 144 vss hvtnfet l=6e-08 w=4e-07 $X=13905 $Y=39402 $D=616
M540 149 144 vss vss hvtnfet l=6e-08 w=4e-07 $X=13905 $Y=45897 $D=616
M541 328 131 vss vss hvtnfet l=6e-08 w=6e-07 $X=13953 $Y=26159 $D=616
M542 538 118 vss vss hvtnfet l=8e-08 w=3.75e-07 $X=14030 $Y=33798 $D=616
M543 vss 138 125 vss hvtnfet l=6e-08 w=3e-07 $X=14093 $Y=31223 $D=616
M544 129 clk_dqa vss vss hvtnfet l=6e-08 w=2e-07 $X=14105 $Y=21427 $D=616
M545 109 clk_dqa_n vss vss hvtnfet l=6e-08 w=2e-07 $X=14105 $Y=23694 $D=616
M546 152 132 vss vss hvtnfet l=6e-08 w=2e-07 $X=14105 $Y=24394 $D=616
M547 126 152 vss vss hvtnfet l=6e-08 w=2e-07 $X=14105 $Y=24904 $D=616
M548 117 115 538 vss hvtnfet l=1.4e-07 w=7.5e-07 $X=14150 $Y=34593 $D=616
M549 vss b_tm_prea_n 22 vss hvtnfet l=6e-08 w=2.5e-07 $X=14160 $Y=17720 $D=616
M550 vss 20 148 vss hvtnfet l=6e-08 w=4e-07 $X=14165 $Y=4836 $D=616
M551 vss b_ma<2> 1087 vss hvtnfet l=6e-08 w=4e-07 $X=14165 $Y=11331 $D=616
M552 vss 22 1088 vss hvtnfet l=6e-08 w=4e-07 $X=14165 $Y=12191 $D=616
M553 vss 23 1089 vss hvtnfet l=6e-08 w=4e-07 $X=14165 $Y=38542 $D=616
M554 vss t_ma<2> 1090 vss hvtnfet l=6e-08 w=4e-07 $X=14165 $Y=39402 $D=616
M555 vss 20 149 vss hvtnfet l=6e-08 w=4e-07 $X=14165 $Y=45897 $D=616
M556 vss 131 328 vss hvtnfet l=6e-08 w=6e-07 $X=14213 $Y=26159 $D=616
M557 vss 118 538 vss hvtnfet l=8e-08 w=3.75e-07 $X=14310 $Y=33798 $D=616
M558 118 saea_n vss vss hvtnfet l=6e-08 w=3e-07 $X=14353 $Y=31223 $D=616
M559 23 t_tm_prea_n vss vss hvtnfet l=6e-08 w=2.5e-07 $X=14420 $Y=17720 $D=616
M560 155 11 vss vss hvtnfet l=6e-08 w=4e-07 $X=14425 $Y=4836 $D=616
M561 1091 b_mb<2> vss vss hvtnfet l=6e-08 w=4e-07 $X=14425 $Y=11331 $D=616
M562 1092 13 vss vss hvtnfet l=6e-08 w=4e-07 $X=14425 $Y=12191 $D=616
M563 1093 14 vss vss hvtnfet l=6e-08 w=4e-07 $X=14425 $Y=38542 $D=616
M564 1094 t_mb<2> vss vss hvtnfet l=6e-08 w=4e-07 $X=14425 $Y=39402 $D=616
M565 156 11 vss vss hvtnfet l=6e-08 w=4e-07 $X=14425 $Y=45897 $D=616
M566 299 155 b_blb<8> vss hvtnfet l=6e-08 w=6e-07 $X=14470 $Y=2941 $D=616
M567 299 155 b_blb<8> vss hvtnfet l=6e-08 w=6e-07 $X=14470 $Y=3201 $D=616
M568 308 148 b_bla_n<8> vss hvtnfet l=6e-08 w=6e-07 $X=14470 $Y=3881 $D=616
M569 308 148 b_bla_n<8> vss hvtnfet l=6e-08 w=6e-07 $X=14470 $Y=4141 $D=616
M570 t_bla_n<8> 149 308 vss hvtnfet l=6e-08 w=6e-07 $X=14470 $Y=46932 $D=616
M571 308 149 t_bla_n<8> vss hvtnfet l=6e-08 w=6e-07 $X=14470 $Y=47192 $D=616
M572 t_blb<8> 156 299 vss hvtnfet l=6e-08 w=6e-07 $X=14470 $Y=47872 $D=616
M573 299 156 t_blb<8> vss hvtnfet l=6e-08 w=6e-07 $X=14470 $Y=48132 $D=616
M574 538 115 117 vss hvtnfet l=1.4e-07 w=7.5e-07 $X=14490 $Y=34593 $D=616
M575 ddqa 117 vss vss hvtnfet l=7e-08 w=3.2e-07 $X=14600 $Y=33798 $D=616
M576 vss t_tm_prea_n 23 vss hvtnfet l=6e-08 w=2.5e-07 $X=14680 $Y=17720 $D=616
M577 vss 153 155 vss hvtnfet l=6e-08 w=4e-07 $X=14685 $Y=4836 $D=616
M578 153 b_cb<0> 1091 vss hvtnfet l=6e-08 w=4e-07 $X=14685 $Y=11331 $D=616
M579 157 153 1092 vss hvtnfet l=6e-08 w=4e-07 $X=14685 $Y=12191 $D=616
M580 158 154 1093 vss hvtnfet l=6e-08 w=4e-07 $X=14685 $Y=38542 $D=616
M581 154 t_cb<0> 1094 vss hvtnfet l=6e-08 w=4e-07 $X=14685 $Y=39402 $D=616
M582 vss 154 156 vss hvtnfet l=6e-08 w=4e-07 $X=14685 $Y=45897 $D=616
M583 544 117 vss vss hvtnfet l=6e-08 w=3e-07 $X=14863 $Y=31223 $D=616
M584 299 166 b_blb<7> vss hvtnfet l=6e-08 w=6e-07 $X=15490 $Y=2941 $D=616
M585 299 166 b_blb<7> vss hvtnfet l=6e-08 w=6e-07 $X=15490 $Y=3201 $D=616
M586 308 176 b_bla_n<7> vss hvtnfet l=6e-08 w=6e-07 $X=15490 $Y=3881 $D=616
M587 308 176 b_bla_n<7> vss hvtnfet l=6e-08 w=6e-07 $X=15490 $Y=4141 $D=616
M588 t_bla_n<7> 177 308 vss hvtnfet l=6e-08 w=6e-07 $X=15490 $Y=46932 $D=616
M589 308 177 t_bla_n<7> vss hvtnfet l=6e-08 w=6e-07 $X=15490 $Y=47192 $D=616
M590 t_blb<7> 167 299 vss hvtnfet l=6e-08 w=6e-07 $X=15490 $Y=47872 $D=616
M591 299 167 t_blb<7> vss hvtnfet l=6e-08 w=6e-07 $X=15490 $Y=48132 $D=616
M592 vss 160 551 vss hvtnfet l=6e-08 w=3e-07 $X=15637 $Y=31223 $D=616
M593 166 163 vss vss hvtnfet l=6e-08 w=4e-07 $X=15815 $Y=4836 $D=616
M594 1095 b_cb<3> 163 vss hvtnfet l=6e-08 w=4e-07 $X=15815 $Y=11331 $D=616
M595 1096 163 161 vss hvtnfet l=6e-08 w=4e-07 $X=15815 $Y=12191 $D=616
M596 1097 164 162 vss hvtnfet l=6e-08 w=4e-07 $X=15815 $Y=38542 $D=616
M597 1098 t_cb<3> 164 vss hvtnfet l=6e-08 w=4e-07 $X=15815 $Y=39402 $D=616
M598 167 164 vss vss hvtnfet l=6e-08 w=4e-07 $X=15815 $Y=45897 $D=616
M599 14 t_tm_preb_n vss vss hvtnfet l=6e-08 w=2.5e-07 $X=15820 $Y=17720 $D=616
M600 vss 160 ddqb vss hvtnfet l=7e-08 w=3.2e-07 $X=15890 $Y=33798 $D=616
M601 160 168 594 vss hvtnfet l=1.4e-07 w=7.5e-07 $X=15930 $Y=34593 $D=616
M602 vss 11 166 vss hvtnfet l=6e-08 w=4e-07 $X=16075 $Y=4836 $D=616
M603 vss b_mb<1> 1095 vss hvtnfet l=6e-08 w=4e-07 $X=16075 $Y=11331 $D=616
M604 vss 13 1096 vss hvtnfet l=6e-08 w=4e-07 $X=16075 $Y=12191 $D=616
M605 vss 14 1097 vss hvtnfet l=6e-08 w=4e-07 $X=16075 $Y=38542 $D=616
M606 vss t_mb<1> 1098 vss hvtnfet l=6e-08 w=4e-07 $X=16075 $Y=39402 $D=616
M607 vss 11 167 vss hvtnfet l=6e-08 w=4e-07 $X=16075 $Y=45897 $D=616
M608 vss t_tm_preb_n 14 vss hvtnfet l=6e-08 w=2.5e-07 $X=16080 $Y=17720 $D=616
M609 vss saeb_n 169 vss hvtnfet l=6e-08 w=3e-07 $X=16147 $Y=31223 $D=616
M610 594 169 vss vss hvtnfet l=8e-08 w=3.75e-07 $X=16170 $Y=33798 $D=616
M611 192 clk_dqb vss vss hvtnfet l=6e-08 w=2e-07 $X=16255 $Y=21427 $D=616
M612 190 clk_dqb_n vss vss hvtnfet l=6e-08 w=2e-07 $X=16255 $Y=23694 $D=616
M613 174 173 vss vss hvtnfet l=6e-08 w=2e-07 $X=16255 $Y=24394 $D=616
M614 200 174 vss vss hvtnfet l=6e-08 w=2e-07 $X=16255 $Y=24904 $D=616
M615 594 168 160 vss hvtnfet l=1.4e-07 w=7.5e-07 $X=16270 $Y=34593 $D=616
M616 299 178 vss vss hvtnfet l=6e-08 w=6e-07 $X=16287 $Y=26159 $D=616
M617 176 20 vss vss hvtnfet l=6e-08 w=4e-07 $X=16335 $Y=4836 $D=616
M618 1099 b_ma<1> vss vss hvtnfet l=6e-08 w=4e-07 $X=16335 $Y=11331 $D=616
M619 1100 22 vss vss hvtnfet l=6e-08 w=4e-07 $X=16335 $Y=12191 $D=616
M620 1101 23 vss vss hvtnfet l=6e-08 w=4e-07 $X=16335 $Y=38542 $D=616
M621 1102 t_ma<1> vss vss hvtnfet l=6e-08 w=4e-07 $X=16335 $Y=39402 $D=616
M622 177 20 vss vss hvtnfet l=6e-08 w=4e-07 $X=16335 $Y=45897 $D=616
M623 13 b_tm_preb_n vss vss hvtnfet l=6e-08 w=2.5e-07 $X=16340 $Y=17720 $D=616
M624 317 166 b_blb_n<7> vss hvtnfet l=6e-08 w=6e-07 $X=16380 $Y=2941 $D=616
M625 317 166 b_blb_n<7> vss hvtnfet l=6e-08 w=6e-07 $X=16380 $Y=3201 $D=616
M626 b_bla<7> 176 328 vss hvtnfet l=6e-08 w=6e-07 $X=16380 $Y=3881 $D=616
M627 b_bla<7> 176 328 vss hvtnfet l=6e-08 w=6e-07 $X=16380 $Y=4141 $D=616
M628 328 177 t_bla<7> vss hvtnfet l=6e-08 w=6e-07 $X=16380 $Y=46932 $D=616
M629 t_bla<7> 177 328 vss hvtnfet l=6e-08 w=6e-07 $X=16380 $Y=47192 $D=616
M630 t_blb_n<7> 167 317 vss hvtnfet l=6e-08 w=6e-07 $X=16380 $Y=47872 $D=616
M631 317 167 t_blb_n<7> vss hvtnfet l=6e-08 w=6e-07 $X=16380 $Y=48132 $D=616
M632 189 194 vss vss hvtnfet l=6e-08 w=3e-07 $X=16407 $Y=31223 $D=616
M633 vss 169 594 vss hvtnfet l=8e-08 w=3.75e-07 $X=16450 $Y=33798 $D=616
M634 vss 178 299 vss hvtnfet l=6e-08 w=6e-07 $X=16547 $Y=26159 $D=616
M635 vss 179 176 vss hvtnfet l=6e-08 w=4e-07 $X=16595 $Y=4836 $D=616
M636 179 b_ca<3> 1099 vss hvtnfet l=6e-08 w=4e-07 $X=16595 $Y=11331 $D=616
M637 184 179 1100 vss hvtnfet l=6e-08 w=4e-07 $X=16595 $Y=12191 $D=616
M638 185 180 1101 vss hvtnfet l=6e-08 w=4e-07 $X=16595 $Y=38542 $D=616
M639 180 t_ca<3> 1102 vss hvtnfet l=6e-08 w=4e-07 $X=16595 $Y=39402 $D=616
M640 vss 180 177 vss hvtnfet l=6e-08 w=4e-07 $X=16595 $Y=45897 $D=616
M641 vss b_tm_preb_n 13 vss hvtnfet l=6e-08 w=2.5e-07 $X=16600 $Y=17720 $D=616
M642 168 160 594 vss hvtnfet l=1.4e-07 w=7.5e-07 $X=16610 $Y=34593 $D=616
M643 594 169 vss vss hvtnfet l=8e-08 w=3.75e-07 $X=16730 $Y=33798 $D=616
M644 594 160 168 vss hvtnfet l=1.4e-07 w=7.5e-07 $X=16950 $Y=34593 $D=616
M645 vss 169 594 vss hvtnfet l=8e-08 w=3.75e-07 $X=17010 $Y=33798 $D=616
M646 qb 189 vss vss hvtnfet l=6e-08 w=4.5e-07 $X=17035 $Y=19812 $D=616
M647 vss 189 qb vss hvtnfet l=6e-08 w=4.5e-07 $X=17035 $Y=20072 $D=616
M648 11 lweb 582 vss hvtnfet l=6e-08 w=8e-07 $X=17067 $Y=26159 $D=616
M649 vss 191 202 vss hvtnfet l=1.4e-07 w=2.1e-07 $X=17085 $Y=14555 $D=616
M650 vss db 195 vss hvtnfet l=1.4e-07 w=2.1e-07 $X=17085 $Y=16755 $D=616
M651 587 vdd vss vss hvtnfet l=6e-08 w=3e-07 $X=17110 $Y=17670 $D=616
M652 1103 201 vss vss hvtnfet l=6e-08 w=3.2e-07 $X=17165 $Y=21012 $D=616
M653 1103 192 178 vss hvtnfet l=6e-08 w=3.2e-07 $X=17165 $Y=21202 $D=616
M654 vss 178 208 vss hvtnfet l=6e-08 w=3.2e-07 $X=17165 $Y=22762 $D=616
M655 1104 202 vss vss hvtnfet l=6e-08 w=3.2e-07 $X=17165 $Y=23729 $D=616
M656 1104 192 173 vss hvtnfet l=6e-08 w=3.2e-07 $X=17165 $Y=23919 $D=616
M657 217 178 vss vss hvtnfet l=6e-08 w=2.1e-07 $X=17275 $Y=21942 $D=616
M658 218 173 vss vss hvtnfet l=6e-08 w=2.1e-07 $X=17275 $Y=24659 $D=616
M659 594 169 vss vss hvtnfet l=8e-08 w=3.75e-07 $X=17290 $Y=33798 $D=616
M660 160 168 594 vss hvtnfet l=1.4e-07 w=7.5e-07 $X=17290 $Y=34593 $D=616
M661 1107 saeb_n vss vss hvtnfet l=6e-08 w=3e-07 $X=17317 $Y=31223 $D=616
M662 582 lweb 11 vss hvtnfet l=6e-08 w=8e-07 $X=17327 $Y=26159 $D=616
M663 1105 217 178 vss hvtnfet l=6e-08 w=1.4e-07 $X=17345 $Y=21477 $D=616
M664 vss 190 1105 vss hvtnfet l=6e-08 w=1.4e-07 $X=17345 $Y=21667 $D=616
M665 1106 218 173 vss hvtnfet l=6e-08 w=1.4e-07 $X=17345 $Y=24194 $D=616
M666 vss 190 1106 vss hvtnfet l=6e-08 w=1.4e-07 $X=17345 $Y=24384 $D=616
M667 vss vdd 587 vss hvtnfet l=6e-08 w=3e-07 $X=17370 $Y=17670 $D=616
M668 317 211 b_blb_n<6> vss hvtnfet l=6e-08 w=6e-07 $X=17400 $Y=2941 $D=616
M669 317 211 b_blb_n<6> vss hvtnfet l=6e-08 w=6e-07 $X=17400 $Y=3201 $D=616
M670 b_bla<6> 205 328 vss hvtnfet l=6e-08 w=6e-07 $X=17400 $Y=3881 $D=616
M671 b_bla<6> 205 328 vss hvtnfet l=6e-08 w=6e-07 $X=17400 $Y=4141 $D=616
M672 328 206 t_bla<6> vss hvtnfet l=6e-08 w=6e-07 $X=17400 $Y=46932 $D=616
M673 t_bla<6> 206 328 vss hvtnfet l=6e-08 w=6e-07 $X=17400 $Y=47192 $D=616
M674 t_blb_n<6> 212 317 vss hvtnfet l=6e-08 w=6e-07 $X=17400 $Y=47872 $D=616
M675 317 212 t_blb_n<6> vss hvtnfet l=6e-08 w=6e-07 $X=17400 $Y=48132 $D=616
M676 191 204 vss vss hvtnfet l=1.4e-07 w=2.1e-07 $X=17425 $Y=14555 $D=616
M677 203 195 vss vss hvtnfet l=1.4e-07 w=2.1e-07 $X=17425 $Y=16755 $D=616
M678 194 189 1107 vss hvtnfet l=6e-08 w=3e-07 $X=17507 $Y=31223 $D=616
M679 vss 169 594 vss hvtnfet l=8e-08 w=3.75e-07 $X=17570 $Y=33798 $D=616
M680 vss 200 582 vss hvtnfet l=6e-08 w=8e-07 $X=17587 $Y=26159 $D=616
M681 587 vdd vss vss hvtnfet l=6e-08 w=3e-07 $X=17630 $Y=17670 $D=616
M682 594 168 160 vss hvtnfet l=1.4e-07 w=7.5e-07 $X=17630 $Y=34593 $D=616
M683 205 196 vss vss hvtnfet l=6e-08 w=4e-07 $X=17725 $Y=4836 $D=616
M684 1108 b_ca<2> 196 vss hvtnfet l=6e-08 w=4e-07 $X=17725 $Y=11331 $D=616
M685 1109 196 198 vss hvtnfet l=6e-08 w=4e-07 $X=17725 $Y=12191 $D=616
M686 1110 197 199 vss hvtnfet l=6e-08 w=4e-07 $X=17725 $Y=38542 $D=616
M687 1111 t_ca<2> 197 vss hvtnfet l=6e-08 w=4e-07 $X=17725 $Y=39402 $D=616
M688 206 197 vss vss hvtnfet l=6e-08 w=4e-07 $X=17725 $Y=45897 $D=616
M689 1112 168 194 vss hvtnfet l=6e-08 w=3e-07 $X=17767 $Y=31223 $D=616
M690 582 200 vss vss hvtnfet l=6e-08 w=8e-07 $X=17847 $Y=26159 $D=616
M691 594 169 vss vss hvtnfet l=8e-08 w=3.75e-07 $X=17850 $Y=33798 $D=616
M692 vss vdd 587 vss hvtnfet l=6e-08 w=3e-07 $X=17890 $Y=17670 $D=616
M693 vss 169 1112 vss hvtnfet l=6e-08 w=3e-07 $X=17957 $Y=31223 $D=616
M694 168 160 594 vss hvtnfet l=1.4e-07 w=7.5e-07 $X=17970 $Y=34593 $D=616
M695 vss 20 205 vss hvtnfet l=6e-08 w=4e-07 $X=17985 $Y=4836 $D=616
M696 vss b_ma<1> 1108 vss hvtnfet l=6e-08 w=4e-07 $X=17985 $Y=11331 $D=616
M697 vss 22 1109 vss hvtnfet l=6e-08 w=4e-07 $X=17985 $Y=12191 $D=616
M698 vss 23 1110 vss hvtnfet l=6e-08 w=4e-07 $X=17985 $Y=38542 $D=616
M699 vss t_ma<1> 1111 vss hvtnfet l=6e-08 w=4e-07 $X=17985 $Y=39402 $D=616
M700 vss 20 206 vss hvtnfet l=6e-08 w=4e-07 $X=17985 $Y=45897 $D=616
M701 vss 207 204 vss hvtnfet l=1.4e-07 w=2.1e-07 $X=18015 $Y=14555 $D=616
M702 vss 203 216 vss hvtnfet l=1.4e-07 w=2.1e-07 $X=18015 $Y=16755 $D=616
M703 vss 169 594 vss hvtnfet l=8e-08 w=3.75e-07 $X=18130 $Y=33798 $D=616
M704 587 vdd vss vss hvtnfet l=6e-08 w=3e-07 $X=18150 $Y=17670 $D=616
M705 211 11 vss vss hvtnfet l=6e-08 w=4e-07 $X=18245 $Y=4836 $D=616
M706 1113 b_mb<1> vss vss hvtnfet l=6e-08 w=4e-07 $X=18245 $Y=11331 $D=616
M707 1114 13 vss vss hvtnfet l=6e-08 w=4e-07 $X=18245 $Y=12191 $D=616
M708 1115 14 vss vss hvtnfet l=6e-08 w=4e-07 $X=18245 $Y=38542 $D=616
M709 1116 t_mb<1> vss vss hvtnfet l=6e-08 w=4e-07 $X=18245 $Y=39402 $D=616
M710 212 11 vss vss hvtnfet l=6e-08 w=4e-07 $X=18245 $Y=45897 $D=616
M711 299 211 b_blb<6> vss hvtnfet l=6e-08 w=6e-07 $X=18290 $Y=2941 $D=616
M712 299 211 b_blb<6> vss hvtnfet l=6e-08 w=6e-07 $X=18290 $Y=3201 $D=616
M713 308 205 b_bla_n<6> vss hvtnfet l=6e-08 w=6e-07 $X=18290 $Y=3881 $D=616
M714 308 205 b_bla_n<6> vss hvtnfet l=6e-08 w=6e-07 $X=18290 $Y=4141 $D=616
M715 t_bla_n<6> 206 308 vss hvtnfet l=6e-08 w=6e-07 $X=18290 $Y=46932 $D=616
M716 308 206 t_bla_n<6> vss hvtnfet l=6e-08 w=6e-07 $X=18290 $Y=47192 $D=616
M717 t_blb<6> 212 299 vss hvtnfet l=6e-08 w=6e-07 $X=18290 $Y=47872 $D=616
M718 299 212 t_blb<6> vss hvtnfet l=6e-08 w=6e-07 $X=18290 $Y=48132 $D=616
M719 594 160 168 vss hvtnfet l=1.4e-07 w=7.5e-07 $X=18310 $Y=34593 $D=616
M720 207 bwenb vss vss hvtnfet l=1.4e-07 w=2.1e-07 $X=18355 $Y=14555 $D=616
M721 201 216 vss vss hvtnfet l=1.4e-07 w=2.1e-07 $X=18355 $Y=16755 $D=616
M722 317 208 vss vss hvtnfet l=6e-08 w=6e-07 $X=18357 $Y=26159 $D=616
M723 vss vdd 587 vss hvtnfet l=6e-08 w=3e-07 $X=18410 $Y=17670 $D=616
M724 ddqb_n 168 vss vss hvtnfet l=7e-08 w=3.2e-07 $X=18420 $Y=33798 $D=616
M725 598 vdd vss vss hvtnfet l=6e-08 w=3e-07 $X=18467 $Y=31223 $D=616
M726 vss 209 211 vss hvtnfet l=6e-08 w=4e-07 $X=18505 $Y=4836 $D=616
M727 209 b_cb<2> 1113 vss hvtnfet l=6e-08 w=4e-07 $X=18505 $Y=11331 $D=616
M728 214 209 1114 vss hvtnfet l=6e-08 w=4e-07 $X=18505 $Y=12191 $D=616
M729 215 210 1115 vss hvtnfet l=6e-08 w=4e-07 $X=18505 $Y=38542 $D=616
M730 210 t_cb<2> 1116 vss hvtnfet l=6e-08 w=4e-07 $X=18505 $Y=39402 $D=616
M731 vss 210 212 vss hvtnfet l=6e-08 w=4e-07 $X=18505 $Y=45897 $D=616
M732 vss 208 317 vss hvtnfet l=6e-08 w=6e-07 $X=18617 $Y=26159 $D=616
M733 299 223 b_blb<5> vss hvtnfet l=6e-08 w=6e-07 $X=19310 $Y=2941 $D=616
M734 299 223 b_blb<5> vss hvtnfet l=6e-08 w=6e-07 $X=19310 $Y=3201 $D=616
M735 308 225 b_bla_n<5> vss hvtnfet l=6e-08 w=6e-07 $X=19310 $Y=3881 $D=616
M736 308 225 b_bla_n<5> vss hvtnfet l=6e-08 w=6e-07 $X=19310 $Y=4141 $D=616
M737 t_bla_n<5> 226 308 vss hvtnfet l=6e-08 w=6e-07 $X=19310 $Y=46932 $D=616
M738 308 226 t_bla_n<5> vss hvtnfet l=6e-08 w=6e-07 $X=19310 $Y=47192 $D=616
M739 t_blb<5> 224 299 vss hvtnfet l=6e-08 w=6e-07 $X=19310 $Y=47872 $D=616
M740 299 224 t_blb<5> vss hvtnfet l=6e-08 w=6e-07 $X=19310 $Y=48132 $D=616
M741 609 vdd vss vss hvtnfet l=6e-08 w=6e-07 $X=19523 $Y=26159 $D=616
M742 223 221 vss vss hvtnfet l=6e-08 w=4e-07 $X=19635 $Y=4836 $D=616
M743 1117 b_cb<1> 221 vss hvtnfet l=6e-08 w=4e-07 $X=19635 $Y=11331 $D=616
M744 1118 221 219 vss hvtnfet l=6e-08 w=4e-07 $X=19635 $Y=12191 $D=616
M745 1119 222 220 vss hvtnfet l=6e-08 w=4e-07 $X=19635 $Y=38542 $D=616
M746 1120 t_cb<1> 222 vss hvtnfet l=6e-08 w=4e-07 $X=19635 $Y=39402 $D=616
M747 224 222 vss vss hvtnfet l=6e-08 w=4e-07 $X=19635 $Y=45897 $D=616
M748 612 vdd vss vss hvtnfet l=1.4e-07 w=2.1e-07 $X=19705 $Y=14550 $D=616
M749 613 vdd vss vss hvtnfet l=1.4e-07 w=2.1e-07 $X=19705 $Y=16760 $D=616
M750 vss vss vss vss hvtnfet l=7e-08 w=3.2e-07 $X=19710 $Y=33798 $D=616
M751 630 vdd vss vss hvtnfet l=6e-08 w=3e-07 $X=19730 $Y=17670 $D=616
M752 vss vss vss vss hvtnfet l=1.4e-07 w=7.5e-07 $X=19750 $Y=34593 $D=616
M753 vss vdd 609 vss hvtnfet l=6e-08 w=6e-07 $X=19783 $Y=26159 $D=616
M754 vss 11 223 vss hvtnfet l=6e-08 w=4e-07 $X=19895 $Y=4836 $D=616
M755 vss b_mb<1> 1117 vss hvtnfet l=6e-08 w=4e-07 $X=19895 $Y=11331 $D=616
M756 vss 13 1118 vss hvtnfet l=6e-08 w=4e-07 $X=19895 $Y=12191 $D=616
M757 vss 14 1119 vss hvtnfet l=6e-08 w=4e-07 $X=19895 $Y=38542 $D=616
M758 vss t_mb<1> 1120 vss hvtnfet l=6e-08 w=4e-07 $X=19895 $Y=39402 $D=616
M759 vss 11 224 vss hvtnfet l=6e-08 w=4e-07 $X=19895 $Y=45897 $D=616
M760 vss vdd 630 vss hvtnfet l=6e-08 w=3e-07 $X=19990 $Y=17670 $D=616
M761 vss vss vss vss hvtnfet l=8e-08 w=3.75e-07 $X=19990 $Y=33798 $D=616
M762 vss vss vss vss hvtnfet l=6e-08 w=3e-07 $X=20043 $Y=31223 $D=616
M763 vss vdd 612 vss hvtnfet l=1.4e-07 w=2.1e-07 $X=20045 $Y=14550 $D=616
M764 vss vdd 613 vss hvtnfet l=1.4e-07 w=2.1e-07 $X=20045 $Y=16760 $D=616
M765 vss vss vss vss hvtnfet l=1.4e-07 w=7.5e-07 $X=20090 $Y=34593 $D=616
M766 225 20 vss vss hvtnfet l=6e-08 w=4e-07 $X=20155 $Y=4836 $D=616
M767 1121 b_ma<1> vss vss hvtnfet l=6e-08 w=4e-07 $X=20155 $Y=11331 $D=616
M768 1122 22 vss vss hvtnfet l=6e-08 w=4e-07 $X=20155 $Y=12191 $D=616
M769 1123 23 vss vss hvtnfet l=6e-08 w=4e-07 $X=20155 $Y=38542 $D=616
M770 1124 t_ma<1> vss vss hvtnfet l=6e-08 w=4e-07 $X=20155 $Y=39402 $D=616
M771 226 20 vss vss hvtnfet l=6e-08 w=4e-07 $X=20155 $Y=45897 $D=616
M772 317 223 b_blb_n<5> vss hvtnfet l=6e-08 w=6e-07 $X=20200 $Y=2941 $D=616
M773 317 223 b_blb_n<5> vss hvtnfet l=6e-08 w=6e-07 $X=20200 $Y=3201 $D=616
M774 b_bla<5> 225 328 vss hvtnfet l=6e-08 w=6e-07 $X=20200 $Y=3881 $D=616
M775 b_bla<5> 225 328 vss hvtnfet l=6e-08 w=6e-07 $X=20200 $Y=4141 $D=616
M776 328 226 t_bla<5> vss hvtnfet l=6e-08 w=6e-07 $X=20200 $Y=46932 $D=616
M777 t_bla<5> 226 328 vss hvtnfet l=6e-08 w=6e-07 $X=20200 $Y=47192 $D=616
M778 t_blb_n<5> 224 317 vss hvtnfet l=6e-08 w=6e-07 $X=20200 $Y=47872 $D=616
M779 317 224 t_blb_n<5> vss hvtnfet l=6e-08 w=6e-07 $X=20200 $Y=48132 $D=616
M780 630 vdd vss vss hvtnfet l=6e-08 w=3e-07 $X=20250 $Y=17670 $D=616
M781 vss vss vss vss hvtnfet l=8e-08 w=3.75e-07 $X=20270 $Y=33798 $D=616
M782 vss vdd 636 vss hvtnfet l=6e-08 w=8e-07 $X=20293 $Y=26159 $D=616
M783 vss vss vss vss hvtnfet l=6e-08 w=3e-07 $X=20303 $Y=31223 $D=616
M784 vss 227 225 vss hvtnfet l=6e-08 w=4e-07 $X=20415 $Y=4836 $D=616
M785 227 b_ca<1> 1121 vss hvtnfet l=6e-08 w=4e-07 $X=20415 $Y=11331 $D=616
M786 229 227 1122 vss hvtnfet l=6e-08 w=4e-07 $X=20415 $Y=12191 $D=616
M787 230 228 1123 vss hvtnfet l=6e-08 w=4e-07 $X=20415 $Y=38542 $D=616
M788 228 t_ca<1> 1124 vss hvtnfet l=6e-08 w=4e-07 $X=20415 $Y=39402 $D=616
M789 vss 228 226 vss hvtnfet l=6e-08 w=4e-07 $X=20415 $Y=45897 $D=616
M790 vss vss vss vss hvtnfet l=1.4e-07 w=7.5e-07 $X=20430 $Y=34593 $D=616
M791 vss vdd 630 vss hvtnfet l=6e-08 w=3e-07 $X=20510 $Y=17670 $D=616
M792 vss vss vss vss hvtnfet l=8e-08 w=3.75e-07 $X=20550 $Y=33798 $D=616
M793 636 vdd vss vss hvtnfet l=6e-08 w=8e-07 $X=20553 $Y=26159 $D=616
M794 vss vss vss vss hvtnfet l=6e-08 w=3e-07 $X=20563 $Y=31223 $D=616
M795 628 vdd vss vss hvtnfet l=1.4e-07 w=2.1e-07 $X=20635 $Y=14550 $D=616
M796 629 vdd vss vss hvtnfet l=1.4e-07 w=2.1e-07 $X=20635 $Y=16760 $D=616
M797 vss vss vss vss hvtnfet l=6e-08 w=3.2e-07 $X=20680 $Y=19812 $D=616
M798 vss vss vss vss hvtnfet l=6e-08 w=3.2e-07 $X=20680 $Y=20072 $D=616
M799 vss vss vss vss hvtnfet l=6e-08 w=3.2e-07 $X=20680 $Y=21162 $D=616
M800 vss vss vss vss hvtnfet l=6e-08 w=3.2e-07 $X=20680 $Y=21422 $D=616
M801 vss vss vss vss hvtnfet l=6e-08 w=3.2e-07 $X=20680 $Y=21682 $D=616
M802 vss vss vss vss hvtnfet l=6e-08 w=3.2e-07 $X=20680 $Y=21942 $D=616
M803 vss vss vss vss hvtnfet l=6e-08 w=3.2e-07 $X=20680 $Y=22762 $D=616
M804 vss vss vss vss hvtnfet l=6e-08 w=3.2e-07 $X=20680 $Y=23879 $D=616
M805 vss vss vss vss hvtnfet l=6e-08 w=3.2e-07 $X=20680 $Y=24139 $D=616
M806 vss vss vss vss hvtnfet l=6e-08 w=3.2e-07 $X=20680 $Y=24399 $D=616
M807 vss vss vss vss hvtnfet l=6e-08 w=3.2e-07 $X=20680 $Y=24659 $D=616
M808 630 vdd vss vss hvtnfet l=6e-08 w=3e-07 $X=20770 $Y=17670 $D=616
M809 vss vss vss vss hvtnfet l=1.4e-07 w=7.5e-07 $X=20770 $Y=34593 $D=616
M810 631 vdd 636 vss hvtnfet l=6e-08 w=8e-07 $X=20813 $Y=26159 $D=616
M811 vss vss vss vss hvtnfet l=6e-08 w=3e-07 $X=20823 $Y=31223 $D=616
M812 vss vss vss vss hvtnfet l=8e-08 w=3.75e-07 $X=20830 $Y=33798 $D=616
M813 vss vdd 628 vss hvtnfet l=1.4e-07 w=2.1e-07 $X=20975 $Y=14550 $D=616
M814 vss vdd 629 vss hvtnfet l=1.4e-07 w=2.1e-07 $X=20975 $Y=16760 $D=616
M815 vss vdd 630 vss hvtnfet l=6e-08 w=3e-07 $X=21030 $Y=17670 $D=616
M816 636 vdd 631 vss hvtnfet l=6e-08 w=8e-07 $X=21073 $Y=26159 $D=616
M817 vss vss vss vss hvtnfet l=8e-08 w=3.75e-07 $X=21110 $Y=33798 $D=616
M818 vss vss vss vss hvtnfet l=1.4e-07 w=7.5e-07 $X=21110 $Y=34593 $D=616
M819 317 239 b_blb_n<4> vss hvtnfet l=6e-08 w=6e-07 $X=21220 $Y=2941 $D=616
M820 317 239 b_blb_n<4> vss hvtnfet l=6e-08 w=6e-07 $X=21220 $Y=3201 $D=616
M821 b_bla<4> 235 328 vss hvtnfet l=6e-08 w=6e-07 $X=21220 $Y=3881 $D=616
M822 b_bla<4> 235 328 vss hvtnfet l=6e-08 w=6e-07 $X=21220 $Y=4141 $D=616
M823 328 236 t_bla<4> vss hvtnfet l=6e-08 w=6e-07 $X=21220 $Y=46932 $D=616
M824 t_bla<4> 236 328 vss hvtnfet l=6e-08 w=6e-07 $X=21220 $Y=47192 $D=616
M825 t_blb_n<4> 240 317 vss hvtnfet l=6e-08 w=6e-07 $X=21220 $Y=47872 $D=616
M826 317 240 t_blb_n<4> vss hvtnfet l=6e-08 w=6e-07 $X=21220 $Y=48132 $D=616
M827 vss vss vss vss hvtnfet l=8e-08 w=3.75e-07 $X=21390 $Y=33798 $D=616
M828 vss vss vss vss hvtnfet l=1.4e-07 w=7.5e-07 $X=21450 $Y=34593 $D=616
M829 654 vdd vss vss hvtnfet l=6e-08 w=2.5e-07 $X=21540 $Y=17720 $D=616
M830 235 231 vss vss hvtnfet l=6e-08 w=4e-07 $X=21545 $Y=4836 $D=616
M831 1125 b_ca<0> 231 vss hvtnfet l=6e-08 w=4e-07 $X=21545 $Y=11331 $D=616
M832 1126 231 233 vss hvtnfet l=6e-08 w=4e-07 $X=21545 $Y=12191 $D=616
M833 1127 232 234 vss hvtnfet l=6e-08 w=4e-07 $X=21545 $Y=38542 $D=616
M834 1128 t_ca<0> 232 vss hvtnfet l=6e-08 w=4e-07 $X=21545 $Y=39402 $D=616
M835 236 232 vss vss hvtnfet l=6e-08 w=4e-07 $X=21545 $Y=45897 $D=616
M836 643 vdd vss vss hvtnfet l=6e-08 w=6e-07 $X=21593 $Y=26159 $D=616
M837 vss vss vss vss hvtnfet l=8e-08 w=3.75e-07 $X=21670 $Y=33798 $D=616
M838 vss vss vss vss hvtnfet l=6e-08 w=3e-07 $X=21733 $Y=31223 $D=616
M839 644 vdd vss vss hvtnfet l=6e-08 w=2e-07 $X=21745 $Y=21427 $D=616
M840 645 vdd vss vss hvtnfet l=6e-08 w=2e-07 $X=21745 $Y=23694 $D=616
M841 646 vdd vss vss hvtnfet l=6e-08 w=2e-07 $X=21745 $Y=24394 $D=616
M842 647 vdd vss vss hvtnfet l=6e-08 w=2e-07 $X=21745 $Y=24904 $D=616
M843 vss vss vss vss hvtnfet l=1.4e-07 w=7.5e-07 $X=21790 $Y=34593 $D=616
M844 vss vdd 654 vss hvtnfet l=6e-08 w=2.5e-07 $X=21800 $Y=17720 $D=616
M845 vss 20 235 vss hvtnfet l=6e-08 w=4e-07 $X=21805 $Y=4836 $D=616
M846 vss b_ma<1> 1125 vss hvtnfet l=6e-08 w=4e-07 $X=21805 $Y=11331 $D=616
M847 vss 22 1126 vss hvtnfet l=6e-08 w=4e-07 $X=21805 $Y=12191 $D=616
M848 vss 23 1127 vss hvtnfet l=6e-08 w=4e-07 $X=21805 $Y=38542 $D=616
M849 vss t_ma<1> 1128 vss hvtnfet l=6e-08 w=4e-07 $X=21805 $Y=39402 $D=616
M850 vss 20 236 vss hvtnfet l=6e-08 w=4e-07 $X=21805 $Y=45897 $D=616
M851 vss vdd 643 vss hvtnfet l=6e-08 w=6e-07 $X=21853 $Y=26159 $D=616
M852 vss vss vss vss hvtnfet l=8e-08 w=3.75e-07 $X=21950 $Y=33798 $D=616
M853 vss vss vss vss hvtnfet l=6e-08 w=3e-07 $X=21993 $Y=31223 $D=616
M854 654 vdd vss vss hvtnfet l=6e-08 w=2.5e-07 $X=22060 $Y=17720 $D=616
M855 239 11 vss vss hvtnfet l=6e-08 w=4e-07 $X=22065 $Y=4836 $D=616
M856 1129 b_mb<1> vss vss hvtnfet l=6e-08 w=4e-07 $X=22065 $Y=11331 $D=616
M857 1130 13 vss vss hvtnfet l=6e-08 w=4e-07 $X=22065 $Y=12191 $D=616
M858 1131 14 vss vss hvtnfet l=6e-08 w=4e-07 $X=22065 $Y=38542 $D=616
M859 1132 t_mb<1> vss vss hvtnfet l=6e-08 w=4e-07 $X=22065 $Y=39402 $D=616
M860 240 11 vss vss hvtnfet l=6e-08 w=4e-07 $X=22065 $Y=45897 $D=616
M861 299 239 b_blb<4> vss hvtnfet l=6e-08 w=6e-07 $X=22110 $Y=2941 $D=616
M862 299 239 b_blb<4> vss hvtnfet l=6e-08 w=6e-07 $X=22110 $Y=3201 $D=616
M863 308 235 b_bla_n<4> vss hvtnfet l=6e-08 w=6e-07 $X=22110 $Y=3881 $D=616
M864 308 235 b_bla_n<4> vss hvtnfet l=6e-08 w=6e-07 $X=22110 $Y=4141 $D=616
M865 t_bla_n<4> 236 308 vss hvtnfet l=6e-08 w=6e-07 $X=22110 $Y=46932 $D=616
M866 308 236 t_bla_n<4> vss hvtnfet l=6e-08 w=6e-07 $X=22110 $Y=47192 $D=616
M867 t_blb<4> 240 299 vss hvtnfet l=6e-08 w=6e-07 $X=22110 $Y=47872 $D=616
M868 299 240 t_blb<4> vss hvtnfet l=6e-08 w=6e-07 $X=22110 $Y=48132 $D=616
M869 vss vss vss vss hvtnfet l=1.4e-07 w=7.5e-07 $X=22130 $Y=34593 $D=616
M870 vss vss vss vss hvtnfet l=7e-08 w=3.2e-07 $X=22240 $Y=33798 $D=616
M871 vss vdd 654 vss hvtnfet l=6e-08 w=2.5e-07 $X=22320 $Y=17720 $D=616
M872 vss 237 239 vss hvtnfet l=6e-08 w=4e-07 $X=22325 $Y=4836 $D=616
M873 237 b_cb<0> 1129 vss hvtnfet l=6e-08 w=4e-07 $X=22325 $Y=11331 $D=616
M874 241 237 1130 vss hvtnfet l=6e-08 w=4e-07 $X=22325 $Y=12191 $D=616
M875 242 238 1131 vss hvtnfet l=6e-08 w=4e-07 $X=22325 $Y=38542 $D=616
M876 238 t_cb<0> 1132 vss hvtnfet l=6e-08 w=4e-07 $X=22325 $Y=39402 $D=616
M877 vss 238 240 vss hvtnfet l=6e-08 w=4e-07 $X=22325 $Y=45897 $D=616
M878 299 247 b_blb<3> vss hvtnfet l=6e-08 w=6e-07 $X=23130 $Y=2941 $D=616
M879 299 247 b_blb<3> vss hvtnfet l=6e-08 w=6e-07 $X=23130 $Y=3201 $D=616
M880 308 251 b_bla_n<3> vss hvtnfet l=6e-08 w=6e-07 $X=23130 $Y=3881 $D=616
M881 308 251 b_bla_n<3> vss hvtnfet l=6e-08 w=6e-07 $X=23130 $Y=4141 $D=616
M882 t_bla_n<3> 252 308 vss hvtnfet l=6e-08 w=6e-07 $X=23130 $Y=46932 $D=616
M883 308 252 t_bla_n<3> vss hvtnfet l=6e-08 w=6e-07 $X=23130 $Y=47192 $D=616
M884 t_blb<3> 248 299 vss hvtnfet l=6e-08 w=6e-07 $X=23130 $Y=47872 $D=616
M885 299 248 t_blb<3> vss hvtnfet l=6e-08 w=6e-07 $X=23130 $Y=48132 $D=616
M886 247 245 vss vss hvtnfet l=6e-08 w=4e-07 $X=23455 $Y=4836 $D=616
M887 1133 b_cb<3> 245 vss hvtnfet l=6e-08 w=4e-07 $X=23455 $Y=11331 $D=616
M888 1134 245 243 vss hvtnfet l=6e-08 w=4e-07 $X=23455 $Y=12191 $D=616
M889 1135 246 244 vss hvtnfet l=6e-08 w=4e-07 $X=23455 $Y=38542 $D=616
M890 1136 t_cb<3> 246 vss hvtnfet l=6e-08 w=4e-07 $X=23455 $Y=39402 $D=616
M891 248 246 vss vss hvtnfet l=6e-08 w=4e-07 $X=23455 $Y=45897 $D=616
M892 682 vdd vss vss hvtnfet l=6e-08 w=2.5e-07 $X=23460 $Y=17720 $D=616
M893 vss vss vss vss hvtnfet l=7e-08 w=3.2e-07 $X=23530 $Y=33798 $D=616
M894 vss vss vss vss hvtnfet l=1.4e-07 w=7.5e-07 $X=23570 $Y=34593 $D=616
M895 vss 11 247 vss hvtnfet l=6e-08 w=4e-07 $X=23715 $Y=4836 $D=616
M896 vss b_mb<0> 1133 vss hvtnfet l=6e-08 w=4e-07 $X=23715 $Y=11331 $D=616
M897 vss 13 1134 vss hvtnfet l=6e-08 w=4e-07 $X=23715 $Y=12191 $D=616
M898 vss 14 1135 vss hvtnfet l=6e-08 w=4e-07 $X=23715 $Y=38542 $D=616
M899 vss t_mb<0> 1136 vss hvtnfet l=6e-08 w=4e-07 $X=23715 $Y=39402 $D=616
M900 vss 11 248 vss hvtnfet l=6e-08 w=4e-07 $X=23715 $Y=45897 $D=616
M901 vss vdd 682 vss hvtnfet l=6e-08 w=2.5e-07 $X=23720 $Y=17720 $D=616
M902 vss vss vss vss hvtnfet l=6e-08 w=3e-07 $X=23787 $Y=31223 $D=616
M903 vss vss vss vss hvtnfet l=8e-08 w=3.75e-07 $X=23810 $Y=33798 $D=616
M904 667 vdd vss vss hvtnfet l=6e-08 w=2e-07 $X=23895 $Y=21427 $D=616
M905 668 vdd vss vss hvtnfet l=6e-08 w=2e-07 $X=23895 $Y=23694 $D=616
M906 669 vdd vss vss hvtnfet l=6e-08 w=2e-07 $X=23895 $Y=24394 $D=616
M907 670 vdd vss vss hvtnfet l=6e-08 w=2e-07 $X=23895 $Y=24904 $D=616
M908 vss vss vss vss hvtnfet l=1.4e-07 w=7.5e-07 $X=23910 $Y=34593 $D=616
M909 681 vdd vss vss hvtnfet l=6e-08 w=6e-07 $X=23927 $Y=26159 $D=616
M910 251 20 vss vss hvtnfet l=6e-08 w=4e-07 $X=23975 $Y=4836 $D=616
M911 1137 b_ma<0> vss vss hvtnfet l=6e-08 w=4e-07 $X=23975 $Y=11331 $D=616
M912 1138 22 vss vss hvtnfet l=6e-08 w=4e-07 $X=23975 $Y=12191 $D=616
M913 1139 23 vss vss hvtnfet l=6e-08 w=4e-07 $X=23975 $Y=38542 $D=616
M914 1140 t_ma<0> vss vss hvtnfet l=6e-08 w=4e-07 $X=23975 $Y=39402 $D=616
M915 252 20 vss vss hvtnfet l=6e-08 w=4e-07 $X=23975 $Y=45897 $D=616
M916 682 vdd vss vss hvtnfet l=6e-08 w=2.5e-07 $X=23980 $Y=17720 $D=616
M917 317 247 b_blb_n<3> vss hvtnfet l=6e-08 w=6e-07 $X=24020 $Y=2941 $D=616
M918 317 247 b_blb_n<3> vss hvtnfet l=6e-08 w=6e-07 $X=24020 $Y=3201 $D=616
M919 b_bla<3> 251 328 vss hvtnfet l=6e-08 w=6e-07 $X=24020 $Y=3881 $D=616
M920 b_bla<3> 251 328 vss hvtnfet l=6e-08 w=6e-07 $X=24020 $Y=4141 $D=616
M921 328 252 t_bla<3> vss hvtnfet l=6e-08 w=6e-07 $X=24020 $Y=46932 $D=616
M922 t_bla<3> 252 328 vss hvtnfet l=6e-08 w=6e-07 $X=24020 $Y=47192 $D=616
M923 t_blb_n<3> 248 317 vss hvtnfet l=6e-08 w=6e-07 $X=24020 $Y=47872 $D=616
M924 317 248 t_blb_n<3> vss hvtnfet l=6e-08 w=6e-07 $X=24020 $Y=48132 $D=616
M925 vss vss vss vss hvtnfet l=6e-08 w=3e-07 $X=24047 $Y=31223 $D=616
M926 vss vss vss vss hvtnfet l=8e-08 w=3.75e-07 $X=24090 $Y=33798 $D=616
M927 vss vdd 681 vss hvtnfet l=6e-08 w=6e-07 $X=24187 $Y=26159 $D=616
M928 vss 253 251 vss hvtnfet l=6e-08 w=4e-07 $X=24235 $Y=4836 $D=616
M929 253 b_ca<3> 1137 vss hvtnfet l=6e-08 w=4e-07 $X=24235 $Y=11331 $D=616
M930 257 253 1138 vss hvtnfet l=6e-08 w=4e-07 $X=24235 $Y=12191 $D=616
M931 258 254 1139 vss hvtnfet l=6e-08 w=4e-07 $X=24235 $Y=38542 $D=616
M932 254 t_ca<3> 1140 vss hvtnfet l=6e-08 w=4e-07 $X=24235 $Y=39402 $D=616
M933 vss 254 252 vss hvtnfet l=6e-08 w=4e-07 $X=24235 $Y=45897 $D=616
M934 vss vdd 682 vss hvtnfet l=6e-08 w=2.5e-07 $X=24240 $Y=17720 $D=616
M935 vss vss vss vss hvtnfet l=1.4e-07 w=7.5e-07 $X=24250 $Y=34593 $D=616
M936 vss vss vss vss hvtnfet l=8e-08 w=3.75e-07 $X=24370 $Y=33798 $D=616
M937 vss vss vss vss hvtnfet l=1.4e-07 w=7.5e-07 $X=24590 $Y=34593 $D=616
M938 vss vss vss vss hvtnfet l=8e-08 w=3.75e-07 $X=24650 $Y=33798 $D=616
M939 703 vdd 706 vss hvtnfet l=6e-08 w=8e-07 $X=24707 $Y=26159 $D=616
M940 697 vdd vss vss hvtnfet l=1.4e-07 w=2.1e-07 $X=24725 $Y=14550 $D=616
M941 698 vdd vss vss hvtnfet l=1.4e-07 w=2.1e-07 $X=24725 $Y=16760 $D=616
M942 713 vdd vss vss hvtnfet l=6e-08 w=3e-07 $X=24750 $Y=17670 $D=616
M943 vss vss vss vss hvtnfet l=6e-08 w=3.2e-07 $X=24840 $Y=19812 $D=616
M944 vss vss vss vss hvtnfet l=6e-08 w=3.2e-07 $X=24840 $Y=20072 $D=616
M945 vss vss vss vss hvtnfet l=6e-08 w=3.2e-07 $X=24840 $Y=21162 $D=616
M946 vss vss vss vss hvtnfet l=6e-08 w=3.2e-07 $X=24840 $Y=21422 $D=616
M947 vss vss vss vss hvtnfet l=6e-08 w=3.2e-07 $X=24840 $Y=21682 $D=616
M948 vss vss vss vss hvtnfet l=6e-08 w=3.2e-07 $X=24840 $Y=21942 $D=616
M949 vss vss vss vss hvtnfet l=6e-08 w=3.2e-07 $X=24840 $Y=22762 $D=616
M950 vss vss vss vss hvtnfet l=6e-08 w=3.2e-07 $X=24840 $Y=23879 $D=616
M951 vss vss vss vss hvtnfet l=6e-08 w=3.2e-07 $X=24840 $Y=24139 $D=616
M952 vss vss vss vss hvtnfet l=6e-08 w=3.2e-07 $X=24840 $Y=24399 $D=616
M953 vss vss vss vss hvtnfet l=6e-08 w=3.2e-07 $X=24840 $Y=24659 $D=616
M954 vss vss vss vss hvtnfet l=8e-08 w=3.75e-07 $X=24930 $Y=33798 $D=616
M955 vss vss vss vss hvtnfet l=1.4e-07 w=7.5e-07 $X=24930 $Y=34593 $D=616
M956 vss vss vss vss hvtnfet l=6e-08 w=3e-07 $X=24957 $Y=31223 $D=616
M957 706 vdd 703 vss hvtnfet l=6e-08 w=8e-07 $X=24967 $Y=26159 $D=616
M958 vss vdd 713 vss hvtnfet l=6e-08 w=3e-07 $X=25010 $Y=17670 $D=616
M959 317 267 b_blb_n<2> vss hvtnfet l=6e-08 w=6e-07 $X=25040 $Y=2941 $D=616
M960 317 267 b_blb_n<2> vss hvtnfet l=6e-08 w=6e-07 $X=25040 $Y=3201 $D=616
M961 b_bla<2> 263 328 vss hvtnfet l=6e-08 w=6e-07 $X=25040 $Y=3881 $D=616
M962 b_bla<2> 263 328 vss hvtnfet l=6e-08 w=6e-07 $X=25040 $Y=4141 $D=616
M963 328 264 t_bla<2> vss hvtnfet l=6e-08 w=6e-07 $X=25040 $Y=46932 $D=616
M964 t_bla<2> 264 328 vss hvtnfet l=6e-08 w=6e-07 $X=25040 $Y=47192 $D=616
M965 t_blb_n<2> 268 317 vss hvtnfet l=6e-08 w=6e-07 $X=25040 $Y=47872 $D=616
M966 317 268 t_blb_n<2> vss hvtnfet l=6e-08 w=6e-07 $X=25040 $Y=48132 $D=616
M967 vss vdd 697 vss hvtnfet l=1.4e-07 w=2.1e-07 $X=25065 $Y=14550 $D=616
M968 vss vdd 698 vss hvtnfet l=1.4e-07 w=2.1e-07 $X=25065 $Y=16760 $D=616
M969 vss vss vss vss hvtnfet l=8e-08 w=3.75e-07 $X=25210 $Y=33798 $D=616
M970 vss vss vss vss hvtnfet l=6e-08 w=3e-07 $X=25217 $Y=31223 $D=616
M971 vss vdd 706 vss hvtnfet l=6e-08 w=8e-07 $X=25227 $Y=26159 $D=616
M972 713 vdd vss vss hvtnfet l=6e-08 w=3e-07 $X=25270 $Y=17670 $D=616
M973 vss vss vss vss hvtnfet l=1.4e-07 w=7.5e-07 $X=25270 $Y=34593 $D=616
M974 263 259 vss vss hvtnfet l=6e-08 w=4e-07 $X=25365 $Y=4836 $D=616
M975 1141 b_ca<2> 259 vss hvtnfet l=6e-08 w=4e-07 $X=25365 $Y=11331 $D=616
M976 1142 259 261 vss hvtnfet l=6e-08 w=4e-07 $X=25365 $Y=12191 $D=616
M977 1143 260 262 vss hvtnfet l=6e-08 w=4e-07 $X=25365 $Y=38542 $D=616
M978 1144 t_ca<2> 260 vss hvtnfet l=6e-08 w=4e-07 $X=25365 $Y=39402 $D=616
M979 264 260 vss vss hvtnfet l=6e-08 w=4e-07 $X=25365 $Y=45897 $D=616
M980 vss vss vss vss hvtnfet l=6e-08 w=3e-07 $X=25477 $Y=31223 $D=616
M981 706 vdd vss vss hvtnfet l=6e-08 w=8e-07 $X=25487 $Y=26159 $D=616
M982 vss vss vss vss hvtnfet l=8e-08 w=3.75e-07 $X=25490 $Y=33798 $D=616
M983 vss vdd 713 vss hvtnfet l=6e-08 w=3e-07 $X=25530 $Y=17670 $D=616
M984 vss vss vss vss hvtnfet l=1.4e-07 w=7.5e-07 $X=25610 $Y=34593 $D=616
M985 vss 20 263 vss hvtnfet l=6e-08 w=4e-07 $X=25625 $Y=4836 $D=616
M986 vss b_ma<0> 1141 vss hvtnfet l=6e-08 w=4e-07 $X=25625 $Y=11331 $D=616
M987 vss 22 1142 vss hvtnfet l=6e-08 w=4e-07 $X=25625 $Y=12191 $D=616
M988 vss 23 1143 vss hvtnfet l=6e-08 w=4e-07 $X=25625 $Y=38542 $D=616
M989 vss t_ma<0> 1144 vss hvtnfet l=6e-08 w=4e-07 $X=25625 $Y=39402 $D=616
M990 vss 20 264 vss hvtnfet l=6e-08 w=4e-07 $X=25625 $Y=45897 $D=616
M991 711 vdd vss vss hvtnfet l=1.4e-07 w=2.1e-07 $X=25655 $Y=14550 $D=616
M992 712 vdd vss vss hvtnfet l=1.4e-07 w=2.1e-07 $X=25655 $Y=16760 $D=616
M993 vss vss vss vss hvtnfet l=6e-08 w=3e-07 $X=25737 $Y=31223 $D=616
M994 vss vss vss vss hvtnfet l=8e-08 w=3.75e-07 $X=25770 $Y=33798 $D=616
M995 713 vdd vss vss hvtnfet l=6e-08 w=3e-07 $X=25790 $Y=17670 $D=616
M996 267 11 vss vss hvtnfet l=6e-08 w=4e-07 $X=25885 $Y=4836 $D=616
M997 1145 b_mb<0> vss vss hvtnfet l=6e-08 w=4e-07 $X=25885 $Y=11331 $D=616
M998 1146 13 vss vss hvtnfet l=6e-08 w=4e-07 $X=25885 $Y=12191 $D=616
M999 1147 14 vss vss hvtnfet l=6e-08 w=4e-07 $X=25885 $Y=38542 $D=616
M1000 1148 t_mb<0> vss vss hvtnfet l=6e-08 w=4e-07 $X=25885 $Y=39402 $D=616
M1001 268 11 vss vss hvtnfet l=6e-08 w=4e-07 $X=25885 $Y=45897 $D=616
M1002 299 267 b_blb<2> vss hvtnfet l=6e-08 w=6e-07 $X=25930 $Y=2941 $D=616
M1003 299 267 b_blb<2> vss hvtnfet l=6e-08 w=6e-07 $X=25930 $Y=3201 $D=616
M1004 308 263 b_bla_n<2> vss hvtnfet l=6e-08 w=6e-07 $X=25930 $Y=3881 $D=616
M1005 308 263 b_bla_n<2> vss hvtnfet l=6e-08 w=6e-07 $X=25930 $Y=4141 $D=616
M1006 t_bla_n<2> 264 308 vss hvtnfet l=6e-08 w=6e-07 $X=25930 $Y=46932 $D=616
M1007 308 264 t_bla_n<2> vss hvtnfet l=6e-08 w=6e-07 $X=25930 $Y=47192 $D=616
M1008 t_blb<2> 268 299 vss hvtnfet l=6e-08 w=6e-07 $X=25930 $Y=47872 $D=616
M1009 299 268 t_blb<2> vss hvtnfet l=6e-08 w=6e-07 $X=25930 $Y=48132 $D=616
M1010 vss vss vss vss hvtnfet l=1.4e-07 w=7.5e-07 $X=25950 $Y=34593 $D=616
M1011 vss vdd 711 vss hvtnfet l=1.4e-07 w=2.1e-07 $X=25995 $Y=14550 $D=616
M1012 vss vdd 712 vss hvtnfet l=1.4e-07 w=2.1e-07 $X=25995 $Y=16760 $D=616
M1013 720 vdd vss vss hvtnfet l=6e-08 w=6e-07 $X=25997 $Y=26159 $D=616
M1014 vss vdd 713 vss hvtnfet l=6e-08 w=3e-07 $X=26050 $Y=17670 $D=616
M1015 vss vss vss vss hvtnfet l=7e-08 w=3.2e-07 $X=26060 $Y=33798 $D=616
M1016 vss 265 267 vss hvtnfet l=6e-08 w=4e-07 $X=26145 $Y=4836 $D=616
M1017 265 b_cb<2> 1145 vss hvtnfet l=6e-08 w=4e-07 $X=26145 $Y=11331 $D=616
M1018 269 265 1146 vss hvtnfet l=6e-08 w=4e-07 $X=26145 $Y=12191 $D=616
M1019 270 266 1147 vss hvtnfet l=6e-08 w=4e-07 $X=26145 $Y=38542 $D=616
M1020 266 t_cb<2> 1148 vss hvtnfet l=6e-08 w=4e-07 $X=26145 $Y=39402 $D=616
M1021 vss 266 268 vss hvtnfet l=6e-08 w=4e-07 $X=26145 $Y=45897 $D=616
M1022 vss vdd 720 vss hvtnfet l=6e-08 w=6e-07 $X=26257 $Y=26159 $D=616
M1023 299 275 b_blb<1> vss hvtnfet l=6e-08 w=6e-07 $X=26950 $Y=2941 $D=616
M1024 299 275 b_blb<1> vss hvtnfet l=6e-08 w=6e-07 $X=26950 $Y=3201 $D=616
M1025 308 277 b_bla_n<1> vss hvtnfet l=6e-08 w=6e-07 $X=26950 $Y=3881 $D=616
M1026 308 277 b_bla_n<1> vss hvtnfet l=6e-08 w=6e-07 $X=26950 $Y=4141 $D=616
M1027 t_bla_n<1> 278 308 vss hvtnfet l=6e-08 w=6e-07 $X=26950 $Y=46932 $D=616
M1028 308 278 t_bla_n<1> vss hvtnfet l=6e-08 w=6e-07 $X=26950 $Y=47192 $D=616
M1029 t_blb<1> 276 299 vss hvtnfet l=6e-08 w=6e-07 $X=26950 $Y=47872 $D=616
M1030 299 276 t_blb<1> vss hvtnfet l=6e-08 w=6e-07 $X=26950 $Y=48132 $D=616
M1031 733 vdd vss vss hvtnfet l=6e-08 w=6e-07 $X=27163 $Y=26159 $D=616
M1032 275 273 vss vss hvtnfet l=6e-08 w=4e-07 $X=27275 $Y=4836 $D=616
M1033 1149 b_cb<1> 273 vss hvtnfet l=6e-08 w=4e-07 $X=27275 $Y=11331 $D=616
M1034 1150 273 271 vss hvtnfet l=6e-08 w=4e-07 $X=27275 $Y=12191 $D=616
M1035 1151 274 272 vss hvtnfet l=6e-08 w=4e-07 $X=27275 $Y=38542 $D=616
M1036 1152 t_cb<1> 274 vss hvtnfet l=6e-08 w=4e-07 $X=27275 $Y=39402 $D=616
M1037 276 274 vss vss hvtnfet l=6e-08 w=4e-07 $X=27275 $Y=45897 $D=616
M1038 736 vdd vss vss hvtnfet l=1.4e-07 w=2.1e-07 $X=27345 $Y=14550 $D=616
M1039 737 vdd vss vss hvtnfet l=1.4e-07 w=2.1e-07 $X=27345 $Y=16760 $D=616
M1040 vss vss vss vss hvtnfet l=7e-08 w=3.2e-07 $X=27350 $Y=33798 $D=616
M1041 754 vdd vss vss hvtnfet l=6e-08 w=3e-07 $X=27370 $Y=17670 $D=616
M1042 vss vss vss vss hvtnfet l=1.4e-07 w=7.5e-07 $X=27390 $Y=34593 $D=616
M1043 vss vdd 733 vss hvtnfet l=6e-08 w=6e-07 $X=27423 $Y=26159 $D=616
M1044 vss 11 275 vss hvtnfet l=6e-08 w=4e-07 $X=27535 $Y=4836 $D=616
M1045 vss b_mb<0> 1149 vss hvtnfet l=6e-08 w=4e-07 $X=27535 $Y=11331 $D=616
M1046 vss 13 1150 vss hvtnfet l=6e-08 w=4e-07 $X=27535 $Y=12191 $D=616
M1047 vss 14 1151 vss hvtnfet l=6e-08 w=4e-07 $X=27535 $Y=38542 $D=616
M1048 vss t_mb<0> 1152 vss hvtnfet l=6e-08 w=4e-07 $X=27535 $Y=39402 $D=616
M1049 vss 11 276 vss hvtnfet l=6e-08 w=4e-07 $X=27535 $Y=45897 $D=616
M1050 vss vdd 754 vss hvtnfet l=6e-08 w=3e-07 $X=27630 $Y=17670 $D=616
M1051 vss vss vss vss hvtnfet l=8e-08 w=3.75e-07 $X=27630 $Y=33798 $D=616
M1052 vss vss vss vss hvtnfet l=6e-08 w=3e-07 $X=27683 $Y=31223 $D=616
M1053 vss vdd 736 vss hvtnfet l=1.4e-07 w=2.1e-07 $X=27685 $Y=14550 $D=616
M1054 vss vdd 737 vss hvtnfet l=1.4e-07 w=2.1e-07 $X=27685 $Y=16760 $D=616
M1055 vss vss vss vss hvtnfet l=1.4e-07 w=7.5e-07 $X=27730 $Y=34593 $D=616
M1056 277 20 vss vss hvtnfet l=6e-08 w=4e-07 $X=27795 $Y=4836 $D=616
M1057 1153 b_ma<0> vss vss hvtnfet l=6e-08 w=4e-07 $X=27795 $Y=11331 $D=616
M1058 1154 22 vss vss hvtnfet l=6e-08 w=4e-07 $X=27795 $Y=12191 $D=616
M1059 1155 23 vss vss hvtnfet l=6e-08 w=4e-07 $X=27795 $Y=38542 $D=616
M1060 1156 t_ma<0> vss vss hvtnfet l=6e-08 w=4e-07 $X=27795 $Y=39402 $D=616
M1061 278 20 vss vss hvtnfet l=6e-08 w=4e-07 $X=27795 $Y=45897 $D=616
M1062 317 275 b_blb_n<1> vss hvtnfet l=6e-08 w=6e-07 $X=27840 $Y=2941 $D=616
M1063 317 275 b_blb_n<1> vss hvtnfet l=6e-08 w=6e-07 $X=27840 $Y=3201 $D=616
M1064 b_bla<1> 277 328 vss hvtnfet l=6e-08 w=6e-07 $X=27840 $Y=3881 $D=616
M1065 b_bla<1> 277 328 vss hvtnfet l=6e-08 w=6e-07 $X=27840 $Y=4141 $D=616
M1066 328 278 t_bla<1> vss hvtnfet l=6e-08 w=6e-07 $X=27840 $Y=46932 $D=616
M1067 t_bla<1> 278 328 vss hvtnfet l=6e-08 w=6e-07 $X=27840 $Y=47192 $D=616
M1068 t_blb_n<1> 276 317 vss hvtnfet l=6e-08 w=6e-07 $X=27840 $Y=47872 $D=616
M1069 317 276 t_blb_n<1> vss hvtnfet l=6e-08 w=6e-07 $X=27840 $Y=48132 $D=616
M1070 754 vdd vss vss hvtnfet l=6e-08 w=3e-07 $X=27890 $Y=17670 $D=616
M1071 vss vss vss vss hvtnfet l=8e-08 w=3.75e-07 $X=27910 $Y=33798 $D=616
M1072 vss vdd 760 vss hvtnfet l=6e-08 w=8e-07 $X=27933 $Y=26159 $D=616
M1073 vss vss vss vss hvtnfet l=6e-08 w=3e-07 $X=27943 $Y=31223 $D=616
M1074 vss 279 277 vss hvtnfet l=6e-08 w=4e-07 $X=28055 $Y=4836 $D=616
M1075 279 b_ca<1> 1153 vss hvtnfet l=6e-08 w=4e-07 $X=28055 $Y=11331 $D=616
M1076 281 279 1154 vss hvtnfet l=6e-08 w=4e-07 $X=28055 $Y=12191 $D=616
M1077 282 280 1155 vss hvtnfet l=6e-08 w=4e-07 $X=28055 $Y=38542 $D=616
M1078 280 t_ca<1> 1156 vss hvtnfet l=6e-08 w=4e-07 $X=28055 $Y=39402 $D=616
M1079 vss 280 278 vss hvtnfet l=6e-08 w=4e-07 $X=28055 $Y=45897 $D=616
M1080 vss vss vss vss hvtnfet l=1.4e-07 w=7.5e-07 $X=28070 $Y=34593 $D=616
M1081 vss vdd 754 vss hvtnfet l=6e-08 w=3e-07 $X=28150 $Y=17670 $D=616
M1082 vss vss vss vss hvtnfet l=8e-08 w=3.75e-07 $X=28190 $Y=33798 $D=616
M1083 760 vdd vss vss hvtnfet l=6e-08 w=8e-07 $X=28193 $Y=26159 $D=616
M1084 vss vss vss vss hvtnfet l=6e-08 w=3e-07 $X=28203 $Y=31223 $D=616
M1085 752 vdd vss vss hvtnfet l=1.4e-07 w=2.1e-07 $X=28275 $Y=14550 $D=616
M1086 753 vdd vss vss hvtnfet l=1.4e-07 w=2.1e-07 $X=28275 $Y=16760 $D=616
M1087 vss vss vss vss hvtnfet l=6e-08 w=3.2e-07 $X=28320 $Y=19812 $D=616
M1088 vss vss vss vss hvtnfet l=6e-08 w=3.2e-07 $X=28320 $Y=20072 $D=616
M1089 vss vss vss vss hvtnfet l=6e-08 w=3.2e-07 $X=28320 $Y=21162 $D=616
M1090 vss vss vss vss hvtnfet l=6e-08 w=3.2e-07 $X=28320 $Y=21422 $D=616
M1091 vss vss vss vss hvtnfet l=6e-08 w=3.2e-07 $X=28320 $Y=21682 $D=616
M1092 vss vss vss vss hvtnfet l=6e-08 w=3.2e-07 $X=28320 $Y=21942 $D=616
M1093 vss vss vss vss hvtnfet l=6e-08 w=3.2e-07 $X=28320 $Y=22762 $D=616
M1094 vss vss vss vss hvtnfet l=6e-08 w=3.2e-07 $X=28320 $Y=23879 $D=616
M1095 vss vss vss vss hvtnfet l=6e-08 w=3.2e-07 $X=28320 $Y=24139 $D=616
M1096 vss vss vss vss hvtnfet l=6e-08 w=3.2e-07 $X=28320 $Y=24399 $D=616
M1097 vss vss vss vss hvtnfet l=6e-08 w=3.2e-07 $X=28320 $Y=24659 $D=616
M1098 754 vdd vss vss hvtnfet l=6e-08 w=3e-07 $X=28410 $Y=17670 $D=616
M1099 vss vss vss vss hvtnfet l=1.4e-07 w=7.5e-07 $X=28410 $Y=34593 $D=616
M1100 755 vdd 760 vss hvtnfet l=6e-08 w=8e-07 $X=28453 $Y=26159 $D=616
M1101 vss vss vss vss hvtnfet l=6e-08 w=3e-07 $X=28463 $Y=31223 $D=616
M1102 vss vss vss vss hvtnfet l=8e-08 w=3.75e-07 $X=28470 $Y=33798 $D=616
M1103 vss vdd 752 vss hvtnfet l=1.4e-07 w=2.1e-07 $X=28615 $Y=14550 $D=616
M1104 vss vdd 753 vss hvtnfet l=1.4e-07 w=2.1e-07 $X=28615 $Y=16760 $D=616
M1105 vss vdd 754 vss hvtnfet l=6e-08 w=3e-07 $X=28670 $Y=17670 $D=616
M1106 760 vdd 755 vss hvtnfet l=6e-08 w=8e-07 $X=28713 $Y=26159 $D=616
M1107 vss vss vss vss hvtnfet l=8e-08 w=3.75e-07 $X=28750 $Y=33798 $D=616
M1108 vss vss vss vss hvtnfet l=1.4e-07 w=7.5e-07 $X=28750 $Y=34593 $D=616
M1109 317 291 b_blb_n<0> vss hvtnfet l=6e-08 w=6e-07 $X=28860 $Y=2941 $D=616
M1110 317 291 b_blb_n<0> vss hvtnfet l=6e-08 w=6e-07 $X=28860 $Y=3201 $D=616
M1111 b_bla<0> 287 328 vss hvtnfet l=6e-08 w=6e-07 $X=28860 $Y=3881 $D=616
M1112 b_bla<0> 287 328 vss hvtnfet l=6e-08 w=6e-07 $X=28860 $Y=4141 $D=616
M1113 328 288 t_bla<0> vss hvtnfet l=6e-08 w=6e-07 $X=28860 $Y=46932 $D=616
M1114 t_bla<0> 288 328 vss hvtnfet l=6e-08 w=6e-07 $X=28860 $Y=47192 $D=616
M1115 t_blb_n<0> 292 317 vss hvtnfet l=6e-08 w=6e-07 $X=28860 $Y=47872 $D=616
M1116 317 292 t_blb_n<0> vss hvtnfet l=6e-08 w=6e-07 $X=28860 $Y=48132 $D=616
M1117 vss vss vss vss hvtnfet l=8e-08 w=3.75e-07 $X=29030 $Y=33798 $D=616
M1118 vss vss vss vss hvtnfet l=1.4e-07 w=7.5e-07 $X=29090 $Y=34593 $D=616
M1119 778 vdd vss vss hvtnfet l=6e-08 w=2.5e-07 $X=29180 $Y=17720 $D=616
M1120 287 283 vss vss hvtnfet l=6e-08 w=4e-07 $X=29185 $Y=4836 $D=616
M1121 1157 b_ca<0> 283 vss hvtnfet l=6e-08 w=4e-07 $X=29185 $Y=11331 $D=616
M1122 1158 283 285 vss hvtnfet l=6e-08 w=4e-07 $X=29185 $Y=12191 $D=616
M1123 1159 284 286 vss hvtnfet l=6e-08 w=4e-07 $X=29185 $Y=38542 $D=616
M1124 1160 t_ca<0> 284 vss hvtnfet l=6e-08 w=4e-07 $X=29185 $Y=39402 $D=616
M1125 288 284 vss vss hvtnfet l=6e-08 w=4e-07 $X=29185 $Y=45897 $D=616
M1126 767 vdd vss vss hvtnfet l=6e-08 w=6e-07 $X=29233 $Y=26159 $D=616
M1127 vss vss vss vss hvtnfet l=8e-08 w=3.75e-07 $X=29310 $Y=33798 $D=616
M1128 vss vss vss vss hvtnfet l=6e-08 w=3e-07 $X=29373 $Y=31223 $D=616
M1129 768 vdd vss vss hvtnfet l=6e-08 w=2e-07 $X=29385 $Y=21427 $D=616
M1130 769 vdd vss vss hvtnfet l=6e-08 w=2e-07 $X=29385 $Y=23694 $D=616
M1131 770 vdd vss vss hvtnfet l=6e-08 w=2e-07 $X=29385 $Y=24394 $D=616
M1132 771 vdd vss vss hvtnfet l=6e-08 w=2e-07 $X=29385 $Y=24904 $D=616
M1133 vss vss vss vss hvtnfet l=1.4e-07 w=7.5e-07 $X=29430 $Y=34593 $D=616
M1134 vss vdd 778 vss hvtnfet l=6e-08 w=2.5e-07 $X=29440 $Y=17720 $D=616
M1135 vss 20 287 vss hvtnfet l=6e-08 w=4e-07 $X=29445 $Y=4836 $D=616
M1136 vss b_ma<0> 1157 vss hvtnfet l=6e-08 w=4e-07 $X=29445 $Y=11331 $D=616
M1137 vss 22 1158 vss hvtnfet l=6e-08 w=4e-07 $X=29445 $Y=12191 $D=616
M1138 vss 23 1159 vss hvtnfet l=6e-08 w=4e-07 $X=29445 $Y=38542 $D=616
M1139 vss t_ma<0> 1160 vss hvtnfet l=6e-08 w=4e-07 $X=29445 $Y=39402 $D=616
M1140 vss 20 288 vss hvtnfet l=6e-08 w=4e-07 $X=29445 $Y=45897 $D=616
M1141 vss vdd 767 vss hvtnfet l=6e-08 w=6e-07 $X=29493 $Y=26159 $D=616
M1142 vss vss vss vss hvtnfet l=8e-08 w=3.75e-07 $X=29590 $Y=33798 $D=616
M1143 vss vss vss vss hvtnfet l=6e-08 w=3e-07 $X=29633 $Y=31223 $D=616
M1144 778 vdd vss vss hvtnfet l=6e-08 w=2.5e-07 $X=29700 $Y=17720 $D=616
M1145 291 11 vss vss hvtnfet l=6e-08 w=4e-07 $X=29705 $Y=4836 $D=616
M1146 1161 b_mb<0> vss vss hvtnfet l=6e-08 w=4e-07 $X=29705 $Y=11331 $D=616
M1147 1162 13 vss vss hvtnfet l=6e-08 w=4e-07 $X=29705 $Y=12191 $D=616
M1148 1163 14 vss vss hvtnfet l=6e-08 w=4e-07 $X=29705 $Y=38542 $D=616
M1149 1164 t_mb<0> vss vss hvtnfet l=6e-08 w=4e-07 $X=29705 $Y=39402 $D=616
M1150 292 11 vss vss hvtnfet l=6e-08 w=4e-07 $X=29705 $Y=45897 $D=616
M1151 299 291 b_blb<0> vss hvtnfet l=6e-08 w=6e-07 $X=29750 $Y=2941 $D=616
M1152 299 291 b_blb<0> vss hvtnfet l=6e-08 w=6e-07 $X=29750 $Y=3201 $D=616
M1153 308 287 b_bla_n<0> vss hvtnfet l=6e-08 w=6e-07 $X=29750 $Y=3881 $D=616
M1154 308 287 b_bla_n<0> vss hvtnfet l=6e-08 w=6e-07 $X=29750 $Y=4141 $D=616
M1155 t_bla_n<0> 288 308 vss hvtnfet l=6e-08 w=6e-07 $X=29750 $Y=46932 $D=616
M1156 308 288 t_bla_n<0> vss hvtnfet l=6e-08 w=6e-07 $X=29750 $Y=47192 $D=616
M1157 t_blb<0> 292 299 vss hvtnfet l=6e-08 w=6e-07 $X=29750 $Y=47872 $D=616
M1158 299 292 t_blb<0> vss hvtnfet l=6e-08 w=6e-07 $X=29750 $Y=48132 $D=616
M1159 vss vss vss vss hvtnfet l=1.4e-07 w=7.5e-07 $X=29770 $Y=34593 $D=616
M1160 vss vss vss vss hvtnfet l=7e-08 w=3.2e-07 $X=29880 $Y=33798 $D=616
M1161 vss vdd 778 vss hvtnfet l=6e-08 w=2.5e-07 $X=29960 $Y=17720 $D=616
M1162 vss 289 291 vss hvtnfet l=6e-08 w=4e-07 $X=29965 $Y=4836 $D=616
M1163 289 b_cb<0> 1161 vss hvtnfet l=6e-08 w=4e-07 $X=29965 $Y=11331 $D=616
M1164 293 289 1162 vss hvtnfet l=6e-08 w=4e-07 $X=29965 $Y=12191 $D=616
M1165 294 290 1163 vss hvtnfet l=6e-08 w=4e-07 $X=29965 $Y=38542 $D=616
M1166 290 t_cb<0> 1164 vss hvtnfet l=6e-08 w=4e-07 $X=29965 $Y=39402 $D=616
M1167 vss 290 292 vss hvtnfet l=6e-08 w=4e-07 $X=29965 $Y=45897 $D=616
M1168 b_blb_n<15> 2 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=187 $Y=-170 $D=636
M1169 t_blb_n<15> 3 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=187 $Y=50503 $D=636
M1170 vdd vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=205 $Y=35893 $D=636
M1171 296 5 b_blb<15> vdd hvtpfet l=6e-08 w=3e-07 $X=210 $Y=1094 $D=636
M1172 b_blb<15> 5 296 vdd hvtpfet l=6e-08 w=3e-07 $X=210 $Y=1354 $D=636
M1173 b_blb_n<15> 5 297 vdd hvtpfet l=6e-08 w=3e-07 $X=210 $Y=1864 $D=636
M1174 297 5 b_blb_n<15> vdd hvtpfet l=6e-08 w=3e-07 $X=210 $Y=2124 $D=636
M1175 t_blb_n<15> 6 297 vdd hvtpfet l=6e-08 w=3e-07 $X=210 $Y=48949 $D=636
M1176 297 6 t_blb_n<15> vdd hvtpfet l=6e-08 w=3e-07 $X=210 $Y=49209 $D=636
M1177 296 6 t_blb<15> vdd hvtpfet l=6e-08 w=3e-07 $X=210 $Y=49719 $D=636
M1178 t_blb<15> 6 296 vdd hvtpfet l=6e-08 w=3e-07 $X=210 $Y=49979 $D=636
M1179 302 vdd vdd vdd hvtpfet l=6e-08 w=4e-07 $X=255 $Y=21427 $D=636
M1180 303 vdd vdd vdd hvtpfet l=6e-08 w=4e-07 $X=255 $Y=23694 $D=636
M1181 304 vdd vdd vdd hvtpfet l=6e-08 w=4e-07 $X=255 $Y=24394 $D=636
M1182 305 vdd vdd vdd hvtpfet l=6e-08 w=4e-07 $X=255 $Y=24904 $D=636
M1183 b_blb<15> 2 b_blb_n<15> vdd hvtpfet l=6e-08 w=8e-07 $X=447 $Y=-170 $D=636
M1184 t_blb<15> 3 t_blb_n<15> vdd hvtpfet l=6e-08 w=8e-07 $X=447 $Y=50503 $D=636
M1185 1169 5 8 vdd hvtpfet l=6e-08 w=8e-07 $X=535 $Y=5556 $D=636
M1186 5 b_cb<3> vdd vdd hvtpfet l=6e-08 w=4e-07 $X=535 $Y=10611 $D=636
M1187 2 5 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=535 $Y=12911 $D=636
M1188 3 6 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=535 $Y=37822 $D=636
M1189 6 t_cb<3> vdd vdd hvtpfet l=6e-08 w=4e-07 $X=535 $Y=40122 $D=636
M1190 1170 6 9 vdd hvtpfet l=6e-08 w=8e-07 $X=535 $Y=44777 $D=636
M1191 319 vdd vdd vdd hvtpfet l=6e-08 w=5e-07 $X=540 $Y=18290 $D=636
M1192 vdd vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=650 $Y=35893 $D=636
M1193 vdd vdd vdd vdd hvtpfet l=1e-07 w=2e-07 $X=685 $Y=36723 $D=636
M1194 vdd 2 b_blb<15> vdd hvtpfet l=6e-08 w=8e-07 $X=707 $Y=-170 $D=636
M1195 vdd 3 t_blb<15> vdd hvtpfet l=6e-08 w=8e-07 $X=707 $Y=50503 $D=636
M1196 vdd 11 1169 vdd hvtpfet l=6e-08 w=8e-07 $X=795 $Y=5556 $D=636
M1197 vdd b_mb<3> 5 vdd hvtpfet l=6e-08 w=4e-07 $X=795 $Y=10611 $D=636
M1198 vdd 13 2 vdd hvtpfet l=6e-08 w=4e-07 $X=795 $Y=12911 $D=636
M1199 vdd 14 3 vdd hvtpfet l=6e-08 w=4e-07 $X=795 $Y=37822 $D=636
M1200 vdd t_mb<3> 6 vdd hvtpfet l=6e-08 w=4e-07 $X=795 $Y=40122 $D=636
M1201 vdd 11 1170 vdd hvtpfet l=6e-08 w=8e-07 $X=795 $Y=44777 $D=636
M1202 vdd vdd 319 vdd hvtpfet l=6e-08 w=5e-07 $X=800 $Y=18290 $D=636
M1203 vdd vdd vdd vdd hvtpfet l=6e-08 w=6e-07 $X=867 $Y=29008 $D=636
M1204 vdd vdd vdd vdd hvtpfet l=1e-07 w=2e-07 $X=985 $Y=36723 $D=636
M1205 vdd vdd vdd vdd hvtpfet l=7e-08 w=3.2e-07 $X=990 $Y=32628 $D=636
M1206 vdd vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=990 $Y=35893 $D=636
M1207 1171 20 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=1055 $Y=5556 $D=636
M1208 18 b_ma<3> vdd vdd hvtpfet l=6e-08 w=4e-07 $X=1055 $Y=10611 $D=636
M1209 25 22 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=1055 $Y=12911 $D=636
M1210 26 23 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=1055 $Y=37822 $D=636
M1211 19 t_ma<3> vdd vdd hvtpfet l=6e-08 w=4e-07 $X=1055 $Y=40122 $D=636
M1212 1172 20 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=1055 $Y=44777 $D=636
M1213 319 vdd vdd vdd hvtpfet l=6e-08 w=5e-07 $X=1060 $Y=18290 $D=636
M1214 vdd vdd vdd vdd hvtpfet l=6e-08 w=6e-07 $X=1127 $Y=29008 $D=636
M1215 b_bla_n<15> 25 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=1143 $Y=-170 $D=636
M1216 t_bla_n<15> 26 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=1143 $Y=50503 $D=636
M1217 vdd vdd 318 vdd hvtpfet l=6e-08 w=6e-07 $X=1267 $Y=27488 $D=636
M1218 vdd vdd vdd vdd hvtpfet l=7e-08 w=3.2e-07 $X=1280 $Y=32628 $D=636
M1219 vdd vdd vdd vdd hvtpfet l=1e-07 w=2e-07 $X=1285 $Y=36723 $D=636
M1220 16 18 1171 vdd hvtpfet l=6e-08 w=8e-07 $X=1315 $Y=5556 $D=636
M1221 vdd b_ca<3> 18 vdd hvtpfet l=6e-08 w=4e-07 $X=1315 $Y=10611 $D=636
M1222 vdd 18 25 vdd hvtpfet l=6e-08 w=4e-07 $X=1315 $Y=12911 $D=636
M1223 vdd 19 26 vdd hvtpfet l=6e-08 w=4e-07 $X=1315 $Y=37822 $D=636
M1224 vdd t_ca<3> 19 vdd hvtpfet l=6e-08 w=4e-07 $X=1315 $Y=40122 $D=636
M1225 17 19 1172 vdd hvtpfet l=6e-08 w=8e-07 $X=1315 $Y=44777 $D=636
M1226 vdd vdd 319 vdd hvtpfet l=6e-08 w=5e-07 $X=1320 $Y=18290 $D=636
M1227 vdd vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=1330 $Y=35893 $D=636
M1228 325 18 b_bla<15> vdd hvtpfet l=6e-08 w=3e-07 $X=1400 $Y=1094 $D=636
M1229 b_bla<15> 18 325 vdd hvtpfet l=6e-08 w=3e-07 $X=1400 $Y=1354 $D=636
M1230 b_bla_n<15> 18 326 vdd hvtpfet l=6e-08 w=3e-07 $X=1400 $Y=1864 $D=636
M1231 326 18 b_bla_n<15> vdd hvtpfet l=6e-08 w=3e-07 $X=1400 $Y=2124 $D=636
M1232 t_bla_n<15> 19 326 vdd hvtpfet l=6e-08 w=3e-07 $X=1400 $Y=48949 $D=636
M1233 326 19 t_bla_n<15> vdd hvtpfet l=6e-08 w=3e-07 $X=1400 $Y=49209 $D=636
M1234 325 19 t_bla<15> vdd hvtpfet l=6e-08 w=3e-07 $X=1400 $Y=49719 $D=636
M1235 t_bla<15> 19 325 vdd hvtpfet l=6e-08 w=3e-07 $X=1400 $Y=49979 $D=636
M1236 b_bla<15> 25 b_bla_n<15> vdd hvtpfet l=6e-08 w=8e-07 $X=1403 $Y=-170 $D=636
M1237 t_bla<15> 26 t_bla_n<15> vdd hvtpfet l=6e-08 w=8e-07 $X=1403 $Y=50503 $D=636
M1238 vdd vdd vdd vdd hvtpfet l=1e-07 w=6e-07 $X=1560 $Y=32628 $D=636
M1239 vdd vdd vdd vdd hvtpfet l=1e-07 w=2e-07 $X=1585 $Y=36723 $D=636
M1240 vdd 25 b_bla<15> vdd hvtpfet l=6e-08 w=8e-07 $X=1663 $Y=-170 $D=636
M1241 vdd 26 t_bla<15> vdd hvtpfet l=6e-08 w=8e-07 $X=1663 $Y=50503 $D=636
M1242 vdd vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=1670 $Y=35893 $D=636
M1243 343 vdd vdd vdd hvtpfet l=6e-08 w=8e-07 $X=1787 $Y=27288 $D=636
M1244 337 vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=1805 $Y=15090 $D=636
M1245 338 vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=1805 $Y=16110 $D=636
M1246 353 vdd vdd vdd hvtpfet l=6e-08 w=6e-07 $X=1830 $Y=18290 $D=636
M1247 vdd vdd vdd vdd hvtpfet l=1e-07 w=6e-07 $X=1860 $Y=32628 $D=636
M1248 vdd vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=2010 $Y=35893 $D=636
M1249 vdd vdd vdd vdd hvtpfet l=6e-08 w=6e-07 $X=2037 $Y=29008 $D=636
M1250 vdd vdd 343 vdd hvtpfet l=6e-08 w=8e-07 $X=2047 $Y=27288 $D=636
M1251 vdd vdd 353 vdd hvtpfet l=6e-08 w=6e-07 $X=2090 $Y=18290 $D=636
M1252 b_bla<14> 33 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=2097 $Y=-170 $D=636
M1253 t_bla<14> 34 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=2097 $Y=50503 $D=636
M1254 325 30 b_bla<14> vdd hvtpfet l=6e-08 w=3e-07 $X=2120 $Y=1094 $D=636
M1255 b_bla<14> 30 325 vdd hvtpfet l=6e-08 w=3e-07 $X=2120 $Y=1354 $D=636
M1256 b_bla_n<14> 30 326 vdd hvtpfet l=6e-08 w=3e-07 $X=2120 $Y=1864 $D=636
M1257 326 30 b_bla_n<14> vdd hvtpfet l=6e-08 w=3e-07 $X=2120 $Y=2124 $D=636
M1258 t_bla_n<14> 31 326 vdd hvtpfet l=6e-08 w=3e-07 $X=2120 $Y=48949 $D=636
M1259 326 31 t_bla_n<14> vdd hvtpfet l=6e-08 w=3e-07 $X=2120 $Y=49209 $D=636
M1260 325 31 t_bla<14> vdd hvtpfet l=6e-08 w=3e-07 $X=2120 $Y=49719 $D=636
M1261 t_bla<14> 31 325 vdd hvtpfet l=6e-08 w=3e-07 $X=2120 $Y=49979 $D=636
M1262 vdd vdd vdd vdd hvtpfet l=1e-07 w=2e-07 $X=2135 $Y=36723 $D=636
M1263 vdd vdd 337 vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=2145 $Y=15090 $D=636
M1264 vdd vdd 338 vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=2145 $Y=16110 $D=636
M1265 vdd vdd vdd vdd hvtpfet l=1e-07 w=6e-07 $X=2160 $Y=32628 $D=636
M1266 vdd vdd vdd vdd hvtpfet l=6e-08 w=6e-07 $X=2297 $Y=29008 $D=636
M1267 343 vdd vdd vdd hvtpfet l=6e-08 w=8e-07 $X=2307 $Y=27288 $D=636
M1268 353 vdd vdd vdd hvtpfet l=6e-08 w=6e-07 $X=2350 $Y=18290 $D=636
M1269 vdd vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=2350 $Y=35893 $D=636
M1270 b_bla_n<14> 33 b_bla<14> vdd hvtpfet l=6e-08 w=8e-07 $X=2357 $Y=-170 $D=636
M1271 t_bla_n<14> 34 t_bla<14> vdd hvtpfet l=6e-08 w=8e-07 $X=2357 $Y=50503 $D=636
M1272 vdd vdd vdd vdd hvtpfet l=1e-07 w=2e-07 $X=2435 $Y=36723 $D=636
M1273 1177 30 35 vdd hvtpfet l=6e-08 w=8e-07 $X=2445 $Y=5556 $D=636
M1274 30 b_ca<2> vdd vdd hvtpfet l=6e-08 w=4e-07 $X=2445 $Y=10611 $D=636
M1275 33 30 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=2445 $Y=12911 $D=636
M1276 34 31 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=2445 $Y=37822 $D=636
M1277 31 t_ca<2> vdd vdd hvtpfet l=6e-08 w=4e-07 $X=2445 $Y=40122 $D=636
M1278 1178 31 36 vdd hvtpfet l=6e-08 w=8e-07 $X=2445 $Y=44777 $D=636
M1279 vdd vdd vdd vdd hvtpfet l=7e-08 w=3.2e-07 $X=2470 $Y=32628 $D=636
M1280 vdd vdd vdd vdd hvtpfet l=6e-08 w=6e-07 $X=2557 $Y=29008 $D=636
M1281 vdd vdd 343 vdd hvtpfet l=6e-08 w=8e-07 $X=2567 $Y=27288 $D=636
M1282 vdd vdd 353 vdd hvtpfet l=6e-08 w=6e-07 $X=2610 $Y=18290 $D=636
M1283 vdd 33 b_bla_n<14> vdd hvtpfet l=6e-08 w=8e-07 $X=2617 $Y=-170 $D=636
M1284 vdd 34 t_bla_n<14> vdd hvtpfet l=6e-08 w=8e-07 $X=2617 $Y=50503 $D=636
M1285 vdd vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=2690 $Y=35893 $D=636
M1286 vdd 20 1177 vdd hvtpfet l=6e-08 w=8e-07 $X=2705 $Y=5556 $D=636
M1287 vdd b_ma<3> 30 vdd hvtpfet l=6e-08 w=4e-07 $X=2705 $Y=10611 $D=636
M1288 vdd 22 33 vdd hvtpfet l=6e-08 w=4e-07 $X=2705 $Y=12911 $D=636
M1289 vdd 23 34 vdd hvtpfet l=6e-08 w=4e-07 $X=2705 $Y=37822 $D=636
M1290 vdd t_ma<3> 31 vdd hvtpfet l=6e-08 w=4e-07 $X=2705 $Y=40122 $D=636
M1291 vdd 20 1178 vdd hvtpfet l=6e-08 w=8e-07 $X=2705 $Y=44777 $D=636
M1292 351 vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=2735 $Y=15090 $D=636
M1293 352 vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=2735 $Y=16110 $D=636
M1294 vdd vdd vdd vdd hvtpfet l=1e-07 w=2e-07 $X=2735 $Y=36723 $D=636
M1295 vdd vdd vdd vdd hvtpfet l=7e-08 w=3.2e-07 $X=2760 $Y=32628 $D=636
M1296 vdd vdd vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=2806 $Y=19812 $D=636
M1297 vdd vdd vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=2806 $Y=20072 $D=636
M1298 vdd vdd vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=2806 $Y=21162 $D=636
M1299 vdd vdd vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=2806 $Y=21422 $D=636
M1300 vdd vdd vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=2806 $Y=21682 $D=636
M1301 vdd vdd vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=2806 $Y=21942 $D=636
M1302 vdd vdd vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=2806 $Y=22762 $D=636
M1303 vdd vdd vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=2806 $Y=23879 $D=636
M1304 vdd vdd vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=2806 $Y=24139 $D=636
M1305 vdd vdd vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=2806 $Y=24399 $D=636
M1306 vdd vdd vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=2806 $Y=24659 $D=636
M1307 vdd vdd vdd vdd hvtpfet l=6e-08 w=6e-07 $X=2817 $Y=29008 $D=636
M1308 353 vdd vdd vdd hvtpfet l=6e-08 w=6e-07 $X=2870 $Y=18290 $D=636
M1309 1179 11 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=2965 $Y=5556 $D=636
M1310 37 b_mb<3> vdd vdd hvtpfet l=6e-08 w=4e-07 $X=2965 $Y=10611 $D=636
M1311 41 13 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=2965 $Y=12911 $D=636
M1312 42 14 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=2965 $Y=37822 $D=636
M1313 38 t_mb<3> vdd vdd hvtpfet l=6e-08 w=4e-07 $X=2965 $Y=40122 $D=636
M1314 1180 11 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=2965 $Y=44777 $D=636
M1315 vdd vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=3030 $Y=35893 $D=636
M1316 vdd vdd vdd vdd hvtpfet l=1e-07 w=2e-07 $X=3035 $Y=36723 $D=636
M1317 b_blb<14> 41 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=3053 $Y=-170 $D=636
M1318 t_blb<14> 42 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=3053 $Y=50503 $D=636
M1319 vdd vdd 351 vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=3075 $Y=15090 $D=636
M1320 vdd vdd 352 vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=3075 $Y=16110 $D=636
M1321 360 vdd vdd vdd hvtpfet l=6e-08 w=6e-07 $X=3077 $Y=27488 $D=636
M1322 vdd vdd 353 vdd hvtpfet l=6e-08 w=6e-07 $X=3130 $Y=18290 $D=636
M1323 39 37 1179 vdd hvtpfet l=6e-08 w=8e-07 $X=3225 $Y=5556 $D=636
M1324 vdd b_cb<2> 37 vdd hvtpfet l=6e-08 w=4e-07 $X=3225 $Y=10611 $D=636
M1325 vdd 37 41 vdd hvtpfet l=6e-08 w=4e-07 $X=3225 $Y=12911 $D=636
M1326 vdd 38 42 vdd hvtpfet l=6e-08 w=4e-07 $X=3225 $Y=37822 $D=636
M1327 vdd t_cb<2> 38 vdd hvtpfet l=6e-08 w=4e-07 $X=3225 $Y=40122 $D=636
M1328 40 38 1180 vdd hvtpfet l=6e-08 w=8e-07 $X=3225 $Y=44777 $D=636
M1329 296 37 b_blb<14> vdd hvtpfet l=6e-08 w=3e-07 $X=3310 $Y=1094 $D=636
M1330 b_blb<14> 37 296 vdd hvtpfet l=6e-08 w=3e-07 $X=3310 $Y=1354 $D=636
M1331 b_blb_n<14> 37 297 vdd hvtpfet l=6e-08 w=3e-07 $X=3310 $Y=1864 $D=636
M1332 297 37 b_blb_n<14> vdd hvtpfet l=6e-08 w=3e-07 $X=3310 $Y=2124 $D=636
M1333 t_blb_n<14> 38 297 vdd hvtpfet l=6e-08 w=3e-07 $X=3310 $Y=48949 $D=636
M1334 297 38 t_blb_n<14> vdd hvtpfet l=6e-08 w=3e-07 $X=3310 $Y=49209 $D=636
M1335 296 38 t_blb<14> vdd hvtpfet l=6e-08 w=3e-07 $X=3310 $Y=49719 $D=636
M1336 t_blb<14> 38 296 vdd hvtpfet l=6e-08 w=3e-07 $X=3310 $Y=49979 $D=636
M1337 b_blb_n<14> 41 b_blb<14> vdd hvtpfet l=6e-08 w=8e-07 $X=3313 $Y=-170 $D=636
M1338 t_blb_n<14> 42 t_blb<14> vdd hvtpfet l=6e-08 w=8e-07 $X=3313 $Y=50503 $D=636
M1339 vdd vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=3475 $Y=35893 $D=636
M1340 vdd 41 b_blb_n<14> vdd hvtpfet l=6e-08 w=8e-07 $X=3573 $Y=-170 $D=636
M1341 vdd 42 t_blb_n<14> vdd hvtpfet l=6e-08 w=8e-07 $X=3573 $Y=50503 $D=636
M1342 b_blb_n<13> 45 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=4007 $Y=-170 $D=636
M1343 t_blb_n<13> 46 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=4007 $Y=50503 $D=636
M1344 vdd vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=4025 $Y=35893 $D=636
M1345 296 48 b_blb<13> vdd hvtpfet l=6e-08 w=3e-07 $X=4030 $Y=1094 $D=636
M1346 b_blb<13> 48 296 vdd hvtpfet l=6e-08 w=3e-07 $X=4030 $Y=1354 $D=636
M1347 b_blb_n<13> 48 297 vdd hvtpfet l=6e-08 w=3e-07 $X=4030 $Y=1864 $D=636
M1348 297 48 b_blb_n<13> vdd hvtpfet l=6e-08 w=3e-07 $X=4030 $Y=2124 $D=636
M1349 t_blb_n<13> 49 297 vdd hvtpfet l=6e-08 w=3e-07 $X=4030 $Y=48949 $D=636
M1350 297 49 t_blb_n<13> vdd hvtpfet l=6e-08 w=3e-07 $X=4030 $Y=49209 $D=636
M1351 296 49 t_blb<13> vdd hvtpfet l=6e-08 w=3e-07 $X=4030 $Y=49719 $D=636
M1352 t_blb<13> 49 296 vdd hvtpfet l=6e-08 w=3e-07 $X=4030 $Y=49979 $D=636
M1353 b_blb<13> 45 b_blb_n<13> vdd hvtpfet l=6e-08 w=8e-07 $X=4267 $Y=-170 $D=636
M1354 t_blb<13> 46 t_blb_n<13> vdd hvtpfet l=6e-08 w=8e-07 $X=4267 $Y=50503 $D=636
M1355 1185 48 51 vdd hvtpfet l=6e-08 w=8e-07 $X=4355 $Y=5556 $D=636
M1356 48 b_cb<1> vdd vdd hvtpfet l=6e-08 w=4e-07 $X=4355 $Y=10611 $D=636
M1357 45 48 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=4355 $Y=12911 $D=636
M1358 46 49 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=4355 $Y=37822 $D=636
M1359 49 t_cb<1> vdd vdd hvtpfet l=6e-08 w=4e-07 $X=4355 $Y=40122 $D=636
M1360 1186 49 52 vdd hvtpfet l=6e-08 w=8e-07 $X=4355 $Y=44777 $D=636
M1361 376 vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=4425 $Y=15090 $D=636
M1362 377 vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=4425 $Y=16110 $D=636
M1363 394 vdd vdd vdd hvtpfet l=6e-08 w=6e-07 $X=4450 $Y=18290 $D=636
M1364 vdd vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=4470 $Y=35893 $D=636
M1365 vdd vdd 373 vdd hvtpfet l=6e-08 w=6e-07 $X=4503 $Y=27488 $D=636
M1366 vdd vdd vdd vdd hvtpfet l=1e-07 w=2e-07 $X=4505 $Y=36723 $D=636
M1367 vdd vdd vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=4514 $Y=19812 $D=636
M1368 vdd vdd vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=4514 $Y=20072 $D=636
M1369 vdd vdd vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=4514 $Y=21162 $D=636
M1370 vdd vdd vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=4514 $Y=21422 $D=636
M1371 vdd vdd vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=4514 $Y=21682 $D=636
M1372 vdd vdd vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=4514 $Y=21942 $D=636
M1373 vdd vdd vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=4514 $Y=22762 $D=636
M1374 vdd vdd vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=4514 $Y=23879 $D=636
M1375 vdd vdd vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=4514 $Y=24139 $D=636
M1376 vdd vdd vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=4514 $Y=24399 $D=636
M1377 vdd vdd vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=4514 $Y=24659 $D=636
M1378 vdd 45 b_blb<13> vdd hvtpfet l=6e-08 w=8e-07 $X=4527 $Y=-170 $D=636
M1379 vdd 46 t_blb<13> vdd hvtpfet l=6e-08 w=8e-07 $X=4527 $Y=50503 $D=636
M1380 vdd 11 1185 vdd hvtpfet l=6e-08 w=8e-07 $X=4615 $Y=5556 $D=636
M1381 vdd b_mb<3> 48 vdd hvtpfet l=6e-08 w=4e-07 $X=4615 $Y=10611 $D=636
M1382 vdd 13 45 vdd hvtpfet l=6e-08 w=4e-07 $X=4615 $Y=12911 $D=636
M1383 vdd 14 46 vdd hvtpfet l=6e-08 w=4e-07 $X=4615 $Y=37822 $D=636
M1384 vdd t_mb<3> 49 vdd hvtpfet l=6e-08 w=4e-07 $X=4615 $Y=40122 $D=636
M1385 vdd 11 1186 vdd hvtpfet l=6e-08 w=8e-07 $X=4615 $Y=44777 $D=636
M1386 vdd vdd 394 vdd hvtpfet l=6e-08 w=6e-07 $X=4710 $Y=18290 $D=636
M1387 vdd vdd vdd vdd hvtpfet l=6e-08 w=6e-07 $X=4763 $Y=29008 $D=636
M1388 vdd vdd 376 vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=4765 $Y=15090 $D=636
M1389 vdd vdd 377 vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=4765 $Y=16110 $D=636
M1390 vdd vdd vdd vdd hvtpfet l=1e-07 w=2e-07 $X=4805 $Y=36723 $D=636
M1391 vdd vdd vdd vdd hvtpfet l=7e-08 w=3.2e-07 $X=4810 $Y=32628 $D=636
M1392 vdd vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=4810 $Y=35893 $D=636
M1393 1187 20 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=4875 $Y=5556 $D=636
M1394 55 b_ma<3> vdd vdd hvtpfet l=6e-08 w=4e-07 $X=4875 $Y=10611 $D=636
M1395 57 22 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=4875 $Y=12911 $D=636
M1396 58 23 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=4875 $Y=37822 $D=636
M1397 56 t_ma<3> vdd vdd hvtpfet l=6e-08 w=4e-07 $X=4875 $Y=40122 $D=636
M1398 1188 20 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=4875 $Y=44777 $D=636
M1399 b_bla_n<13> 57 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=4963 $Y=-170 $D=636
M1400 t_bla_n<13> 58 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=4963 $Y=50503 $D=636
M1401 394 vdd vdd vdd hvtpfet l=6e-08 w=6e-07 $X=4970 $Y=18290 $D=636
M1402 395 vdd vdd vdd hvtpfet l=6e-08 w=8e-07 $X=5013 $Y=27288 $D=636
M1403 vdd vdd vdd vdd hvtpfet l=6e-08 w=6e-07 $X=5023 $Y=29008 $D=636
M1404 vdd vdd vdd vdd hvtpfet l=7e-08 w=3.2e-07 $X=5100 $Y=32628 $D=636
M1405 vdd vdd vdd vdd hvtpfet l=1e-07 w=2e-07 $X=5105 $Y=36723 $D=636
M1406 53 55 1187 vdd hvtpfet l=6e-08 w=8e-07 $X=5135 $Y=5556 $D=636
M1407 vdd b_ca<1> 55 vdd hvtpfet l=6e-08 w=4e-07 $X=5135 $Y=10611 $D=636
M1408 vdd 55 57 vdd hvtpfet l=6e-08 w=4e-07 $X=5135 $Y=12911 $D=636
M1409 vdd 56 58 vdd hvtpfet l=6e-08 w=4e-07 $X=5135 $Y=37822 $D=636
M1410 vdd t_ca<1> 56 vdd hvtpfet l=6e-08 w=4e-07 $X=5135 $Y=40122 $D=636
M1411 54 56 1188 vdd hvtpfet l=6e-08 w=8e-07 $X=5135 $Y=44777 $D=636
M1412 vdd vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=5150 $Y=35893 $D=636
M1413 325 55 b_bla<13> vdd hvtpfet l=6e-08 w=3e-07 $X=5220 $Y=1094 $D=636
M1414 b_bla<13> 55 325 vdd hvtpfet l=6e-08 w=3e-07 $X=5220 $Y=1354 $D=636
M1415 b_bla_n<13> 55 326 vdd hvtpfet l=6e-08 w=3e-07 $X=5220 $Y=1864 $D=636
M1416 326 55 b_bla_n<13> vdd hvtpfet l=6e-08 w=3e-07 $X=5220 $Y=2124 $D=636
M1417 t_bla_n<13> 56 326 vdd hvtpfet l=6e-08 w=3e-07 $X=5220 $Y=48949 $D=636
M1418 326 56 t_bla_n<13> vdd hvtpfet l=6e-08 w=3e-07 $X=5220 $Y=49209 $D=636
M1419 325 56 t_bla<13> vdd hvtpfet l=6e-08 w=3e-07 $X=5220 $Y=49719 $D=636
M1420 t_bla<13> 56 325 vdd hvtpfet l=6e-08 w=3e-07 $X=5220 $Y=49979 $D=636
M1421 b_bla<13> 57 b_bla_n<13> vdd hvtpfet l=6e-08 w=8e-07 $X=5223 $Y=-170 $D=636
M1422 t_bla<13> 58 t_bla_n<13> vdd hvtpfet l=6e-08 w=8e-07 $X=5223 $Y=50503 $D=636
M1423 vdd vdd 394 vdd hvtpfet l=6e-08 w=6e-07 $X=5230 $Y=18290 $D=636
M1424 vdd vdd 395 vdd hvtpfet l=6e-08 w=8e-07 $X=5273 $Y=27288 $D=636
M1425 vdd vdd vdd vdd hvtpfet l=6e-08 w=6e-07 $X=5283 $Y=29008 $D=636
M1426 392 vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=5355 $Y=15090 $D=636
M1427 393 vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=5355 $Y=16110 $D=636
M1428 vdd vdd vdd vdd hvtpfet l=1e-07 w=6e-07 $X=5380 $Y=32628 $D=636
M1429 vdd vdd vdd vdd hvtpfet l=1e-07 w=2e-07 $X=5405 $Y=36723 $D=636
M1430 vdd 57 b_bla<13> vdd hvtpfet l=6e-08 w=8e-07 $X=5483 $Y=-170 $D=636
M1431 vdd 58 t_bla<13> vdd hvtpfet l=6e-08 w=8e-07 $X=5483 $Y=50503 $D=636
M1432 394 vdd vdd vdd hvtpfet l=6e-08 w=6e-07 $X=5490 $Y=18290 $D=636
M1433 vdd vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=5490 $Y=35893 $D=636
M1434 395 vdd vdd vdd hvtpfet l=6e-08 w=8e-07 $X=5533 $Y=27288 $D=636
M1435 vdd vdd vdd vdd hvtpfet l=6e-08 w=6e-07 $X=5543 $Y=29008 $D=636
M1436 vdd vdd vdd vdd hvtpfet l=1e-07 w=6e-07 $X=5680 $Y=32628 $D=636
M1437 vdd vdd 392 vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=5695 $Y=15090 $D=636
M1438 vdd vdd 393 vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=5695 $Y=16110 $D=636
M1439 vdd vdd 394 vdd hvtpfet l=6e-08 w=6e-07 $X=5750 $Y=18290 $D=636
M1440 vdd vdd 395 vdd hvtpfet l=6e-08 w=8e-07 $X=5793 $Y=27288 $D=636
M1441 vdd vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=5830 $Y=35893 $D=636
M1442 b_bla<12> 65 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=5917 $Y=-170 $D=636
M1443 t_bla<12> 66 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=5917 $Y=50503 $D=636
M1444 325 62 b_bla<12> vdd hvtpfet l=6e-08 w=3e-07 $X=5940 $Y=1094 $D=636
M1445 b_bla<12> 62 325 vdd hvtpfet l=6e-08 w=3e-07 $X=5940 $Y=1354 $D=636
M1446 b_bla_n<12> 62 326 vdd hvtpfet l=6e-08 w=3e-07 $X=5940 $Y=1864 $D=636
M1447 326 62 b_bla_n<12> vdd hvtpfet l=6e-08 w=3e-07 $X=5940 $Y=2124 $D=636
M1448 t_bla_n<12> 63 326 vdd hvtpfet l=6e-08 w=3e-07 $X=5940 $Y=48949 $D=636
M1449 326 63 t_bla_n<12> vdd hvtpfet l=6e-08 w=3e-07 $X=5940 $Y=49209 $D=636
M1450 325 63 t_bla<12> vdd hvtpfet l=6e-08 w=3e-07 $X=5940 $Y=49719 $D=636
M1451 t_bla<12> 63 325 vdd hvtpfet l=6e-08 w=3e-07 $X=5940 $Y=49979 $D=636
M1452 vdd vdd vdd vdd hvtpfet l=1e-07 w=2e-07 $X=5955 $Y=36723 $D=636
M1453 vdd vdd vdd vdd hvtpfet l=1e-07 w=6e-07 $X=5980 $Y=32628 $D=636
M1454 vdd vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=6170 $Y=35893 $D=636
M1455 b_bla_n<12> 65 b_bla<12> vdd hvtpfet l=6e-08 w=8e-07 $X=6177 $Y=-170 $D=636
M1456 t_bla_n<12> 66 t_bla<12> vdd hvtpfet l=6e-08 w=8e-07 $X=6177 $Y=50503 $D=636
M1457 vdd vdd vdd vdd hvtpfet l=1e-07 w=2e-07 $X=6255 $Y=36723 $D=636
M1458 418 vdd vdd vdd hvtpfet l=6e-08 w=5e-07 $X=6260 $Y=18290 $D=636
M1459 1193 62 67 vdd hvtpfet l=6e-08 w=8e-07 $X=6265 $Y=5556 $D=636
M1460 62 b_ca<0> vdd vdd hvtpfet l=6e-08 w=4e-07 $X=6265 $Y=10611 $D=636
M1461 65 62 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=6265 $Y=12911 $D=636
M1462 66 63 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=6265 $Y=37822 $D=636
M1463 63 t_ca<0> vdd vdd hvtpfet l=6e-08 w=4e-07 $X=6265 $Y=40122 $D=636
M1464 1194 63 68 vdd hvtpfet l=6e-08 w=8e-07 $X=6265 $Y=44777 $D=636
M1465 vdd vdd vdd vdd hvtpfet l=7e-08 w=3.2e-07 $X=6290 $Y=32628 $D=636
M1466 407 vdd vdd vdd hvtpfet l=6e-08 w=6e-07 $X=6313 $Y=27488 $D=636
M1467 vdd 65 b_bla_n<12> vdd hvtpfet l=6e-08 w=8e-07 $X=6437 $Y=-170 $D=636
M1468 vdd 66 t_bla_n<12> vdd hvtpfet l=6e-08 w=8e-07 $X=6437 $Y=50503 $D=636
M1469 vdd vdd vdd vdd hvtpfet l=6e-08 w=6e-07 $X=6453 $Y=29008 $D=636
M1470 vdd vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=6510 $Y=35893 $D=636
M1471 vdd vdd 418 vdd hvtpfet l=6e-08 w=5e-07 $X=6520 $Y=18290 $D=636
M1472 vdd 20 1193 vdd hvtpfet l=6e-08 w=8e-07 $X=6525 $Y=5556 $D=636
M1473 vdd b_ma<3> 62 vdd hvtpfet l=6e-08 w=4e-07 $X=6525 $Y=10611 $D=636
M1474 vdd 22 65 vdd hvtpfet l=6e-08 w=4e-07 $X=6525 $Y=12911 $D=636
M1475 vdd 23 66 vdd hvtpfet l=6e-08 w=4e-07 $X=6525 $Y=37822 $D=636
M1476 vdd t_ma<3> 63 vdd hvtpfet l=6e-08 w=4e-07 $X=6525 $Y=40122 $D=636
M1477 vdd 20 1194 vdd hvtpfet l=6e-08 w=8e-07 $X=6525 $Y=44777 $D=636
M1478 vdd vdd vdd vdd hvtpfet l=1e-07 w=2e-07 $X=6555 $Y=36723 $D=636
M1479 vdd vdd vdd vdd hvtpfet l=7e-08 w=3.2e-07 $X=6580 $Y=32628 $D=636
M1480 vdd vdd vdd vdd hvtpfet l=6e-08 w=6e-07 $X=6713 $Y=29008 $D=636
M1481 418 vdd vdd vdd hvtpfet l=6e-08 w=5e-07 $X=6780 $Y=18290 $D=636
M1482 1195 11 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=6785 $Y=5556 $D=636
M1483 69 b_mb<3> vdd vdd hvtpfet l=6e-08 w=4e-07 $X=6785 $Y=10611 $D=636
M1484 73 13 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=6785 $Y=12911 $D=636
M1485 74 14 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=6785 $Y=37822 $D=636
M1486 70 t_mb<3> vdd vdd hvtpfet l=6e-08 w=4e-07 $X=6785 $Y=40122 $D=636
M1487 1196 11 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=6785 $Y=44777 $D=636
M1488 vdd vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=6850 $Y=35893 $D=636
M1489 vdd vdd vdd vdd hvtpfet l=1e-07 w=2e-07 $X=6855 $Y=36723 $D=636
M1490 b_blb<12> 73 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=6873 $Y=-170 $D=636
M1491 t_blb<12> 74 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=6873 $Y=50503 $D=636
M1492 408 vdd vdd vdd hvtpfet l=6e-08 w=4e-07 $X=6985 $Y=21427 $D=636
M1493 409 vdd vdd vdd hvtpfet l=6e-08 w=4e-07 $X=6985 $Y=23694 $D=636
M1494 410 vdd vdd vdd hvtpfet l=6e-08 w=4e-07 $X=6985 $Y=24394 $D=636
M1495 411 vdd vdd vdd hvtpfet l=6e-08 w=4e-07 $X=6985 $Y=24904 $D=636
M1496 vdd vdd 418 vdd hvtpfet l=6e-08 w=5e-07 $X=7040 $Y=18290 $D=636
M1497 71 69 1195 vdd hvtpfet l=6e-08 w=8e-07 $X=7045 $Y=5556 $D=636
M1498 vdd b_cb<0> 69 vdd hvtpfet l=6e-08 w=4e-07 $X=7045 $Y=10611 $D=636
M1499 vdd 69 73 vdd hvtpfet l=6e-08 w=4e-07 $X=7045 $Y=12911 $D=636
M1500 vdd 70 74 vdd hvtpfet l=6e-08 w=4e-07 $X=7045 $Y=37822 $D=636
M1501 vdd t_cb<0> 70 vdd hvtpfet l=6e-08 w=4e-07 $X=7045 $Y=40122 $D=636
M1502 72 70 1196 vdd hvtpfet l=6e-08 w=8e-07 $X=7045 $Y=44777 $D=636
M1503 296 69 b_blb<12> vdd hvtpfet l=6e-08 w=3e-07 $X=7130 $Y=1094 $D=636
M1504 b_blb<12> 69 296 vdd hvtpfet l=6e-08 w=3e-07 $X=7130 $Y=1354 $D=636
M1505 b_blb_n<12> 69 297 vdd hvtpfet l=6e-08 w=3e-07 $X=7130 $Y=1864 $D=636
M1506 297 69 b_blb_n<12> vdd hvtpfet l=6e-08 w=3e-07 $X=7130 $Y=2124 $D=636
M1507 t_blb_n<12> 70 297 vdd hvtpfet l=6e-08 w=3e-07 $X=7130 $Y=48949 $D=636
M1508 297 70 t_blb_n<12> vdd hvtpfet l=6e-08 w=3e-07 $X=7130 $Y=49209 $D=636
M1509 296 70 t_blb<12> vdd hvtpfet l=6e-08 w=3e-07 $X=7130 $Y=49719 $D=636
M1510 t_blb<12> 70 296 vdd hvtpfet l=6e-08 w=3e-07 $X=7130 $Y=49979 $D=636
M1511 b_blb_n<12> 73 b_blb<12> vdd hvtpfet l=6e-08 w=8e-07 $X=7133 $Y=-170 $D=636
M1512 t_blb_n<12> 74 t_blb<12> vdd hvtpfet l=6e-08 w=8e-07 $X=7133 $Y=50503 $D=636
M1513 vdd vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=7295 $Y=35893 $D=636
M1514 vdd 73 b_blb_n<12> vdd hvtpfet l=6e-08 w=8e-07 $X=7393 $Y=-170 $D=636
M1515 vdd 74 t_blb_n<12> vdd hvtpfet l=6e-08 w=8e-07 $X=7393 $Y=50503 $D=636
M1516 b_blb_n<11> 77 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=7827 $Y=-170 $D=636
M1517 t_blb_n<11> 78 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=7827 $Y=50503 $D=636
M1518 vdd vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=7845 $Y=35893 $D=636
M1519 296 79 b_blb<11> vdd hvtpfet l=6e-08 w=3e-07 $X=7850 $Y=1094 $D=636
M1520 b_blb<11> 79 296 vdd hvtpfet l=6e-08 w=3e-07 $X=7850 $Y=1354 $D=636
M1521 b_blb_n<11> 79 297 vdd hvtpfet l=6e-08 w=3e-07 $X=7850 $Y=1864 $D=636
M1522 297 79 b_blb_n<11> vdd hvtpfet l=6e-08 w=3e-07 $X=7850 $Y=2124 $D=636
M1523 t_blb_n<11> 80 297 vdd hvtpfet l=6e-08 w=3e-07 $X=7850 $Y=48949 $D=636
M1524 297 80 t_blb_n<11> vdd hvtpfet l=6e-08 w=3e-07 $X=7850 $Y=49209 $D=636
M1525 296 80 t_blb<11> vdd hvtpfet l=6e-08 w=3e-07 $X=7850 $Y=49719 $D=636
M1526 t_blb<11> 80 296 vdd hvtpfet l=6e-08 w=3e-07 $X=7850 $Y=49979 $D=636
M1527 431 vdd vdd vdd hvtpfet l=6e-08 w=4e-07 $X=7895 $Y=21427 $D=636
M1528 432 vdd vdd vdd hvtpfet l=6e-08 w=4e-07 $X=7895 $Y=23694 $D=636
M1529 433 vdd vdd vdd hvtpfet l=6e-08 w=4e-07 $X=7895 $Y=24394 $D=636
M1530 434 vdd vdd vdd hvtpfet l=6e-08 w=4e-07 $X=7895 $Y=24904 $D=636
M1531 b_blb<11> 77 b_blb_n<11> vdd hvtpfet l=6e-08 w=8e-07 $X=8087 $Y=-170 $D=636
M1532 t_blb<11> 78 t_blb_n<11> vdd hvtpfet l=6e-08 w=8e-07 $X=8087 $Y=50503 $D=636
M1533 1201 79 81 vdd hvtpfet l=6e-08 w=8e-07 $X=8175 $Y=5556 $D=636
M1534 79 b_cb<3> vdd vdd hvtpfet l=6e-08 w=4e-07 $X=8175 $Y=10611 $D=636
M1535 77 79 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=8175 $Y=12911 $D=636
M1536 78 80 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=8175 $Y=37822 $D=636
M1537 80 t_cb<3> vdd vdd hvtpfet l=6e-08 w=4e-07 $X=8175 $Y=40122 $D=636
M1538 1202 80 82 vdd hvtpfet l=6e-08 w=8e-07 $X=8175 $Y=44777 $D=636
M1539 446 vdd vdd vdd hvtpfet l=6e-08 w=5e-07 $X=8180 $Y=18290 $D=636
M1540 vdd vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=8290 $Y=35893 $D=636
M1541 vdd vdd vdd vdd hvtpfet l=1e-07 w=2e-07 $X=8325 $Y=36723 $D=636
M1542 vdd 77 b_blb<11> vdd hvtpfet l=6e-08 w=8e-07 $X=8347 $Y=-170 $D=636
M1543 vdd 78 t_blb<11> vdd hvtpfet l=6e-08 w=8e-07 $X=8347 $Y=50503 $D=636
M1544 vdd 11 1201 vdd hvtpfet l=6e-08 w=8e-07 $X=8435 $Y=5556 $D=636
M1545 vdd b_mb<2> 79 vdd hvtpfet l=6e-08 w=4e-07 $X=8435 $Y=10611 $D=636
M1546 vdd 13 77 vdd hvtpfet l=6e-08 w=4e-07 $X=8435 $Y=12911 $D=636
M1547 vdd 14 78 vdd hvtpfet l=6e-08 w=4e-07 $X=8435 $Y=37822 $D=636
M1548 vdd t_mb<2> 80 vdd hvtpfet l=6e-08 w=4e-07 $X=8435 $Y=40122 $D=636
M1549 vdd 11 1202 vdd hvtpfet l=6e-08 w=8e-07 $X=8435 $Y=44777 $D=636
M1550 vdd vdd 446 vdd hvtpfet l=6e-08 w=5e-07 $X=8440 $Y=18290 $D=636
M1551 vdd vdd vdd vdd hvtpfet l=6e-08 w=6e-07 $X=8507 $Y=29008 $D=636
M1552 vdd vdd vdd vdd hvtpfet l=1e-07 w=2e-07 $X=8625 $Y=36723 $D=636
M1553 vdd vdd vdd vdd hvtpfet l=7e-08 w=3.2e-07 $X=8630 $Y=32628 $D=636
M1554 vdd vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=8630 $Y=35893 $D=636
M1555 1203 20 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=8695 $Y=5556 $D=636
M1556 87 b_ma<2> vdd vdd hvtpfet l=6e-08 w=4e-07 $X=8695 $Y=10611 $D=636
M1557 91 22 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=8695 $Y=12911 $D=636
M1558 92 23 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=8695 $Y=37822 $D=636
M1559 88 t_ma<2> vdd vdd hvtpfet l=6e-08 w=4e-07 $X=8695 $Y=40122 $D=636
M1560 1204 20 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=8695 $Y=44777 $D=636
M1561 446 vdd vdd vdd hvtpfet l=6e-08 w=5e-07 $X=8700 $Y=18290 $D=636
M1562 vdd vdd vdd vdd hvtpfet l=6e-08 w=6e-07 $X=8767 $Y=29008 $D=636
M1563 b_bla_n<11> 91 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=8783 $Y=-170 $D=636
M1564 t_bla_n<11> 92 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=8783 $Y=50503 $D=636
M1565 vdd vdd 445 vdd hvtpfet l=6e-08 w=6e-07 $X=8907 $Y=27488 $D=636
M1566 vdd vdd vdd vdd hvtpfet l=7e-08 w=3.2e-07 $X=8920 $Y=32628 $D=636
M1567 vdd vdd vdd vdd hvtpfet l=1e-07 w=2e-07 $X=8925 $Y=36723 $D=636
M1568 85 87 1203 vdd hvtpfet l=6e-08 w=8e-07 $X=8955 $Y=5556 $D=636
M1569 vdd b_ca<3> 87 vdd hvtpfet l=6e-08 w=4e-07 $X=8955 $Y=10611 $D=636
M1570 vdd 87 91 vdd hvtpfet l=6e-08 w=4e-07 $X=8955 $Y=12911 $D=636
M1571 vdd 88 92 vdd hvtpfet l=6e-08 w=4e-07 $X=8955 $Y=37822 $D=636
M1572 vdd t_ca<3> 88 vdd hvtpfet l=6e-08 w=4e-07 $X=8955 $Y=40122 $D=636
M1573 86 88 1204 vdd hvtpfet l=6e-08 w=8e-07 $X=8955 $Y=44777 $D=636
M1574 vdd vdd 446 vdd hvtpfet l=6e-08 w=5e-07 $X=8960 $Y=18290 $D=636
M1575 vdd vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=8970 $Y=35893 $D=636
M1576 325 87 b_bla<11> vdd hvtpfet l=6e-08 w=3e-07 $X=9040 $Y=1094 $D=636
M1577 b_bla<11> 87 325 vdd hvtpfet l=6e-08 w=3e-07 $X=9040 $Y=1354 $D=636
M1578 b_bla_n<11> 87 326 vdd hvtpfet l=6e-08 w=3e-07 $X=9040 $Y=1864 $D=636
M1579 326 87 b_bla_n<11> vdd hvtpfet l=6e-08 w=3e-07 $X=9040 $Y=2124 $D=636
M1580 t_bla_n<11> 88 326 vdd hvtpfet l=6e-08 w=3e-07 $X=9040 $Y=48949 $D=636
M1581 326 88 t_bla_n<11> vdd hvtpfet l=6e-08 w=3e-07 $X=9040 $Y=49209 $D=636
M1582 325 88 t_bla<11> vdd hvtpfet l=6e-08 w=3e-07 $X=9040 $Y=49719 $D=636
M1583 t_bla<11> 88 325 vdd hvtpfet l=6e-08 w=3e-07 $X=9040 $Y=49979 $D=636
M1584 b_bla<11> 91 b_bla_n<11> vdd hvtpfet l=6e-08 w=8e-07 $X=9043 $Y=-170 $D=636
M1585 t_bla<11> 92 t_bla_n<11> vdd hvtpfet l=6e-08 w=8e-07 $X=9043 $Y=50503 $D=636
M1586 vdd vdd vdd vdd hvtpfet l=1e-07 w=6e-07 $X=9200 $Y=32628 $D=636
M1587 vdd vdd vdd vdd hvtpfet l=1e-07 w=2e-07 $X=9225 $Y=36723 $D=636
M1588 vdd 91 b_bla<11> vdd hvtpfet l=6e-08 w=8e-07 $X=9303 $Y=-170 $D=636
M1589 vdd 92 t_bla<11> vdd hvtpfet l=6e-08 w=8e-07 $X=9303 $Y=50503 $D=636
M1590 vdd vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=9310 $Y=35893 $D=636
M1591 467 vdd vdd vdd hvtpfet l=6e-08 w=8e-07 $X=9427 $Y=27288 $D=636
M1592 461 vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=9445 $Y=15090 $D=636
M1593 462 vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=9445 $Y=16110 $D=636
M1594 477 vdd vdd vdd hvtpfet l=6e-08 w=6e-07 $X=9470 $Y=18290 $D=636
M1595 vdd vdd vdd vdd hvtpfet l=1e-07 w=6e-07 $X=9500 $Y=32628 $D=636
M1596 vdd vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=9650 $Y=35893 $D=636
M1597 vdd vdd vdd vdd hvtpfet l=6e-08 w=6e-07 $X=9677 $Y=29008 $D=636
M1598 vdd vdd 467 vdd hvtpfet l=6e-08 w=8e-07 $X=9687 $Y=27288 $D=636
M1599 vdd vdd 477 vdd hvtpfet l=6e-08 w=6e-07 $X=9730 $Y=18290 $D=636
M1600 b_bla<10> 95 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=9737 $Y=-170 $D=636
M1601 t_bla<10> 96 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=9737 $Y=50503 $D=636
M1602 325 93 b_bla<10> vdd hvtpfet l=6e-08 w=3e-07 $X=9760 $Y=1094 $D=636
M1603 b_bla<10> 93 325 vdd hvtpfet l=6e-08 w=3e-07 $X=9760 $Y=1354 $D=636
M1604 b_bla_n<10> 93 326 vdd hvtpfet l=6e-08 w=3e-07 $X=9760 $Y=1864 $D=636
M1605 326 93 b_bla_n<10> vdd hvtpfet l=6e-08 w=3e-07 $X=9760 $Y=2124 $D=636
M1606 t_bla_n<10> 94 326 vdd hvtpfet l=6e-08 w=3e-07 $X=9760 $Y=48949 $D=636
M1607 326 94 t_bla_n<10> vdd hvtpfet l=6e-08 w=3e-07 $X=9760 $Y=49209 $D=636
M1608 325 94 t_bla<10> vdd hvtpfet l=6e-08 w=3e-07 $X=9760 $Y=49719 $D=636
M1609 t_bla<10> 94 325 vdd hvtpfet l=6e-08 w=3e-07 $X=9760 $Y=49979 $D=636
M1610 vdd vdd vdd vdd hvtpfet l=1e-07 w=2e-07 $X=9775 $Y=36723 $D=636
M1611 vdd vdd 461 vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=9785 $Y=15090 $D=636
M1612 vdd vdd 462 vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=9785 $Y=16110 $D=636
M1613 vdd vdd vdd vdd hvtpfet l=1e-07 w=6e-07 $X=9800 $Y=32628 $D=636
M1614 vdd vdd vdd vdd hvtpfet l=6e-08 w=6e-07 $X=9937 $Y=29008 $D=636
M1615 467 vdd vdd vdd hvtpfet l=6e-08 w=8e-07 $X=9947 $Y=27288 $D=636
M1616 477 vdd vdd vdd hvtpfet l=6e-08 w=6e-07 $X=9990 $Y=18290 $D=636
M1617 vdd vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=9990 $Y=35893 $D=636
M1618 b_bla_n<10> 95 b_bla<10> vdd hvtpfet l=6e-08 w=8e-07 $X=9997 $Y=-170 $D=636
M1619 t_bla_n<10> 96 t_bla<10> vdd hvtpfet l=6e-08 w=8e-07 $X=9997 $Y=50503 $D=636
M1620 vdd vdd vdd vdd hvtpfet l=1e-07 w=2e-07 $X=10075 $Y=36723 $D=636
M1621 1209 93 97 vdd hvtpfet l=6e-08 w=8e-07 $X=10085 $Y=5556 $D=636
M1622 93 b_ca<2> vdd vdd hvtpfet l=6e-08 w=4e-07 $X=10085 $Y=10611 $D=636
M1623 95 93 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=10085 $Y=12911 $D=636
M1624 96 94 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=10085 $Y=37822 $D=636
M1625 94 t_ca<2> vdd vdd hvtpfet l=6e-08 w=4e-07 $X=10085 $Y=40122 $D=636
M1626 1210 94 98 vdd hvtpfet l=6e-08 w=8e-07 $X=10085 $Y=44777 $D=636
M1627 vdd vdd vdd vdd hvtpfet l=7e-08 w=3.2e-07 $X=10110 $Y=32628 $D=636
M1628 vdd vdd vdd vdd hvtpfet l=6e-08 w=6e-07 $X=10197 $Y=29008 $D=636
M1629 vdd vdd 467 vdd hvtpfet l=6e-08 w=8e-07 $X=10207 $Y=27288 $D=636
M1630 vdd vdd 477 vdd hvtpfet l=6e-08 w=6e-07 $X=10250 $Y=18290 $D=636
M1631 vdd 95 b_bla_n<10> vdd hvtpfet l=6e-08 w=8e-07 $X=10257 $Y=-170 $D=636
M1632 vdd 96 t_bla_n<10> vdd hvtpfet l=6e-08 w=8e-07 $X=10257 $Y=50503 $D=636
M1633 vdd vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=10330 $Y=35893 $D=636
M1634 vdd 20 1209 vdd hvtpfet l=6e-08 w=8e-07 $X=10345 $Y=5556 $D=636
M1635 vdd b_ma<2> 93 vdd hvtpfet l=6e-08 w=4e-07 $X=10345 $Y=10611 $D=636
M1636 vdd 22 95 vdd hvtpfet l=6e-08 w=4e-07 $X=10345 $Y=12911 $D=636
M1637 vdd 23 96 vdd hvtpfet l=6e-08 w=4e-07 $X=10345 $Y=37822 $D=636
M1638 vdd t_ma<2> 94 vdd hvtpfet l=6e-08 w=4e-07 $X=10345 $Y=40122 $D=636
M1639 vdd 20 1210 vdd hvtpfet l=6e-08 w=8e-07 $X=10345 $Y=44777 $D=636
M1640 475 vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=10375 $Y=15090 $D=636
M1641 476 vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=10375 $Y=16110 $D=636
M1642 vdd vdd vdd vdd hvtpfet l=1e-07 w=2e-07 $X=10375 $Y=36723 $D=636
M1643 vdd vdd vdd vdd hvtpfet l=7e-08 w=3.2e-07 $X=10400 $Y=32628 $D=636
M1644 vdd vdd vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=10446 $Y=19812 $D=636
M1645 vdd vdd vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=10446 $Y=20072 $D=636
M1646 vdd vdd vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=10446 $Y=21162 $D=636
M1647 vdd vdd vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=10446 $Y=21422 $D=636
M1648 vdd vdd vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=10446 $Y=21682 $D=636
M1649 vdd vdd vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=10446 $Y=21942 $D=636
M1650 vdd vdd vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=10446 $Y=22762 $D=636
M1651 vdd vdd vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=10446 $Y=23879 $D=636
M1652 vdd vdd vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=10446 $Y=24139 $D=636
M1653 vdd vdd vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=10446 $Y=24399 $D=636
M1654 vdd vdd vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=10446 $Y=24659 $D=636
M1655 vdd vdd vdd vdd hvtpfet l=6e-08 w=6e-07 $X=10457 $Y=29008 $D=636
M1656 477 vdd vdd vdd hvtpfet l=6e-08 w=6e-07 $X=10510 $Y=18290 $D=636
M1657 1211 11 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=10605 $Y=5556 $D=636
M1658 99 b_mb<2> vdd vdd hvtpfet l=6e-08 w=4e-07 $X=10605 $Y=10611 $D=636
M1659 103 13 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=10605 $Y=12911 $D=636
M1660 104 14 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=10605 $Y=37822 $D=636
M1661 100 t_mb<2> vdd vdd hvtpfet l=6e-08 w=4e-07 $X=10605 $Y=40122 $D=636
M1662 1212 11 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=10605 $Y=44777 $D=636
M1663 vdd vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=10670 $Y=35893 $D=636
M1664 vdd vdd vdd vdd hvtpfet l=1e-07 w=2e-07 $X=10675 $Y=36723 $D=636
M1665 b_blb<10> 103 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=10693 $Y=-170 $D=636
M1666 t_blb<10> 104 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=10693 $Y=50503 $D=636
M1667 vdd vdd 475 vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=10715 $Y=15090 $D=636
M1668 vdd vdd 476 vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=10715 $Y=16110 $D=636
M1669 484 vdd vdd vdd hvtpfet l=6e-08 w=6e-07 $X=10717 $Y=27488 $D=636
M1670 vdd vdd 477 vdd hvtpfet l=6e-08 w=6e-07 $X=10770 $Y=18290 $D=636
M1671 101 99 1211 vdd hvtpfet l=6e-08 w=8e-07 $X=10865 $Y=5556 $D=636
M1672 vdd b_cb<2> 99 vdd hvtpfet l=6e-08 w=4e-07 $X=10865 $Y=10611 $D=636
M1673 vdd 99 103 vdd hvtpfet l=6e-08 w=4e-07 $X=10865 $Y=12911 $D=636
M1674 vdd 100 104 vdd hvtpfet l=6e-08 w=4e-07 $X=10865 $Y=37822 $D=636
M1675 vdd t_cb<2> 100 vdd hvtpfet l=6e-08 w=4e-07 $X=10865 $Y=40122 $D=636
M1676 102 100 1212 vdd hvtpfet l=6e-08 w=8e-07 $X=10865 $Y=44777 $D=636
M1677 296 99 b_blb<10> vdd hvtpfet l=6e-08 w=3e-07 $X=10950 $Y=1094 $D=636
M1678 b_blb<10> 99 296 vdd hvtpfet l=6e-08 w=3e-07 $X=10950 $Y=1354 $D=636
M1679 b_blb_n<10> 99 297 vdd hvtpfet l=6e-08 w=3e-07 $X=10950 $Y=1864 $D=636
M1680 297 99 b_blb_n<10> vdd hvtpfet l=6e-08 w=3e-07 $X=10950 $Y=2124 $D=636
M1681 t_blb_n<10> 100 297 vdd hvtpfet l=6e-08 w=3e-07 $X=10950 $Y=48949 $D=636
M1682 297 100 t_blb_n<10> vdd hvtpfet l=6e-08 w=3e-07 $X=10950 $Y=49209 $D=636
M1683 296 100 t_blb<10> vdd hvtpfet l=6e-08 w=3e-07 $X=10950 $Y=49719 $D=636
M1684 t_blb<10> 100 296 vdd hvtpfet l=6e-08 w=3e-07 $X=10950 $Y=49979 $D=636
M1685 b_blb_n<10> 103 b_blb<10> vdd hvtpfet l=6e-08 w=8e-07 $X=10953 $Y=-170 $D=636
M1686 t_blb_n<10> 104 t_blb<10> vdd hvtpfet l=6e-08 w=8e-07 $X=10953 $Y=50503 $D=636
M1687 vdd vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=11115 $Y=35893 $D=636
M1688 vdd 103 b_blb_n<10> vdd hvtpfet l=6e-08 w=8e-07 $X=11213 $Y=-170 $D=636
M1689 vdd 104 t_blb_n<10> vdd hvtpfet l=6e-08 w=8e-07 $X=11213 $Y=50503 $D=636
M1690 b_blb_n<9> 105 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=11647 $Y=-170 $D=636
M1691 t_blb_n<9> 106 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=11647 $Y=50503 $D=636
M1692 vdd vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=11665 $Y=35893 $D=636
M1693 296 107 b_blb<9> vdd hvtpfet l=6e-08 w=3e-07 $X=11670 $Y=1094 $D=636
M1694 b_blb<9> 107 296 vdd hvtpfet l=6e-08 w=3e-07 $X=11670 $Y=1354 $D=636
M1695 b_blb_n<9> 107 297 vdd hvtpfet l=6e-08 w=3e-07 $X=11670 $Y=1864 $D=636
M1696 297 107 b_blb_n<9> vdd hvtpfet l=6e-08 w=3e-07 $X=11670 $Y=2124 $D=636
M1697 t_blb_n<9> 108 297 vdd hvtpfet l=6e-08 w=3e-07 $X=11670 $Y=48949 $D=636
M1698 297 108 t_blb_n<9> vdd hvtpfet l=6e-08 w=3e-07 $X=11670 $Y=49209 $D=636
M1699 296 108 t_blb<9> vdd hvtpfet l=6e-08 w=3e-07 $X=11670 $Y=49719 $D=636
M1700 t_blb<9> 108 296 vdd hvtpfet l=6e-08 w=3e-07 $X=11670 $Y=49979 $D=636
M1701 qa 125 vdd vdd hvtpfet l=6e-08 w=9e-07 $X=11758 $Y=19812 $D=636
M1702 qa 125 vdd vdd hvtpfet l=6e-08 w=9e-07 $X=11758 $Y=20072 $D=636
M1703 b_blb<9> 105 b_blb_n<9> vdd hvtpfet l=6e-08 w=8e-07 $X=11907 $Y=-170 $D=636
M1704 t_blb<9> 106 t_blb_n<9> vdd hvtpfet l=6e-08 w=8e-07 $X=11907 $Y=50503 $D=636
M1705 1217 107 112 vdd hvtpfet l=6e-08 w=8e-07 $X=11995 $Y=5556 $D=636
M1706 107 b_cb<1> vdd vdd hvtpfet l=6e-08 w=4e-07 $X=11995 $Y=10611 $D=636
M1707 105 107 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=11995 $Y=12911 $D=636
M1708 106 108 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=11995 $Y=37822 $D=636
M1709 108 t_cb<1> vdd vdd hvtpfet l=6e-08 w=4e-07 $X=11995 $Y=40122 $D=636
M1710 1218 108 113 vdd hvtpfet l=6e-08 w=8e-07 $X=11995 $Y=44777 $D=636
M1711 vdd vdd 498 vdd hvtpfet l=6e-08 w=6e-07 $X=12033 $Y=29008 $D=636
M1712 vdd bwena 122 vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=12065 $Y=15085 $D=636
M1713 vdd 114 134 vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=12065 $Y=16115 $D=636
M1714 516 vdd vdd vdd hvtpfet l=6e-08 w=6e-07 $X=12090 $Y=18290 $D=636
M1715 115 117 vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=12110 $Y=35893 $D=636
M1716 1219 134 vdd vdd hvtpfet l=6e-08 w=4.8e-07 $X=12113 $Y=21012 $D=636
M1717 1219 109 131 vdd hvtpfet l=6e-08 w=4.8e-07 $X=12113 $Y=21202 $D=636
M1718 119 131 vdd vdd hvtpfet l=6e-08 w=4.8e-07 $X=12113 $Y=22762 $D=636
M1719 1220 135 vdd vdd hvtpfet l=6e-08 w=4.8e-07 $X=12113 $Y=23729 $D=636
M1720 1220 109 132 vdd hvtpfet l=6e-08 w=4.8e-07 $X=12113 $Y=23919 $D=636
M1721 vdd 119 308 vdd hvtpfet l=6e-08 w=6e-07 $X=12143 $Y=27488 $D=636
M1722 115 118 325 vdd hvtpfet l=1e-07 w=2e-07 $X=12145 $Y=36723 $D=636
M1723 vdd 105 b_blb<9> vdd hvtpfet l=6e-08 w=8e-07 $X=12167 $Y=-170 $D=636
M1724 vdd 106 t_blb<9> vdd hvtpfet l=6e-08 w=8e-07 $X=12167 $Y=50503 $D=636
M1725 vdd 11 1217 vdd hvtpfet l=6e-08 w=8e-07 $X=12255 $Y=5556 $D=636
M1726 vdd b_mb<2> 107 vdd hvtpfet l=6e-08 w=4e-07 $X=12255 $Y=10611 $D=636
M1727 vdd 13 105 vdd hvtpfet l=6e-08 w=4e-07 $X=12255 $Y=12911 $D=636
M1728 vdd 14 106 vdd hvtpfet l=6e-08 w=4e-07 $X=12255 $Y=37822 $D=636
M1729 vdd t_mb<2> 108 vdd hvtpfet l=6e-08 w=4e-07 $X=12255 $Y=40122 $D=636
M1730 vdd 11 1218 vdd hvtpfet l=6e-08 w=8e-07 $X=12255 $Y=44777 $D=636
M1731 vdd 131 111 vdd hvtpfet l=6e-08 w=3.2e-07 $X=12273 $Y=21942 $D=636
M1732 vdd 132 110 vdd hvtpfet l=6e-08 w=3.2e-07 $X=12273 $Y=24659 $D=636
M1733 vdd vdd 516 vdd hvtpfet l=6e-08 w=6e-07 $X=12350 $Y=18290 $D=636
M1734 1221 111 131 vdd hvtpfet l=6e-08 w=2.1e-07 $X=12383 $Y=21477 $D=636
M1735 1221 129 vdd vdd hvtpfet l=6e-08 w=2.1e-07 $X=12383 $Y=21667 $D=636
M1736 1222 110 132 vdd hvtpfet l=6e-08 w=2.1e-07 $X=12383 $Y=24194 $D=636
M1737 1222 129 vdd vdd hvtpfet l=6e-08 w=2.1e-07 $X=12383 $Y=24384 $D=636
M1738 130 122 vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=12405 $Y=15085 $D=636
M1739 114 133 vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=12405 $Y=16115 $D=636
M1740 325 118 115 vdd hvtpfet l=1e-07 w=2e-07 $X=12445 $Y=36723 $D=636
M1741 ddqa_n 115 vdd vdd hvtpfet l=7e-08 w=3.2e-07 $X=12450 $Y=32628 $D=636
M1742 vdd 117 115 vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=12450 $Y=35893 $D=636
M1743 1223 20 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=12515 $Y=5556 $D=636
M1744 123 b_ma<2> vdd vdd hvtpfet l=6e-08 w=4e-07 $X=12515 $Y=10611 $D=636
M1745 127 22 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=12515 $Y=12911 $D=636
M1746 128 23 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=12515 $Y=37822 $D=636
M1747 124 t_ma<2> vdd vdd hvtpfet l=6e-08 w=4e-07 $X=12515 $Y=40122 $D=636
M1748 1224 20 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=12515 $Y=44777 $D=636
M1749 1225 118 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=12543 $Y=29008 $D=636
M1750 b_bla_n<9> 127 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=12603 $Y=-170 $D=636
M1751 t_bla_n<9> 128 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=12603 $Y=50503 $D=636
M1752 516 vdd vdd vdd hvtpfet l=6e-08 w=6e-07 $X=12610 $Y=18290 $D=636
M1753 20 126 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=12653 $Y=27288 $D=636
M1754 138 125 1225 vdd hvtpfet l=6e-08 w=6e-07 $X=12733 $Y=29008 $D=636
M1755 vdd 115 ddqa_n vdd hvtpfet l=7e-08 w=3.2e-07 $X=12740 $Y=32628 $D=636
M1756 115 118 325 vdd hvtpfet l=1e-07 w=2e-07 $X=12745 $Y=36723 $D=636
M1757 120 123 1223 vdd hvtpfet l=6e-08 w=8e-07 $X=12775 $Y=5556 $D=636
M1758 vdd b_ca<1> 123 vdd hvtpfet l=6e-08 w=4e-07 $X=12775 $Y=10611 $D=636
M1759 vdd 123 127 vdd hvtpfet l=6e-08 w=4e-07 $X=12775 $Y=12911 $D=636
M1760 vdd 124 128 vdd hvtpfet l=6e-08 w=4e-07 $X=12775 $Y=37822 $D=636
M1761 vdd t_ca<1> 124 vdd hvtpfet l=6e-08 w=4e-07 $X=12775 $Y=40122 $D=636
M1762 121 124 1224 vdd hvtpfet l=6e-08 w=8e-07 $X=12775 $Y=44777 $D=636
M1763 117 115 vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=12790 $Y=35893 $D=636
M1764 325 123 b_bla<9> vdd hvtpfet l=6e-08 w=3e-07 $X=12860 $Y=1094 $D=636
M1765 b_bla<9> 123 325 vdd hvtpfet l=6e-08 w=3e-07 $X=12860 $Y=1354 $D=636
M1766 b_bla_n<9> 123 326 vdd hvtpfet l=6e-08 w=3e-07 $X=12860 $Y=1864 $D=636
M1767 326 123 b_bla_n<9> vdd hvtpfet l=6e-08 w=3e-07 $X=12860 $Y=2124 $D=636
M1768 t_bla_n<9> 124 326 vdd hvtpfet l=6e-08 w=3e-07 $X=12860 $Y=48949 $D=636
M1769 326 124 t_bla_n<9> vdd hvtpfet l=6e-08 w=3e-07 $X=12860 $Y=49209 $D=636
M1770 325 124 t_bla<9> vdd hvtpfet l=6e-08 w=3e-07 $X=12860 $Y=49719 $D=636
M1771 t_bla<9> 124 325 vdd hvtpfet l=6e-08 w=3e-07 $X=12860 $Y=49979 $D=636
M1772 b_bla<9> 127 b_bla_n<9> vdd hvtpfet l=6e-08 w=8e-07 $X=12863 $Y=-170 $D=636
M1773 t_bla<9> 128 t_bla_n<9> vdd hvtpfet l=6e-08 w=8e-07 $X=12863 $Y=50503 $D=636
M1774 vdd vdd 516 vdd hvtpfet l=6e-08 w=6e-07 $X=12870 $Y=18290 $D=636
M1775 vdd 126 20 vdd hvtpfet l=6e-08 w=8e-07 $X=12913 $Y=27288 $D=636
M1776 1226 115 138 vdd hvtpfet l=6e-08 w=6e-07 $X=12993 $Y=29008 $D=636
M1777 vdd 130 141 vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=12995 $Y=15085 $D=636
M1778 vdd 136 133 vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=12995 $Y=16115 $D=636
M1779 115 sa_prea_n vdd vdd hvtpfet l=1e-07 w=6e-07 $X=13020 $Y=32628 $D=636
M1780 325 118 115 vdd hvtpfet l=1e-07 w=2e-07 $X=13045 $Y=36723 $D=636
M1781 vdd 127 b_bla<9> vdd hvtpfet l=6e-08 w=8e-07 $X=13123 $Y=-170 $D=636
M1782 vdd 128 t_bla<9> vdd hvtpfet l=6e-08 w=8e-07 $X=13123 $Y=50503 $D=636
M1783 516 vdd vdd vdd hvtpfet l=6e-08 w=6e-07 $X=13130 $Y=18290 $D=636
M1784 vdd 115 117 vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=13130 $Y=35893 $D=636
M1785 20 lwea vdd vdd hvtpfet l=6e-08 w=8e-07 $X=13173 $Y=27288 $D=636
M1786 vdd saea_n 1226 vdd hvtpfet l=6e-08 w=6e-07 $X=13183 $Y=29008 $D=636
M1787 117 sa_prea_n 115 vdd hvtpfet l=1e-07 w=6e-07 $X=13320 $Y=32628 $D=636
M1788 135 141 vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=13335 $Y=15085 $D=636
M1789 136 da vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=13335 $Y=16115 $D=636
M1790 vdd vdd 516 vdd hvtpfet l=6e-08 w=6e-07 $X=13390 $Y=18290 $D=636
M1791 vdd lwea 20 vdd hvtpfet l=6e-08 w=8e-07 $X=13433 $Y=27288 $D=636
M1792 115 117 vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=13470 $Y=35893 $D=636
M1793 b_bla<8> 145 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=13557 $Y=-170 $D=636
M1794 t_bla<8> 146 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=13557 $Y=50503 $D=636
M1795 325 143 b_bla<8> vdd hvtpfet l=6e-08 w=3e-07 $X=13580 $Y=1094 $D=636
M1796 b_bla<8> 143 325 vdd hvtpfet l=6e-08 w=3e-07 $X=13580 $Y=1354 $D=636
M1797 b_bla_n<8> 143 326 vdd hvtpfet l=6e-08 w=3e-07 $X=13580 $Y=1864 $D=636
M1798 326 143 b_bla_n<8> vdd hvtpfet l=6e-08 w=3e-07 $X=13580 $Y=2124 $D=636
M1799 t_bla_n<8> 144 326 vdd hvtpfet l=6e-08 w=3e-07 $X=13580 $Y=48949 $D=636
M1800 326 144 t_bla_n<8> vdd hvtpfet l=6e-08 w=3e-07 $X=13580 $Y=49209 $D=636
M1801 325 144 t_bla<8> vdd hvtpfet l=6e-08 w=3e-07 $X=13580 $Y=49719 $D=636
M1802 t_bla<8> 144 325 vdd hvtpfet l=6e-08 w=3e-07 $X=13580 $Y=49979 $D=636
M1803 117 118 326 vdd hvtpfet l=1e-07 w=2e-07 $X=13595 $Y=36723 $D=636
M1804 vdd sa_prea_n 117 vdd hvtpfet l=1e-07 w=6e-07 $X=13620 $Y=32628 $D=636
M1805 vdd 117 115 vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=13810 $Y=35893 $D=636
M1806 b_bla_n<8> 145 b_bla<8> vdd hvtpfet l=6e-08 w=8e-07 $X=13817 $Y=-170 $D=636
M1807 t_bla_n<8> 146 t_bla<8> vdd hvtpfet l=6e-08 w=8e-07 $X=13817 $Y=50503 $D=636
M1808 326 118 117 vdd hvtpfet l=1e-07 w=2e-07 $X=13895 $Y=36723 $D=636
M1809 22 b_tm_prea_n vdd vdd hvtpfet l=6e-08 w=5e-07 $X=13900 $Y=18290 $D=636
M1810 1231 143 148 vdd hvtpfet l=6e-08 w=8e-07 $X=13905 $Y=5556 $D=636
M1811 143 b_ca<0> vdd vdd hvtpfet l=6e-08 w=4e-07 $X=13905 $Y=10611 $D=636
M1812 145 143 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=13905 $Y=12911 $D=636
M1813 146 144 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=13905 $Y=37822 $D=636
M1814 144 t_ca<0> vdd vdd hvtpfet l=6e-08 w=4e-07 $X=13905 $Y=40122 $D=636
M1815 1232 144 149 vdd hvtpfet l=6e-08 w=8e-07 $X=13905 $Y=44777 $D=636
M1816 ddqa 117 vdd vdd hvtpfet l=7e-08 w=3.2e-07 $X=13930 $Y=32628 $D=636
M1817 328 131 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=13953 $Y=27488 $D=636
M1818 vdd 145 b_bla_n<8> vdd hvtpfet l=6e-08 w=8e-07 $X=14077 $Y=-170 $D=636
M1819 vdd 146 t_bla_n<8> vdd hvtpfet l=6e-08 w=8e-07 $X=14077 $Y=50503 $D=636
M1820 vdd 138 125 vdd hvtpfet l=6e-08 w=6e-07 $X=14093 $Y=29008 $D=636
M1821 117 115 vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=14150 $Y=35893 $D=636
M1822 vdd b_tm_prea_n 22 vdd hvtpfet l=6e-08 w=5e-07 $X=14160 $Y=18290 $D=636
M1823 vdd 20 1231 vdd hvtpfet l=6e-08 w=8e-07 $X=14165 $Y=5556 $D=636
M1824 vdd b_ma<2> 143 vdd hvtpfet l=6e-08 w=4e-07 $X=14165 $Y=10611 $D=636
M1825 vdd 22 145 vdd hvtpfet l=6e-08 w=4e-07 $X=14165 $Y=12911 $D=636
M1826 vdd 23 146 vdd hvtpfet l=6e-08 w=4e-07 $X=14165 $Y=37822 $D=636
M1827 vdd t_ma<2> 144 vdd hvtpfet l=6e-08 w=4e-07 $X=14165 $Y=40122 $D=636
M1828 vdd 20 1232 vdd hvtpfet l=6e-08 w=8e-07 $X=14165 $Y=44777 $D=636
M1829 117 118 326 vdd hvtpfet l=1e-07 w=2e-07 $X=14195 $Y=36723 $D=636
M1830 vdd 117 ddqa vdd hvtpfet l=7e-08 w=3.2e-07 $X=14220 $Y=32628 $D=636
M1831 118 saea_n vdd vdd hvtpfet l=6e-08 w=6e-07 $X=14353 $Y=29008 $D=636
M1832 23 t_tm_prea_n vdd vdd hvtpfet l=6e-08 w=5e-07 $X=14420 $Y=18290 $D=636
M1833 1233 11 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=14425 $Y=5556 $D=636
M1834 153 b_mb<2> vdd vdd hvtpfet l=6e-08 w=4e-07 $X=14425 $Y=10611 $D=636
M1835 157 13 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=14425 $Y=12911 $D=636
M1836 158 14 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=14425 $Y=37822 $D=636
M1837 154 t_mb<2> vdd vdd hvtpfet l=6e-08 w=4e-07 $X=14425 $Y=40122 $D=636
M1838 1234 11 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=14425 $Y=44777 $D=636
M1839 vdd 115 117 vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=14490 $Y=35893 $D=636
M1840 326 118 117 vdd hvtpfet l=1e-07 w=2e-07 $X=14495 $Y=36723 $D=636
M1841 b_blb<8> 157 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=14513 $Y=-170 $D=636
M1842 t_blb<8> 158 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=14513 $Y=50503 $D=636
M1843 129 clk_dqa vdd vdd hvtpfet l=6e-08 w=4e-07 $X=14625 $Y=21427 $D=636
M1844 109 clk_dqa_n vdd vdd hvtpfet l=6e-08 w=4e-07 $X=14625 $Y=23694 $D=636
M1845 152 132 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=14625 $Y=24394 $D=636
M1846 126 152 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=14625 $Y=24904 $D=636
M1847 vdd t_tm_prea_n 23 vdd hvtpfet l=6e-08 w=5e-07 $X=14680 $Y=18290 $D=636
M1848 155 153 1233 vdd hvtpfet l=6e-08 w=8e-07 $X=14685 $Y=5556 $D=636
M1849 vdd b_cb<0> 153 vdd hvtpfet l=6e-08 w=4e-07 $X=14685 $Y=10611 $D=636
M1850 vdd 153 157 vdd hvtpfet l=6e-08 w=4e-07 $X=14685 $Y=12911 $D=636
M1851 vdd 154 158 vdd hvtpfet l=6e-08 w=4e-07 $X=14685 $Y=37822 $D=636
M1852 vdd t_cb<0> 154 vdd hvtpfet l=6e-08 w=4e-07 $X=14685 $Y=40122 $D=636
M1853 156 154 1234 vdd hvtpfet l=6e-08 w=8e-07 $X=14685 $Y=44777 $D=636
M1854 296 153 b_blb<8> vdd hvtpfet l=6e-08 w=3e-07 $X=14770 $Y=1094 $D=636
M1855 b_blb<8> 153 296 vdd hvtpfet l=6e-08 w=3e-07 $X=14770 $Y=1354 $D=636
M1856 b_blb_n<8> 153 297 vdd hvtpfet l=6e-08 w=3e-07 $X=14770 $Y=1864 $D=636
M1857 297 153 b_blb_n<8> vdd hvtpfet l=6e-08 w=3e-07 $X=14770 $Y=2124 $D=636
M1858 t_blb_n<8> 154 297 vdd hvtpfet l=6e-08 w=3e-07 $X=14770 $Y=48949 $D=636
M1859 297 154 t_blb_n<8> vdd hvtpfet l=6e-08 w=3e-07 $X=14770 $Y=49209 $D=636
M1860 296 154 t_blb<8> vdd hvtpfet l=6e-08 w=3e-07 $X=14770 $Y=49719 $D=636
M1861 t_blb<8> 154 296 vdd hvtpfet l=6e-08 w=3e-07 $X=14770 $Y=49979 $D=636
M1862 b_blb_n<8> 157 b_blb<8> vdd hvtpfet l=6e-08 w=8e-07 $X=14773 $Y=-170 $D=636
M1863 t_blb_n<8> 158 t_blb<8> vdd hvtpfet l=6e-08 w=8e-07 $X=14773 $Y=50503 $D=636
M1864 544 117 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=14863 $Y=29008 $D=636
M1865 vdd vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=14935 $Y=35893 $D=636
M1866 vdd 157 b_blb_n<8> vdd hvtpfet l=6e-08 w=8e-07 $X=15033 $Y=-170 $D=636
M1867 vdd 158 t_blb_n<8> vdd hvtpfet l=6e-08 w=8e-07 $X=15033 $Y=50503 $D=636
M1868 b_blb_n<7> 161 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=15467 $Y=-170 $D=636
M1869 t_blb_n<7> 162 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=15467 $Y=50503 $D=636
M1870 vdd vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=15485 $Y=35893 $D=636
M1871 296 163 b_blb<7> vdd hvtpfet l=6e-08 w=3e-07 $X=15490 $Y=1094 $D=636
M1872 b_blb<7> 163 296 vdd hvtpfet l=6e-08 w=3e-07 $X=15490 $Y=1354 $D=636
M1873 b_blb_n<7> 163 297 vdd hvtpfet l=6e-08 w=3e-07 $X=15490 $Y=1864 $D=636
M1874 297 163 b_blb_n<7> vdd hvtpfet l=6e-08 w=3e-07 $X=15490 $Y=2124 $D=636
M1875 t_blb_n<7> 164 297 vdd hvtpfet l=6e-08 w=3e-07 $X=15490 $Y=48949 $D=636
M1876 297 164 t_blb_n<7> vdd hvtpfet l=6e-08 w=3e-07 $X=15490 $Y=49209 $D=636
M1877 296 164 t_blb<7> vdd hvtpfet l=6e-08 w=3e-07 $X=15490 $Y=49719 $D=636
M1878 t_blb<7> 164 296 vdd hvtpfet l=6e-08 w=3e-07 $X=15490 $Y=49979 $D=636
M1879 192 clk_dqb vdd vdd hvtpfet l=6e-08 w=4e-07 $X=15535 $Y=21427 $D=636
M1880 190 clk_dqb_n vdd vdd hvtpfet l=6e-08 w=4e-07 $X=15535 $Y=23694 $D=636
M1881 174 173 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=15535 $Y=24394 $D=636
M1882 200 174 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=15535 $Y=24904 $D=636
M1883 vdd 160 551 vdd hvtpfet l=6e-08 w=6e-07 $X=15637 $Y=29008 $D=636
M1884 b_blb<7> 161 b_blb_n<7> vdd hvtpfet l=6e-08 w=8e-07 $X=15727 $Y=-170 $D=636
M1885 t_blb<7> 162 t_blb_n<7> vdd hvtpfet l=6e-08 w=8e-07 $X=15727 $Y=50503 $D=636
M1886 1239 163 166 vdd hvtpfet l=6e-08 w=8e-07 $X=15815 $Y=5556 $D=636
M1887 163 b_cb<3> vdd vdd hvtpfet l=6e-08 w=4e-07 $X=15815 $Y=10611 $D=636
M1888 161 163 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=15815 $Y=12911 $D=636
M1889 162 164 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=15815 $Y=37822 $D=636
M1890 164 t_cb<3> vdd vdd hvtpfet l=6e-08 w=4e-07 $X=15815 $Y=40122 $D=636
M1891 1240 164 167 vdd hvtpfet l=6e-08 w=8e-07 $X=15815 $Y=44777 $D=636
M1892 14 t_tm_preb_n vdd vdd hvtpfet l=6e-08 w=5e-07 $X=15820 $Y=18290 $D=636
M1893 160 168 vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=15930 $Y=35893 $D=636
M1894 160 169 297 vdd hvtpfet l=1e-07 w=2e-07 $X=15965 $Y=36723 $D=636
M1895 vdd 161 b_blb<7> vdd hvtpfet l=6e-08 w=8e-07 $X=15987 $Y=-170 $D=636
M1896 vdd 162 t_blb<7> vdd hvtpfet l=6e-08 w=8e-07 $X=15987 $Y=50503 $D=636
M1897 vdd 11 1239 vdd hvtpfet l=6e-08 w=8e-07 $X=16075 $Y=5556 $D=636
M1898 vdd b_mb<1> 163 vdd hvtpfet l=6e-08 w=4e-07 $X=16075 $Y=10611 $D=636
M1899 vdd 13 161 vdd hvtpfet l=6e-08 w=4e-07 $X=16075 $Y=12911 $D=636
M1900 vdd 14 162 vdd hvtpfet l=6e-08 w=4e-07 $X=16075 $Y=37822 $D=636
M1901 vdd t_mb<1> 164 vdd hvtpfet l=6e-08 w=4e-07 $X=16075 $Y=40122 $D=636
M1902 vdd 11 1240 vdd hvtpfet l=6e-08 w=8e-07 $X=16075 $Y=44777 $D=636
M1903 vdd t_tm_preb_n 14 vdd hvtpfet l=6e-08 w=5e-07 $X=16080 $Y=18290 $D=636
M1904 vdd saeb_n 169 vdd hvtpfet l=6e-08 w=6e-07 $X=16147 $Y=29008 $D=636
M1905 297 169 160 vdd hvtpfet l=1e-07 w=2e-07 $X=16265 $Y=36723 $D=636
M1906 ddqb 160 vdd vdd hvtpfet l=7e-08 w=3.2e-07 $X=16270 $Y=32628 $D=636
M1907 vdd 168 160 vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=16270 $Y=35893 $D=636
M1908 1241 20 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=16335 $Y=5556 $D=636
M1909 179 b_ma<1> vdd vdd hvtpfet l=6e-08 w=4e-07 $X=16335 $Y=10611 $D=636
M1910 184 22 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=16335 $Y=12911 $D=636
M1911 185 23 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=16335 $Y=37822 $D=636
M1912 180 t_ma<1> vdd vdd hvtpfet l=6e-08 w=4e-07 $X=16335 $Y=40122 $D=636
M1913 1242 20 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=16335 $Y=44777 $D=636
M1914 13 b_tm_preb_n vdd vdd hvtpfet l=6e-08 w=5e-07 $X=16340 $Y=18290 $D=636
M1915 189 194 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=16407 $Y=29008 $D=636
M1916 b_bla_n<7> 184 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=16423 $Y=-170 $D=636
M1917 t_bla_n<7> 185 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=16423 $Y=50503 $D=636
M1918 vdd 178 299 vdd hvtpfet l=6e-08 w=6e-07 $X=16547 $Y=27488 $D=636
M1919 vdd 160 ddqb vdd hvtpfet l=7e-08 w=3.2e-07 $X=16560 $Y=32628 $D=636
M1920 160 169 297 vdd hvtpfet l=1e-07 w=2e-07 $X=16565 $Y=36723 $D=636
M1921 176 179 1241 vdd hvtpfet l=6e-08 w=8e-07 $X=16595 $Y=5556 $D=636
M1922 vdd b_ca<3> 179 vdd hvtpfet l=6e-08 w=4e-07 $X=16595 $Y=10611 $D=636
M1923 vdd 179 184 vdd hvtpfet l=6e-08 w=4e-07 $X=16595 $Y=12911 $D=636
M1924 vdd 180 185 vdd hvtpfet l=6e-08 w=4e-07 $X=16595 $Y=37822 $D=636
M1925 vdd t_ca<3> 180 vdd hvtpfet l=6e-08 w=4e-07 $X=16595 $Y=40122 $D=636
M1926 177 180 1242 vdd hvtpfet l=6e-08 w=8e-07 $X=16595 $Y=44777 $D=636
M1927 vdd b_tm_preb_n 13 vdd hvtpfet l=6e-08 w=5e-07 $X=16600 $Y=18290 $D=636
M1928 168 160 vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=16610 $Y=35893 $D=636
M1929 325 179 b_bla<7> vdd hvtpfet l=6e-08 w=3e-07 $X=16680 $Y=1094 $D=636
M1930 b_bla<7> 179 325 vdd hvtpfet l=6e-08 w=3e-07 $X=16680 $Y=1354 $D=636
M1931 b_bla_n<7> 179 326 vdd hvtpfet l=6e-08 w=3e-07 $X=16680 $Y=1864 $D=636
M1932 326 179 b_bla_n<7> vdd hvtpfet l=6e-08 w=3e-07 $X=16680 $Y=2124 $D=636
M1933 t_bla_n<7> 180 326 vdd hvtpfet l=6e-08 w=3e-07 $X=16680 $Y=48949 $D=636
M1934 326 180 t_bla_n<7> vdd hvtpfet l=6e-08 w=3e-07 $X=16680 $Y=49209 $D=636
M1935 325 180 t_bla<7> vdd hvtpfet l=6e-08 w=3e-07 $X=16680 $Y=49719 $D=636
M1936 t_bla<7> 180 325 vdd hvtpfet l=6e-08 w=3e-07 $X=16680 $Y=49979 $D=636
M1937 b_bla<7> 184 b_bla_n<7> vdd hvtpfet l=6e-08 w=8e-07 $X=16683 $Y=-170 $D=636
M1938 t_bla<7> 185 t_bla_n<7> vdd hvtpfet l=6e-08 w=8e-07 $X=16683 $Y=50503 $D=636
M1939 160 sa_preb_n vdd vdd hvtpfet l=1e-07 w=6e-07 $X=16840 $Y=32628 $D=636
M1940 297 169 160 vdd hvtpfet l=1e-07 w=2e-07 $X=16865 $Y=36723 $D=636
M1941 vdd 184 b_bla<7> vdd hvtpfet l=6e-08 w=8e-07 $X=16943 $Y=-170 $D=636
M1942 vdd 185 t_bla<7> vdd hvtpfet l=6e-08 w=8e-07 $X=16943 $Y=50503 $D=636
M1943 vdd 160 168 vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=16950 $Y=35893 $D=636
M1944 11 lweb vdd vdd hvtpfet l=6e-08 w=8e-07 $X=17067 $Y=27288 $D=636
M1945 vdd 191 202 vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=17085 $Y=15085 $D=636
M1946 vdd db 195 vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=17085 $Y=16115 $D=636
M1947 587 vdd vdd vdd hvtpfet l=6e-08 w=6e-07 $X=17110 $Y=18290 $D=636
M1948 168 sa_preb_n 160 vdd hvtpfet l=1e-07 w=6e-07 $X=17140 $Y=32628 $D=636
M1949 160 168 vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=17290 $Y=35893 $D=636
M1950 1243 saeb_n vdd vdd hvtpfet l=6e-08 w=6e-07 $X=17317 $Y=29008 $D=636
M1951 vdd lweb 11 vdd hvtpfet l=6e-08 w=8e-07 $X=17327 $Y=27288 $D=636
M1952 vdd vdd 587 vdd hvtpfet l=6e-08 w=6e-07 $X=17370 $Y=18290 $D=636
M1953 b_bla<6> 198 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=17377 $Y=-170 $D=636
M1954 t_bla<6> 199 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=17377 $Y=50503 $D=636
M1955 325 196 b_bla<6> vdd hvtpfet l=6e-08 w=3e-07 $X=17400 $Y=1094 $D=636
M1956 b_bla<6> 196 325 vdd hvtpfet l=6e-08 w=3e-07 $X=17400 $Y=1354 $D=636
M1957 b_bla_n<6> 196 326 vdd hvtpfet l=6e-08 w=3e-07 $X=17400 $Y=1864 $D=636
M1958 326 196 b_bla_n<6> vdd hvtpfet l=6e-08 w=3e-07 $X=17400 $Y=2124 $D=636
M1959 t_bla_n<6> 197 326 vdd hvtpfet l=6e-08 w=3e-07 $X=17400 $Y=48949 $D=636
M1960 326 197 t_bla_n<6> vdd hvtpfet l=6e-08 w=3e-07 $X=17400 $Y=49209 $D=636
M1961 325 197 t_bla<6> vdd hvtpfet l=6e-08 w=3e-07 $X=17400 $Y=49719 $D=636
M1962 t_bla<6> 197 325 vdd hvtpfet l=6e-08 w=3e-07 $X=17400 $Y=49979 $D=636
M1963 168 169 296 vdd hvtpfet l=1e-07 w=2e-07 $X=17415 $Y=36723 $D=636
M1964 191 204 vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=17425 $Y=15085 $D=636
M1965 203 195 vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=17425 $Y=16115 $D=636
M1966 vdd sa_preb_n 168 vdd hvtpfet l=1e-07 w=6e-07 $X=17440 $Y=32628 $D=636
M1967 194 168 1243 vdd hvtpfet l=6e-08 w=6e-07 $X=17507 $Y=29008 $D=636
M1968 11 200 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=17587 $Y=27288 $D=636
M1969 587 vdd vdd vdd hvtpfet l=6e-08 w=6e-07 $X=17630 $Y=18290 $D=636
M1970 vdd 168 160 vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=17630 $Y=35893 $D=636
M1971 b_bla_n<6> 198 b_bla<6> vdd hvtpfet l=6e-08 w=8e-07 $X=17637 $Y=-170 $D=636
M1972 t_bla_n<6> 199 t_bla<6> vdd hvtpfet l=6e-08 w=8e-07 $X=17637 $Y=50503 $D=636
M1973 296 169 168 vdd hvtpfet l=1e-07 w=2e-07 $X=17715 $Y=36723 $D=636
M1974 1248 196 205 vdd hvtpfet l=6e-08 w=8e-07 $X=17725 $Y=5556 $D=636
M1975 196 b_ca<2> vdd vdd hvtpfet l=6e-08 w=4e-07 $X=17725 $Y=10611 $D=636
M1976 198 196 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=17725 $Y=12911 $D=636
M1977 199 197 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=17725 $Y=37822 $D=636
M1978 197 t_ca<2> vdd vdd hvtpfet l=6e-08 w=4e-07 $X=17725 $Y=40122 $D=636
M1979 1249 197 206 vdd hvtpfet l=6e-08 w=8e-07 $X=17725 $Y=44777 $D=636
M1980 ddqb_n 168 vdd vdd hvtpfet l=7e-08 w=3.2e-07 $X=17750 $Y=32628 $D=636
M1981 1250 189 194 vdd hvtpfet l=6e-08 w=6e-07 $X=17767 $Y=29008 $D=636
M1982 vdd 200 11 vdd hvtpfet l=6e-08 w=8e-07 $X=17847 $Y=27288 $D=636
M1983 vdd vdd 587 vdd hvtpfet l=6e-08 w=6e-07 $X=17890 $Y=18290 $D=636
M1984 vdd 198 b_bla_n<6> vdd hvtpfet l=6e-08 w=8e-07 $X=17897 $Y=-170 $D=636
M1985 vdd 199 t_bla_n<6> vdd hvtpfet l=6e-08 w=8e-07 $X=17897 $Y=50503 $D=636
M1986 qb 189 vdd vdd hvtpfet l=6e-08 w=9e-07 $X=17902 $Y=19812 $D=636
M1987 qb 189 vdd vdd hvtpfet l=6e-08 w=9e-07 $X=17902 $Y=20072 $D=636
M1988 vdd 169 1250 vdd hvtpfet l=6e-08 w=6e-07 $X=17957 $Y=29008 $D=636
M1989 1251 201 vdd vdd hvtpfet l=6e-08 w=4.8e-07 $X=17967 $Y=21012 $D=636
M1990 1251 190 178 vdd hvtpfet l=6e-08 w=4.8e-07 $X=17967 $Y=21202 $D=636
M1991 1252 217 178 vdd hvtpfet l=6e-08 w=2.1e-07 $X=17967 $Y=21477 $D=636
M1992 1252 192 vdd vdd hvtpfet l=6e-08 w=2.1e-07 $X=17967 $Y=21667 $D=636
M1993 vdd 178 217 vdd hvtpfet l=6e-08 w=3.2e-07 $X=17967 $Y=21942 $D=636
M1994 208 178 vdd vdd hvtpfet l=6e-08 w=4.8e-07 $X=17967 $Y=22762 $D=636
M1995 1253 202 vdd vdd hvtpfet l=6e-08 w=4.8e-07 $X=17967 $Y=23729 $D=636
M1996 1253 190 173 vdd hvtpfet l=6e-08 w=4.8e-07 $X=17967 $Y=23919 $D=636
M1997 1254 218 173 vdd hvtpfet l=6e-08 w=2.1e-07 $X=17967 $Y=24194 $D=636
M1998 1254 192 vdd vdd hvtpfet l=6e-08 w=2.1e-07 $X=17967 $Y=24384 $D=636
M1999 vdd 173 218 vdd hvtpfet l=6e-08 w=3.2e-07 $X=17967 $Y=24659 $D=636
M2000 168 160 vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=17970 $Y=35893 $D=636
M2001 vdd 20 1248 vdd hvtpfet l=6e-08 w=8e-07 $X=17985 $Y=5556 $D=636
M2002 vdd b_ma<1> 196 vdd hvtpfet l=6e-08 w=4e-07 $X=17985 $Y=10611 $D=636
M2003 vdd 22 198 vdd hvtpfet l=6e-08 w=4e-07 $X=17985 $Y=12911 $D=636
M2004 vdd 23 199 vdd hvtpfet l=6e-08 w=4e-07 $X=17985 $Y=37822 $D=636
M2005 vdd t_ma<1> 197 vdd hvtpfet l=6e-08 w=4e-07 $X=17985 $Y=40122 $D=636
M2006 vdd 20 1249 vdd hvtpfet l=6e-08 w=8e-07 $X=17985 $Y=44777 $D=636
M2007 vdd 207 204 vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=18015 $Y=15085 $D=636
M2008 vdd 203 216 vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=18015 $Y=16115 $D=636
M2009 168 169 296 vdd hvtpfet l=1e-07 w=2e-07 $X=18015 $Y=36723 $D=636
M2010 vdd 168 ddqb_n vdd hvtpfet l=7e-08 w=3.2e-07 $X=18040 $Y=32628 $D=636
M2011 587 vdd vdd vdd hvtpfet l=6e-08 w=6e-07 $X=18150 $Y=18290 $D=636
M2012 1255 11 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=18245 $Y=5556 $D=636
M2013 209 b_mb<1> vdd vdd hvtpfet l=6e-08 w=4e-07 $X=18245 $Y=10611 $D=636
M2014 214 13 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=18245 $Y=12911 $D=636
M2015 215 14 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=18245 $Y=37822 $D=636
M2016 210 t_mb<1> vdd vdd hvtpfet l=6e-08 w=4e-07 $X=18245 $Y=40122 $D=636
M2017 1256 11 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=18245 $Y=44777 $D=636
M2018 vdd 160 168 vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=18310 $Y=35893 $D=636
M2019 296 169 168 vdd hvtpfet l=1e-07 w=2e-07 $X=18315 $Y=36723 $D=636
M2020 b_blb<6> 214 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=18333 $Y=-170 $D=636
M2021 t_blb<6> 215 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=18333 $Y=50503 $D=636
M2022 207 bwenb vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=18355 $Y=15085 $D=636
M2023 201 216 vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=18355 $Y=16115 $D=636
M2024 317 208 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=18357 $Y=27488 $D=636
M2025 vdd vdd 587 vdd hvtpfet l=6e-08 w=6e-07 $X=18410 $Y=18290 $D=636
M2026 598 vdd vdd vdd hvtpfet l=6e-08 w=6e-07 $X=18467 $Y=29008 $D=636
M2027 211 209 1255 vdd hvtpfet l=6e-08 w=8e-07 $X=18505 $Y=5556 $D=636
M2028 vdd b_cb<2> 209 vdd hvtpfet l=6e-08 w=4e-07 $X=18505 $Y=10611 $D=636
M2029 vdd 209 214 vdd hvtpfet l=6e-08 w=4e-07 $X=18505 $Y=12911 $D=636
M2030 vdd 210 215 vdd hvtpfet l=6e-08 w=4e-07 $X=18505 $Y=37822 $D=636
M2031 vdd t_cb<2> 210 vdd hvtpfet l=6e-08 w=4e-07 $X=18505 $Y=40122 $D=636
M2032 212 210 1256 vdd hvtpfet l=6e-08 w=8e-07 $X=18505 $Y=44777 $D=636
M2033 296 209 b_blb<6> vdd hvtpfet l=6e-08 w=3e-07 $X=18590 $Y=1094 $D=636
M2034 b_blb<6> 209 296 vdd hvtpfet l=6e-08 w=3e-07 $X=18590 $Y=1354 $D=636
M2035 b_blb_n<6> 209 297 vdd hvtpfet l=6e-08 w=3e-07 $X=18590 $Y=1864 $D=636
M2036 297 209 b_blb_n<6> vdd hvtpfet l=6e-08 w=3e-07 $X=18590 $Y=2124 $D=636
M2037 t_blb_n<6> 210 297 vdd hvtpfet l=6e-08 w=3e-07 $X=18590 $Y=48949 $D=636
M2038 297 210 t_blb_n<6> vdd hvtpfet l=6e-08 w=3e-07 $X=18590 $Y=49209 $D=636
M2039 296 210 t_blb<6> vdd hvtpfet l=6e-08 w=3e-07 $X=18590 $Y=49719 $D=636
M2040 t_blb<6> 210 296 vdd hvtpfet l=6e-08 w=3e-07 $X=18590 $Y=49979 $D=636
M2041 b_blb_n<6> 214 b_blb<6> vdd hvtpfet l=6e-08 w=8e-07 $X=18593 $Y=-170 $D=636
M2042 t_blb_n<6> 215 t_blb<6> vdd hvtpfet l=6e-08 w=8e-07 $X=18593 $Y=50503 $D=636
M2043 vdd vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=18755 $Y=35893 $D=636
M2044 vdd 214 b_blb_n<6> vdd hvtpfet l=6e-08 w=8e-07 $X=18853 $Y=-170 $D=636
M2045 vdd 215 t_blb_n<6> vdd hvtpfet l=6e-08 w=8e-07 $X=18853 $Y=50503 $D=636
M2046 b_blb_n<5> 219 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=19287 $Y=-170 $D=636
M2047 t_blb_n<5> 220 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=19287 $Y=50503 $D=636
M2048 vdd vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=19305 $Y=35893 $D=636
M2049 296 221 b_blb<5> vdd hvtpfet l=6e-08 w=3e-07 $X=19310 $Y=1094 $D=636
M2050 b_blb<5> 221 296 vdd hvtpfet l=6e-08 w=3e-07 $X=19310 $Y=1354 $D=636
M2051 b_blb_n<5> 221 297 vdd hvtpfet l=6e-08 w=3e-07 $X=19310 $Y=1864 $D=636
M2052 297 221 b_blb_n<5> vdd hvtpfet l=6e-08 w=3e-07 $X=19310 $Y=2124 $D=636
M2053 t_blb_n<5> 222 297 vdd hvtpfet l=6e-08 w=3e-07 $X=19310 $Y=48949 $D=636
M2054 297 222 t_blb_n<5> vdd hvtpfet l=6e-08 w=3e-07 $X=19310 $Y=49209 $D=636
M2055 296 222 t_blb<5> vdd hvtpfet l=6e-08 w=3e-07 $X=19310 $Y=49719 $D=636
M2056 t_blb<5> 222 296 vdd hvtpfet l=6e-08 w=3e-07 $X=19310 $Y=49979 $D=636
M2057 b_blb<5> 219 b_blb_n<5> vdd hvtpfet l=6e-08 w=8e-07 $X=19547 $Y=-170 $D=636
M2058 t_blb<5> 220 t_blb_n<5> vdd hvtpfet l=6e-08 w=8e-07 $X=19547 $Y=50503 $D=636
M2059 1261 221 223 vdd hvtpfet l=6e-08 w=8e-07 $X=19635 $Y=5556 $D=636
M2060 221 b_cb<1> vdd vdd hvtpfet l=6e-08 w=4e-07 $X=19635 $Y=10611 $D=636
M2061 219 221 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=19635 $Y=12911 $D=636
M2062 220 222 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=19635 $Y=37822 $D=636
M2063 222 t_cb<1> vdd vdd hvtpfet l=6e-08 w=4e-07 $X=19635 $Y=40122 $D=636
M2064 1262 222 224 vdd hvtpfet l=6e-08 w=8e-07 $X=19635 $Y=44777 $D=636
M2065 612 vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=19705 $Y=15090 $D=636
M2066 613 vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=19705 $Y=16110 $D=636
M2067 630 vdd vdd vdd hvtpfet l=6e-08 w=6e-07 $X=19730 $Y=18290 $D=636
M2068 vdd vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=19750 $Y=35893 $D=636
M2069 vdd vdd 609 vdd hvtpfet l=6e-08 w=6e-07 $X=19783 $Y=27488 $D=636
M2070 vdd vdd vdd vdd hvtpfet l=1e-07 w=2e-07 $X=19785 $Y=36723 $D=636
M2071 vdd vdd vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=19794 $Y=19812 $D=636
M2072 vdd vdd vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=19794 $Y=20072 $D=636
M2073 vdd vdd vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=19794 $Y=21162 $D=636
M2074 vdd vdd vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=19794 $Y=21422 $D=636
M2075 vdd vdd vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=19794 $Y=21682 $D=636
M2076 vdd vdd vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=19794 $Y=21942 $D=636
M2077 vdd vdd vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=19794 $Y=22762 $D=636
M2078 vdd vdd vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=19794 $Y=23879 $D=636
M2079 vdd vdd vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=19794 $Y=24139 $D=636
M2080 vdd vdd vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=19794 $Y=24399 $D=636
M2081 vdd vdd vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=19794 $Y=24659 $D=636
M2082 vdd 219 b_blb<5> vdd hvtpfet l=6e-08 w=8e-07 $X=19807 $Y=-170 $D=636
M2083 vdd 220 t_blb<5> vdd hvtpfet l=6e-08 w=8e-07 $X=19807 $Y=50503 $D=636
M2084 vdd 11 1261 vdd hvtpfet l=6e-08 w=8e-07 $X=19895 $Y=5556 $D=636
M2085 vdd b_mb<1> 221 vdd hvtpfet l=6e-08 w=4e-07 $X=19895 $Y=10611 $D=636
M2086 vdd 13 219 vdd hvtpfet l=6e-08 w=4e-07 $X=19895 $Y=12911 $D=636
M2087 vdd 14 220 vdd hvtpfet l=6e-08 w=4e-07 $X=19895 $Y=37822 $D=636
M2088 vdd t_mb<1> 222 vdd hvtpfet l=6e-08 w=4e-07 $X=19895 $Y=40122 $D=636
M2089 vdd 11 1262 vdd hvtpfet l=6e-08 w=8e-07 $X=19895 $Y=44777 $D=636
M2090 vdd vdd 630 vdd hvtpfet l=6e-08 w=6e-07 $X=19990 $Y=18290 $D=636
M2091 vdd vdd vdd vdd hvtpfet l=6e-08 w=6e-07 $X=20043 $Y=29008 $D=636
M2092 vdd vdd 612 vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=20045 $Y=15090 $D=636
M2093 vdd vdd 613 vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=20045 $Y=16110 $D=636
M2094 vdd vdd vdd vdd hvtpfet l=1e-07 w=2e-07 $X=20085 $Y=36723 $D=636
M2095 vdd vdd vdd vdd hvtpfet l=7e-08 w=3.2e-07 $X=20090 $Y=32628 $D=636
M2096 vdd vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=20090 $Y=35893 $D=636
M2097 1263 20 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=20155 $Y=5556 $D=636
M2098 227 b_ma<1> vdd vdd hvtpfet l=6e-08 w=4e-07 $X=20155 $Y=10611 $D=636
M2099 229 22 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=20155 $Y=12911 $D=636
M2100 230 23 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=20155 $Y=37822 $D=636
M2101 228 t_ma<1> vdd vdd hvtpfet l=6e-08 w=4e-07 $X=20155 $Y=40122 $D=636
M2102 1264 20 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=20155 $Y=44777 $D=636
M2103 b_bla_n<5> 229 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=20243 $Y=-170 $D=636
M2104 t_bla_n<5> 230 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=20243 $Y=50503 $D=636
M2105 630 vdd vdd vdd hvtpfet l=6e-08 w=6e-07 $X=20250 $Y=18290 $D=636
M2106 631 vdd vdd vdd hvtpfet l=6e-08 w=8e-07 $X=20293 $Y=27288 $D=636
M2107 vdd vdd vdd vdd hvtpfet l=6e-08 w=6e-07 $X=20303 $Y=29008 $D=636
M2108 vdd vdd vdd vdd hvtpfet l=7e-08 w=3.2e-07 $X=20380 $Y=32628 $D=636
M2109 vdd vdd vdd vdd hvtpfet l=1e-07 w=2e-07 $X=20385 $Y=36723 $D=636
M2110 225 227 1263 vdd hvtpfet l=6e-08 w=8e-07 $X=20415 $Y=5556 $D=636
M2111 vdd b_ca<1> 227 vdd hvtpfet l=6e-08 w=4e-07 $X=20415 $Y=10611 $D=636
M2112 vdd 227 229 vdd hvtpfet l=6e-08 w=4e-07 $X=20415 $Y=12911 $D=636
M2113 vdd 228 230 vdd hvtpfet l=6e-08 w=4e-07 $X=20415 $Y=37822 $D=636
M2114 vdd t_ca<1> 228 vdd hvtpfet l=6e-08 w=4e-07 $X=20415 $Y=40122 $D=636
M2115 226 228 1264 vdd hvtpfet l=6e-08 w=8e-07 $X=20415 $Y=44777 $D=636
M2116 vdd vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=20430 $Y=35893 $D=636
M2117 325 227 b_bla<5> vdd hvtpfet l=6e-08 w=3e-07 $X=20500 $Y=1094 $D=636
M2118 b_bla<5> 227 325 vdd hvtpfet l=6e-08 w=3e-07 $X=20500 $Y=1354 $D=636
M2119 b_bla_n<5> 227 326 vdd hvtpfet l=6e-08 w=3e-07 $X=20500 $Y=1864 $D=636
M2120 326 227 b_bla_n<5> vdd hvtpfet l=6e-08 w=3e-07 $X=20500 $Y=2124 $D=636
M2121 t_bla_n<5> 228 326 vdd hvtpfet l=6e-08 w=3e-07 $X=20500 $Y=48949 $D=636
M2122 326 228 t_bla_n<5> vdd hvtpfet l=6e-08 w=3e-07 $X=20500 $Y=49209 $D=636
M2123 325 228 t_bla<5> vdd hvtpfet l=6e-08 w=3e-07 $X=20500 $Y=49719 $D=636
M2124 t_bla<5> 228 325 vdd hvtpfet l=6e-08 w=3e-07 $X=20500 $Y=49979 $D=636
M2125 b_bla<5> 229 b_bla_n<5> vdd hvtpfet l=6e-08 w=8e-07 $X=20503 $Y=-170 $D=636
M2126 t_bla<5> 230 t_bla_n<5> vdd hvtpfet l=6e-08 w=8e-07 $X=20503 $Y=50503 $D=636
M2127 vdd vdd 630 vdd hvtpfet l=6e-08 w=6e-07 $X=20510 $Y=18290 $D=636
M2128 vdd vdd 631 vdd hvtpfet l=6e-08 w=8e-07 $X=20553 $Y=27288 $D=636
M2129 vdd vdd vdd vdd hvtpfet l=6e-08 w=6e-07 $X=20563 $Y=29008 $D=636
M2130 628 vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=20635 $Y=15090 $D=636
M2131 629 vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=20635 $Y=16110 $D=636
M2132 vdd vdd vdd vdd hvtpfet l=1e-07 w=6e-07 $X=20660 $Y=32628 $D=636
M2133 vdd vdd vdd vdd hvtpfet l=1e-07 w=2e-07 $X=20685 $Y=36723 $D=636
M2134 vdd 229 b_bla<5> vdd hvtpfet l=6e-08 w=8e-07 $X=20763 $Y=-170 $D=636
M2135 vdd 230 t_bla<5> vdd hvtpfet l=6e-08 w=8e-07 $X=20763 $Y=50503 $D=636
M2136 630 vdd vdd vdd hvtpfet l=6e-08 w=6e-07 $X=20770 $Y=18290 $D=636
M2137 vdd vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=20770 $Y=35893 $D=636
M2138 631 vdd vdd vdd hvtpfet l=6e-08 w=8e-07 $X=20813 $Y=27288 $D=636
M2139 vdd vdd vdd vdd hvtpfet l=6e-08 w=6e-07 $X=20823 $Y=29008 $D=636
M2140 vdd vdd vdd vdd hvtpfet l=1e-07 w=6e-07 $X=20960 $Y=32628 $D=636
M2141 vdd vdd 628 vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=20975 $Y=15090 $D=636
M2142 vdd vdd 629 vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=20975 $Y=16110 $D=636
M2143 vdd vdd 630 vdd hvtpfet l=6e-08 w=6e-07 $X=21030 $Y=18290 $D=636
M2144 vdd vdd 631 vdd hvtpfet l=6e-08 w=8e-07 $X=21073 $Y=27288 $D=636
M2145 vdd vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=21110 $Y=35893 $D=636
M2146 b_bla<4> 233 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=21197 $Y=-170 $D=636
M2147 t_bla<4> 234 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=21197 $Y=50503 $D=636
M2148 325 231 b_bla<4> vdd hvtpfet l=6e-08 w=3e-07 $X=21220 $Y=1094 $D=636
M2149 b_bla<4> 231 325 vdd hvtpfet l=6e-08 w=3e-07 $X=21220 $Y=1354 $D=636
M2150 b_bla_n<4> 231 326 vdd hvtpfet l=6e-08 w=3e-07 $X=21220 $Y=1864 $D=636
M2151 326 231 b_bla_n<4> vdd hvtpfet l=6e-08 w=3e-07 $X=21220 $Y=2124 $D=636
M2152 t_bla_n<4> 232 326 vdd hvtpfet l=6e-08 w=3e-07 $X=21220 $Y=48949 $D=636
M2153 326 232 t_bla_n<4> vdd hvtpfet l=6e-08 w=3e-07 $X=21220 $Y=49209 $D=636
M2154 325 232 t_bla<4> vdd hvtpfet l=6e-08 w=3e-07 $X=21220 $Y=49719 $D=636
M2155 t_bla<4> 232 325 vdd hvtpfet l=6e-08 w=3e-07 $X=21220 $Y=49979 $D=636
M2156 vdd vdd vdd vdd hvtpfet l=1e-07 w=2e-07 $X=21235 $Y=36723 $D=636
M2157 vdd vdd vdd vdd hvtpfet l=1e-07 w=6e-07 $X=21260 $Y=32628 $D=636
M2158 vdd vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=21450 $Y=35893 $D=636
M2159 b_bla_n<4> 233 b_bla<4> vdd hvtpfet l=6e-08 w=8e-07 $X=21457 $Y=-170 $D=636
M2160 t_bla_n<4> 234 t_bla<4> vdd hvtpfet l=6e-08 w=8e-07 $X=21457 $Y=50503 $D=636
M2161 vdd vdd vdd vdd hvtpfet l=1e-07 w=2e-07 $X=21535 $Y=36723 $D=636
M2162 654 vdd vdd vdd hvtpfet l=6e-08 w=5e-07 $X=21540 $Y=18290 $D=636
M2163 1269 231 235 vdd hvtpfet l=6e-08 w=8e-07 $X=21545 $Y=5556 $D=636
M2164 231 b_ca<0> vdd vdd hvtpfet l=6e-08 w=4e-07 $X=21545 $Y=10611 $D=636
M2165 233 231 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=21545 $Y=12911 $D=636
M2166 234 232 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=21545 $Y=37822 $D=636
M2167 232 t_ca<0> vdd vdd hvtpfet l=6e-08 w=4e-07 $X=21545 $Y=40122 $D=636
M2168 1270 232 236 vdd hvtpfet l=6e-08 w=8e-07 $X=21545 $Y=44777 $D=636
M2169 vdd vdd vdd vdd hvtpfet l=7e-08 w=3.2e-07 $X=21570 $Y=32628 $D=636
M2170 643 vdd vdd vdd hvtpfet l=6e-08 w=6e-07 $X=21593 $Y=27488 $D=636
M2171 vdd 233 b_bla_n<4> vdd hvtpfet l=6e-08 w=8e-07 $X=21717 $Y=-170 $D=636
M2172 vdd 234 t_bla_n<4> vdd hvtpfet l=6e-08 w=8e-07 $X=21717 $Y=50503 $D=636
M2173 vdd vdd vdd vdd hvtpfet l=6e-08 w=6e-07 $X=21733 $Y=29008 $D=636
M2174 vdd vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=21790 $Y=35893 $D=636
M2175 vdd vdd 654 vdd hvtpfet l=6e-08 w=5e-07 $X=21800 $Y=18290 $D=636
M2176 vdd 20 1269 vdd hvtpfet l=6e-08 w=8e-07 $X=21805 $Y=5556 $D=636
M2177 vdd b_ma<1> 231 vdd hvtpfet l=6e-08 w=4e-07 $X=21805 $Y=10611 $D=636
M2178 vdd 22 233 vdd hvtpfet l=6e-08 w=4e-07 $X=21805 $Y=12911 $D=636
M2179 vdd 23 234 vdd hvtpfet l=6e-08 w=4e-07 $X=21805 $Y=37822 $D=636
M2180 vdd t_ma<1> 232 vdd hvtpfet l=6e-08 w=4e-07 $X=21805 $Y=40122 $D=636
M2181 vdd 20 1270 vdd hvtpfet l=6e-08 w=8e-07 $X=21805 $Y=44777 $D=636
M2182 vdd vdd vdd vdd hvtpfet l=1e-07 w=2e-07 $X=21835 $Y=36723 $D=636
M2183 vdd vdd vdd vdd hvtpfet l=7e-08 w=3.2e-07 $X=21860 $Y=32628 $D=636
M2184 vdd vdd vdd vdd hvtpfet l=6e-08 w=6e-07 $X=21993 $Y=29008 $D=636
M2185 654 vdd vdd vdd hvtpfet l=6e-08 w=5e-07 $X=22060 $Y=18290 $D=636
M2186 1271 11 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=22065 $Y=5556 $D=636
M2187 237 b_mb<1> vdd vdd hvtpfet l=6e-08 w=4e-07 $X=22065 $Y=10611 $D=636
M2188 241 13 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=22065 $Y=12911 $D=636
M2189 242 14 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=22065 $Y=37822 $D=636
M2190 238 t_mb<1> vdd vdd hvtpfet l=6e-08 w=4e-07 $X=22065 $Y=40122 $D=636
M2191 1272 11 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=22065 $Y=44777 $D=636
M2192 vdd vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=22130 $Y=35893 $D=636
M2193 vdd vdd vdd vdd hvtpfet l=1e-07 w=2e-07 $X=22135 $Y=36723 $D=636
M2194 b_blb<4> 241 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=22153 $Y=-170 $D=636
M2195 t_blb<4> 242 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=22153 $Y=50503 $D=636
M2196 644 vdd vdd vdd hvtpfet l=6e-08 w=4e-07 $X=22265 $Y=21427 $D=636
M2197 645 vdd vdd vdd hvtpfet l=6e-08 w=4e-07 $X=22265 $Y=23694 $D=636
M2198 646 vdd vdd vdd hvtpfet l=6e-08 w=4e-07 $X=22265 $Y=24394 $D=636
M2199 647 vdd vdd vdd hvtpfet l=6e-08 w=4e-07 $X=22265 $Y=24904 $D=636
M2200 vdd vdd 654 vdd hvtpfet l=6e-08 w=5e-07 $X=22320 $Y=18290 $D=636
M2201 239 237 1271 vdd hvtpfet l=6e-08 w=8e-07 $X=22325 $Y=5556 $D=636
M2202 vdd b_cb<0> 237 vdd hvtpfet l=6e-08 w=4e-07 $X=22325 $Y=10611 $D=636
M2203 vdd 237 241 vdd hvtpfet l=6e-08 w=4e-07 $X=22325 $Y=12911 $D=636
M2204 vdd 238 242 vdd hvtpfet l=6e-08 w=4e-07 $X=22325 $Y=37822 $D=636
M2205 vdd t_cb<0> 238 vdd hvtpfet l=6e-08 w=4e-07 $X=22325 $Y=40122 $D=636
M2206 240 238 1272 vdd hvtpfet l=6e-08 w=8e-07 $X=22325 $Y=44777 $D=636
M2207 296 237 b_blb<4> vdd hvtpfet l=6e-08 w=3e-07 $X=22410 $Y=1094 $D=636
M2208 b_blb<4> 237 296 vdd hvtpfet l=6e-08 w=3e-07 $X=22410 $Y=1354 $D=636
M2209 b_blb_n<4> 237 297 vdd hvtpfet l=6e-08 w=3e-07 $X=22410 $Y=1864 $D=636
M2210 297 237 b_blb_n<4> vdd hvtpfet l=6e-08 w=3e-07 $X=22410 $Y=2124 $D=636
M2211 t_blb_n<4> 238 297 vdd hvtpfet l=6e-08 w=3e-07 $X=22410 $Y=48949 $D=636
M2212 297 238 t_blb_n<4> vdd hvtpfet l=6e-08 w=3e-07 $X=22410 $Y=49209 $D=636
M2213 296 238 t_blb<4> vdd hvtpfet l=6e-08 w=3e-07 $X=22410 $Y=49719 $D=636
M2214 t_blb<4> 238 296 vdd hvtpfet l=6e-08 w=3e-07 $X=22410 $Y=49979 $D=636
M2215 b_blb_n<4> 241 b_blb<4> vdd hvtpfet l=6e-08 w=8e-07 $X=22413 $Y=-170 $D=636
M2216 t_blb_n<4> 242 t_blb<4> vdd hvtpfet l=6e-08 w=8e-07 $X=22413 $Y=50503 $D=636
M2217 vdd vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=22575 $Y=35893 $D=636
M2218 vdd 241 b_blb_n<4> vdd hvtpfet l=6e-08 w=8e-07 $X=22673 $Y=-170 $D=636
M2219 vdd 242 t_blb_n<4> vdd hvtpfet l=6e-08 w=8e-07 $X=22673 $Y=50503 $D=636
M2220 b_blb_n<3> 243 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=23107 $Y=-170 $D=636
M2221 t_blb_n<3> 244 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=23107 $Y=50503 $D=636
M2222 vdd vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=23125 $Y=35893 $D=636
M2223 296 245 b_blb<3> vdd hvtpfet l=6e-08 w=3e-07 $X=23130 $Y=1094 $D=636
M2224 b_blb<3> 245 296 vdd hvtpfet l=6e-08 w=3e-07 $X=23130 $Y=1354 $D=636
M2225 b_blb_n<3> 245 297 vdd hvtpfet l=6e-08 w=3e-07 $X=23130 $Y=1864 $D=636
M2226 297 245 b_blb_n<3> vdd hvtpfet l=6e-08 w=3e-07 $X=23130 $Y=2124 $D=636
M2227 t_blb_n<3> 246 297 vdd hvtpfet l=6e-08 w=3e-07 $X=23130 $Y=48949 $D=636
M2228 297 246 t_blb_n<3> vdd hvtpfet l=6e-08 w=3e-07 $X=23130 $Y=49209 $D=636
M2229 296 246 t_blb<3> vdd hvtpfet l=6e-08 w=3e-07 $X=23130 $Y=49719 $D=636
M2230 t_blb<3> 246 296 vdd hvtpfet l=6e-08 w=3e-07 $X=23130 $Y=49979 $D=636
M2231 667 vdd vdd vdd hvtpfet l=6e-08 w=4e-07 $X=23175 $Y=21427 $D=636
M2232 668 vdd vdd vdd hvtpfet l=6e-08 w=4e-07 $X=23175 $Y=23694 $D=636
M2233 669 vdd vdd vdd hvtpfet l=6e-08 w=4e-07 $X=23175 $Y=24394 $D=636
M2234 670 vdd vdd vdd hvtpfet l=6e-08 w=4e-07 $X=23175 $Y=24904 $D=636
M2235 b_blb<3> 243 b_blb_n<3> vdd hvtpfet l=6e-08 w=8e-07 $X=23367 $Y=-170 $D=636
M2236 t_blb<3> 244 t_blb_n<3> vdd hvtpfet l=6e-08 w=8e-07 $X=23367 $Y=50503 $D=636
M2237 1277 245 247 vdd hvtpfet l=6e-08 w=8e-07 $X=23455 $Y=5556 $D=636
M2238 245 b_cb<3> vdd vdd hvtpfet l=6e-08 w=4e-07 $X=23455 $Y=10611 $D=636
M2239 243 245 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=23455 $Y=12911 $D=636
M2240 244 246 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=23455 $Y=37822 $D=636
M2241 246 t_cb<3> vdd vdd hvtpfet l=6e-08 w=4e-07 $X=23455 $Y=40122 $D=636
M2242 1278 246 248 vdd hvtpfet l=6e-08 w=8e-07 $X=23455 $Y=44777 $D=636
M2243 682 vdd vdd vdd hvtpfet l=6e-08 w=5e-07 $X=23460 $Y=18290 $D=636
M2244 vdd vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=23570 $Y=35893 $D=636
M2245 vdd vdd vdd vdd hvtpfet l=1e-07 w=2e-07 $X=23605 $Y=36723 $D=636
M2246 vdd 243 b_blb<3> vdd hvtpfet l=6e-08 w=8e-07 $X=23627 $Y=-170 $D=636
M2247 vdd 244 t_blb<3> vdd hvtpfet l=6e-08 w=8e-07 $X=23627 $Y=50503 $D=636
M2248 vdd 11 1277 vdd hvtpfet l=6e-08 w=8e-07 $X=23715 $Y=5556 $D=636
M2249 vdd b_mb<0> 245 vdd hvtpfet l=6e-08 w=4e-07 $X=23715 $Y=10611 $D=636
M2250 vdd 13 243 vdd hvtpfet l=6e-08 w=4e-07 $X=23715 $Y=12911 $D=636
M2251 vdd 14 244 vdd hvtpfet l=6e-08 w=4e-07 $X=23715 $Y=37822 $D=636
M2252 vdd t_mb<0> 246 vdd hvtpfet l=6e-08 w=4e-07 $X=23715 $Y=40122 $D=636
M2253 vdd 11 1278 vdd hvtpfet l=6e-08 w=8e-07 $X=23715 $Y=44777 $D=636
M2254 vdd vdd 682 vdd hvtpfet l=6e-08 w=5e-07 $X=23720 $Y=18290 $D=636
M2255 vdd vdd vdd vdd hvtpfet l=6e-08 w=6e-07 $X=23787 $Y=29008 $D=636
M2256 vdd vdd vdd vdd hvtpfet l=1e-07 w=2e-07 $X=23905 $Y=36723 $D=636
M2257 vdd vdd vdd vdd hvtpfet l=7e-08 w=3.2e-07 $X=23910 $Y=32628 $D=636
M2258 vdd vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=23910 $Y=35893 $D=636
M2259 1279 20 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=23975 $Y=5556 $D=636
M2260 253 b_ma<0> vdd vdd hvtpfet l=6e-08 w=4e-07 $X=23975 $Y=10611 $D=636
M2261 257 22 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=23975 $Y=12911 $D=636
M2262 258 23 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=23975 $Y=37822 $D=636
M2263 254 t_ma<0> vdd vdd hvtpfet l=6e-08 w=4e-07 $X=23975 $Y=40122 $D=636
M2264 1280 20 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=23975 $Y=44777 $D=636
M2265 682 vdd vdd vdd hvtpfet l=6e-08 w=5e-07 $X=23980 $Y=18290 $D=636
M2266 vdd vdd vdd vdd hvtpfet l=6e-08 w=6e-07 $X=24047 $Y=29008 $D=636
M2267 b_bla_n<3> 257 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=24063 $Y=-170 $D=636
M2268 t_bla_n<3> 258 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=24063 $Y=50503 $D=636
M2269 vdd vdd 681 vdd hvtpfet l=6e-08 w=6e-07 $X=24187 $Y=27488 $D=636
M2270 vdd vdd vdd vdd hvtpfet l=7e-08 w=3.2e-07 $X=24200 $Y=32628 $D=636
M2271 vdd vdd vdd vdd hvtpfet l=1e-07 w=2e-07 $X=24205 $Y=36723 $D=636
M2272 251 253 1279 vdd hvtpfet l=6e-08 w=8e-07 $X=24235 $Y=5556 $D=636
M2273 vdd b_ca<3> 253 vdd hvtpfet l=6e-08 w=4e-07 $X=24235 $Y=10611 $D=636
M2274 vdd 253 257 vdd hvtpfet l=6e-08 w=4e-07 $X=24235 $Y=12911 $D=636
M2275 vdd 254 258 vdd hvtpfet l=6e-08 w=4e-07 $X=24235 $Y=37822 $D=636
M2276 vdd t_ca<3> 254 vdd hvtpfet l=6e-08 w=4e-07 $X=24235 $Y=40122 $D=636
M2277 252 254 1280 vdd hvtpfet l=6e-08 w=8e-07 $X=24235 $Y=44777 $D=636
M2278 vdd vdd 682 vdd hvtpfet l=6e-08 w=5e-07 $X=24240 $Y=18290 $D=636
M2279 vdd vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=24250 $Y=35893 $D=636
M2280 325 253 b_bla<3> vdd hvtpfet l=6e-08 w=3e-07 $X=24320 $Y=1094 $D=636
M2281 b_bla<3> 253 325 vdd hvtpfet l=6e-08 w=3e-07 $X=24320 $Y=1354 $D=636
M2282 b_bla_n<3> 253 326 vdd hvtpfet l=6e-08 w=3e-07 $X=24320 $Y=1864 $D=636
M2283 326 253 b_bla_n<3> vdd hvtpfet l=6e-08 w=3e-07 $X=24320 $Y=2124 $D=636
M2284 t_bla_n<3> 254 326 vdd hvtpfet l=6e-08 w=3e-07 $X=24320 $Y=48949 $D=636
M2285 326 254 t_bla_n<3> vdd hvtpfet l=6e-08 w=3e-07 $X=24320 $Y=49209 $D=636
M2286 325 254 t_bla<3> vdd hvtpfet l=6e-08 w=3e-07 $X=24320 $Y=49719 $D=636
M2287 t_bla<3> 254 325 vdd hvtpfet l=6e-08 w=3e-07 $X=24320 $Y=49979 $D=636
M2288 b_bla<3> 257 b_bla_n<3> vdd hvtpfet l=6e-08 w=8e-07 $X=24323 $Y=-170 $D=636
M2289 t_bla<3> 258 t_bla_n<3> vdd hvtpfet l=6e-08 w=8e-07 $X=24323 $Y=50503 $D=636
M2290 vdd vdd vdd vdd hvtpfet l=1e-07 w=6e-07 $X=24480 $Y=32628 $D=636
M2291 vdd vdd vdd vdd hvtpfet l=1e-07 w=2e-07 $X=24505 $Y=36723 $D=636
M2292 vdd 257 b_bla<3> vdd hvtpfet l=6e-08 w=8e-07 $X=24583 $Y=-170 $D=636
M2293 vdd 258 t_bla<3> vdd hvtpfet l=6e-08 w=8e-07 $X=24583 $Y=50503 $D=636
M2294 vdd vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=24590 $Y=35893 $D=636
M2295 703 vdd vdd vdd hvtpfet l=6e-08 w=8e-07 $X=24707 $Y=27288 $D=636
M2296 697 vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=24725 $Y=15090 $D=636
M2297 698 vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=24725 $Y=16110 $D=636
M2298 713 vdd vdd vdd hvtpfet l=6e-08 w=6e-07 $X=24750 $Y=18290 $D=636
M2299 vdd vdd vdd vdd hvtpfet l=1e-07 w=6e-07 $X=24780 $Y=32628 $D=636
M2300 vdd vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=24930 $Y=35893 $D=636
M2301 vdd vdd vdd vdd hvtpfet l=6e-08 w=6e-07 $X=24957 $Y=29008 $D=636
M2302 vdd vdd 703 vdd hvtpfet l=6e-08 w=8e-07 $X=24967 $Y=27288 $D=636
M2303 vdd vdd 713 vdd hvtpfet l=6e-08 w=6e-07 $X=25010 $Y=18290 $D=636
M2304 b_bla<2> 261 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=25017 $Y=-170 $D=636
M2305 t_bla<2> 262 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=25017 $Y=50503 $D=636
M2306 325 259 b_bla<2> vdd hvtpfet l=6e-08 w=3e-07 $X=25040 $Y=1094 $D=636
M2307 b_bla<2> 259 325 vdd hvtpfet l=6e-08 w=3e-07 $X=25040 $Y=1354 $D=636
M2308 b_bla_n<2> 259 326 vdd hvtpfet l=6e-08 w=3e-07 $X=25040 $Y=1864 $D=636
M2309 326 259 b_bla_n<2> vdd hvtpfet l=6e-08 w=3e-07 $X=25040 $Y=2124 $D=636
M2310 t_bla_n<2> 260 326 vdd hvtpfet l=6e-08 w=3e-07 $X=25040 $Y=48949 $D=636
M2311 326 260 t_bla_n<2> vdd hvtpfet l=6e-08 w=3e-07 $X=25040 $Y=49209 $D=636
M2312 325 260 t_bla<2> vdd hvtpfet l=6e-08 w=3e-07 $X=25040 $Y=49719 $D=636
M2313 t_bla<2> 260 325 vdd hvtpfet l=6e-08 w=3e-07 $X=25040 $Y=49979 $D=636
M2314 vdd vdd vdd vdd hvtpfet l=1e-07 w=2e-07 $X=25055 $Y=36723 $D=636
M2315 vdd vdd 697 vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=25065 $Y=15090 $D=636
M2316 vdd vdd 698 vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=25065 $Y=16110 $D=636
M2317 vdd vdd vdd vdd hvtpfet l=1e-07 w=6e-07 $X=25080 $Y=32628 $D=636
M2318 vdd vdd vdd vdd hvtpfet l=6e-08 w=6e-07 $X=25217 $Y=29008 $D=636
M2319 703 vdd vdd vdd hvtpfet l=6e-08 w=8e-07 $X=25227 $Y=27288 $D=636
M2320 713 vdd vdd vdd hvtpfet l=6e-08 w=6e-07 $X=25270 $Y=18290 $D=636
M2321 vdd vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=25270 $Y=35893 $D=636
M2322 b_bla_n<2> 261 b_bla<2> vdd hvtpfet l=6e-08 w=8e-07 $X=25277 $Y=-170 $D=636
M2323 t_bla_n<2> 262 t_bla<2> vdd hvtpfet l=6e-08 w=8e-07 $X=25277 $Y=50503 $D=636
M2324 vdd vdd vdd vdd hvtpfet l=1e-07 w=2e-07 $X=25355 $Y=36723 $D=636
M2325 1285 259 263 vdd hvtpfet l=6e-08 w=8e-07 $X=25365 $Y=5556 $D=636
M2326 259 b_ca<2> vdd vdd hvtpfet l=6e-08 w=4e-07 $X=25365 $Y=10611 $D=636
M2327 261 259 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=25365 $Y=12911 $D=636
M2328 262 260 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=25365 $Y=37822 $D=636
M2329 260 t_ca<2> vdd vdd hvtpfet l=6e-08 w=4e-07 $X=25365 $Y=40122 $D=636
M2330 1286 260 264 vdd hvtpfet l=6e-08 w=8e-07 $X=25365 $Y=44777 $D=636
M2331 vdd vdd vdd vdd hvtpfet l=7e-08 w=3.2e-07 $X=25390 $Y=32628 $D=636
M2332 vdd vdd vdd vdd hvtpfet l=6e-08 w=6e-07 $X=25477 $Y=29008 $D=636
M2333 vdd vdd 703 vdd hvtpfet l=6e-08 w=8e-07 $X=25487 $Y=27288 $D=636
M2334 vdd vdd 713 vdd hvtpfet l=6e-08 w=6e-07 $X=25530 $Y=18290 $D=636
M2335 vdd 261 b_bla_n<2> vdd hvtpfet l=6e-08 w=8e-07 $X=25537 $Y=-170 $D=636
M2336 vdd 262 t_bla_n<2> vdd hvtpfet l=6e-08 w=8e-07 $X=25537 $Y=50503 $D=636
M2337 vdd vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=25610 $Y=35893 $D=636
M2338 vdd 20 1285 vdd hvtpfet l=6e-08 w=8e-07 $X=25625 $Y=5556 $D=636
M2339 vdd b_ma<0> 259 vdd hvtpfet l=6e-08 w=4e-07 $X=25625 $Y=10611 $D=636
M2340 vdd 22 261 vdd hvtpfet l=6e-08 w=4e-07 $X=25625 $Y=12911 $D=636
M2341 vdd 23 262 vdd hvtpfet l=6e-08 w=4e-07 $X=25625 $Y=37822 $D=636
M2342 vdd t_ma<0> 260 vdd hvtpfet l=6e-08 w=4e-07 $X=25625 $Y=40122 $D=636
M2343 vdd 20 1286 vdd hvtpfet l=6e-08 w=8e-07 $X=25625 $Y=44777 $D=636
M2344 711 vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=25655 $Y=15090 $D=636
M2345 712 vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=25655 $Y=16110 $D=636
M2346 vdd vdd vdd vdd hvtpfet l=1e-07 w=2e-07 $X=25655 $Y=36723 $D=636
M2347 vdd vdd vdd vdd hvtpfet l=7e-08 w=3.2e-07 $X=25680 $Y=32628 $D=636
M2348 vdd vdd vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=25726 $Y=19812 $D=636
M2349 vdd vdd vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=25726 $Y=20072 $D=636
M2350 vdd vdd vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=25726 $Y=21162 $D=636
M2351 vdd vdd vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=25726 $Y=21422 $D=636
M2352 vdd vdd vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=25726 $Y=21682 $D=636
M2353 vdd vdd vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=25726 $Y=21942 $D=636
M2354 vdd vdd vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=25726 $Y=22762 $D=636
M2355 vdd vdd vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=25726 $Y=23879 $D=636
M2356 vdd vdd vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=25726 $Y=24139 $D=636
M2357 vdd vdd vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=25726 $Y=24399 $D=636
M2358 vdd vdd vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=25726 $Y=24659 $D=636
M2359 vdd vdd vdd vdd hvtpfet l=6e-08 w=6e-07 $X=25737 $Y=29008 $D=636
M2360 713 vdd vdd vdd hvtpfet l=6e-08 w=6e-07 $X=25790 $Y=18290 $D=636
M2361 1287 11 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=25885 $Y=5556 $D=636
M2362 265 b_mb<0> vdd vdd hvtpfet l=6e-08 w=4e-07 $X=25885 $Y=10611 $D=636
M2363 269 13 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=25885 $Y=12911 $D=636
M2364 270 14 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=25885 $Y=37822 $D=636
M2365 266 t_mb<0> vdd vdd hvtpfet l=6e-08 w=4e-07 $X=25885 $Y=40122 $D=636
M2366 1288 11 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=25885 $Y=44777 $D=636
M2367 vdd vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=25950 $Y=35893 $D=636
M2368 vdd vdd vdd vdd hvtpfet l=1e-07 w=2e-07 $X=25955 $Y=36723 $D=636
M2369 b_blb<2> 269 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=25973 $Y=-170 $D=636
M2370 t_blb<2> 270 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=25973 $Y=50503 $D=636
M2371 vdd vdd 711 vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=25995 $Y=15090 $D=636
M2372 vdd vdd 712 vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=25995 $Y=16110 $D=636
M2373 720 vdd vdd vdd hvtpfet l=6e-08 w=6e-07 $X=25997 $Y=27488 $D=636
M2374 vdd vdd 713 vdd hvtpfet l=6e-08 w=6e-07 $X=26050 $Y=18290 $D=636
M2375 267 265 1287 vdd hvtpfet l=6e-08 w=8e-07 $X=26145 $Y=5556 $D=636
M2376 vdd b_cb<2> 265 vdd hvtpfet l=6e-08 w=4e-07 $X=26145 $Y=10611 $D=636
M2377 vdd 265 269 vdd hvtpfet l=6e-08 w=4e-07 $X=26145 $Y=12911 $D=636
M2378 vdd 266 270 vdd hvtpfet l=6e-08 w=4e-07 $X=26145 $Y=37822 $D=636
M2379 vdd t_cb<2> 266 vdd hvtpfet l=6e-08 w=4e-07 $X=26145 $Y=40122 $D=636
M2380 268 266 1288 vdd hvtpfet l=6e-08 w=8e-07 $X=26145 $Y=44777 $D=636
M2381 296 265 b_blb<2> vdd hvtpfet l=6e-08 w=3e-07 $X=26230 $Y=1094 $D=636
M2382 b_blb<2> 265 296 vdd hvtpfet l=6e-08 w=3e-07 $X=26230 $Y=1354 $D=636
M2383 b_blb_n<2> 265 297 vdd hvtpfet l=6e-08 w=3e-07 $X=26230 $Y=1864 $D=636
M2384 297 265 b_blb_n<2> vdd hvtpfet l=6e-08 w=3e-07 $X=26230 $Y=2124 $D=636
M2385 t_blb_n<2> 266 297 vdd hvtpfet l=6e-08 w=3e-07 $X=26230 $Y=48949 $D=636
M2386 297 266 t_blb_n<2> vdd hvtpfet l=6e-08 w=3e-07 $X=26230 $Y=49209 $D=636
M2387 296 266 t_blb<2> vdd hvtpfet l=6e-08 w=3e-07 $X=26230 $Y=49719 $D=636
M2388 t_blb<2> 266 296 vdd hvtpfet l=6e-08 w=3e-07 $X=26230 $Y=49979 $D=636
M2389 b_blb_n<2> 269 b_blb<2> vdd hvtpfet l=6e-08 w=8e-07 $X=26233 $Y=-170 $D=636
M2390 t_blb_n<2> 270 t_blb<2> vdd hvtpfet l=6e-08 w=8e-07 $X=26233 $Y=50503 $D=636
M2391 vdd vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=26395 $Y=35893 $D=636
M2392 vdd 269 b_blb_n<2> vdd hvtpfet l=6e-08 w=8e-07 $X=26493 $Y=-170 $D=636
M2393 vdd 270 t_blb_n<2> vdd hvtpfet l=6e-08 w=8e-07 $X=26493 $Y=50503 $D=636
M2394 b_blb_n<1> 271 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=26927 $Y=-170 $D=636
M2395 t_blb_n<1> 272 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=26927 $Y=50503 $D=636
M2396 vdd vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=26945 $Y=35893 $D=636
M2397 296 273 b_blb<1> vdd hvtpfet l=6e-08 w=3e-07 $X=26950 $Y=1094 $D=636
M2398 b_blb<1> 273 296 vdd hvtpfet l=6e-08 w=3e-07 $X=26950 $Y=1354 $D=636
M2399 b_blb_n<1> 273 297 vdd hvtpfet l=6e-08 w=3e-07 $X=26950 $Y=1864 $D=636
M2400 297 273 b_blb_n<1> vdd hvtpfet l=6e-08 w=3e-07 $X=26950 $Y=2124 $D=636
M2401 t_blb_n<1> 274 297 vdd hvtpfet l=6e-08 w=3e-07 $X=26950 $Y=48949 $D=636
M2402 297 274 t_blb_n<1> vdd hvtpfet l=6e-08 w=3e-07 $X=26950 $Y=49209 $D=636
M2403 296 274 t_blb<1> vdd hvtpfet l=6e-08 w=3e-07 $X=26950 $Y=49719 $D=636
M2404 t_blb<1> 274 296 vdd hvtpfet l=6e-08 w=3e-07 $X=26950 $Y=49979 $D=636
M2405 b_blb<1> 271 b_blb_n<1> vdd hvtpfet l=6e-08 w=8e-07 $X=27187 $Y=-170 $D=636
M2406 t_blb<1> 272 t_blb_n<1> vdd hvtpfet l=6e-08 w=8e-07 $X=27187 $Y=50503 $D=636
M2407 1293 273 275 vdd hvtpfet l=6e-08 w=8e-07 $X=27275 $Y=5556 $D=636
M2408 273 b_cb<1> vdd vdd hvtpfet l=6e-08 w=4e-07 $X=27275 $Y=10611 $D=636
M2409 271 273 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=27275 $Y=12911 $D=636
M2410 272 274 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=27275 $Y=37822 $D=636
M2411 274 t_cb<1> vdd vdd hvtpfet l=6e-08 w=4e-07 $X=27275 $Y=40122 $D=636
M2412 1294 274 276 vdd hvtpfet l=6e-08 w=8e-07 $X=27275 $Y=44777 $D=636
M2413 736 vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=27345 $Y=15090 $D=636
M2414 737 vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=27345 $Y=16110 $D=636
M2415 754 vdd vdd vdd hvtpfet l=6e-08 w=6e-07 $X=27370 $Y=18290 $D=636
M2416 vdd vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=27390 $Y=35893 $D=636
M2417 vdd vdd 733 vdd hvtpfet l=6e-08 w=6e-07 $X=27423 $Y=27488 $D=636
M2418 vdd vdd vdd vdd hvtpfet l=1e-07 w=2e-07 $X=27425 $Y=36723 $D=636
M2419 vdd vdd vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=27434 $Y=19812 $D=636
M2420 vdd vdd vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=27434 $Y=20072 $D=636
M2421 vdd vdd vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=27434 $Y=21162 $D=636
M2422 vdd vdd vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=27434 $Y=21422 $D=636
M2423 vdd vdd vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=27434 $Y=21682 $D=636
M2424 vdd vdd vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=27434 $Y=21942 $D=636
M2425 vdd vdd vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=27434 $Y=22762 $D=636
M2426 vdd vdd vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=27434 $Y=23879 $D=636
M2427 vdd vdd vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=27434 $Y=24139 $D=636
M2428 vdd vdd vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=27434 $Y=24399 $D=636
M2429 vdd vdd vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=27434 $Y=24659 $D=636
M2430 vdd 271 b_blb<1> vdd hvtpfet l=6e-08 w=8e-07 $X=27447 $Y=-170 $D=636
M2431 vdd 272 t_blb<1> vdd hvtpfet l=6e-08 w=8e-07 $X=27447 $Y=50503 $D=636
M2432 vdd 11 1293 vdd hvtpfet l=6e-08 w=8e-07 $X=27535 $Y=5556 $D=636
M2433 vdd b_mb<0> 273 vdd hvtpfet l=6e-08 w=4e-07 $X=27535 $Y=10611 $D=636
M2434 vdd 13 271 vdd hvtpfet l=6e-08 w=4e-07 $X=27535 $Y=12911 $D=636
M2435 vdd 14 272 vdd hvtpfet l=6e-08 w=4e-07 $X=27535 $Y=37822 $D=636
M2436 vdd t_mb<0> 274 vdd hvtpfet l=6e-08 w=4e-07 $X=27535 $Y=40122 $D=636
M2437 vdd 11 1294 vdd hvtpfet l=6e-08 w=8e-07 $X=27535 $Y=44777 $D=636
M2438 vdd vdd 754 vdd hvtpfet l=6e-08 w=6e-07 $X=27630 $Y=18290 $D=636
M2439 vdd vdd vdd vdd hvtpfet l=6e-08 w=6e-07 $X=27683 $Y=29008 $D=636
M2440 vdd vdd 736 vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=27685 $Y=15090 $D=636
M2441 vdd vdd 737 vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=27685 $Y=16110 $D=636
M2442 vdd vdd vdd vdd hvtpfet l=1e-07 w=2e-07 $X=27725 $Y=36723 $D=636
M2443 vdd vdd vdd vdd hvtpfet l=7e-08 w=3.2e-07 $X=27730 $Y=32628 $D=636
M2444 vdd vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=27730 $Y=35893 $D=636
M2445 1295 20 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=27795 $Y=5556 $D=636
M2446 279 b_ma<0> vdd vdd hvtpfet l=6e-08 w=4e-07 $X=27795 $Y=10611 $D=636
M2447 281 22 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=27795 $Y=12911 $D=636
M2448 282 23 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=27795 $Y=37822 $D=636
M2449 280 t_ma<0> vdd vdd hvtpfet l=6e-08 w=4e-07 $X=27795 $Y=40122 $D=636
M2450 1296 20 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=27795 $Y=44777 $D=636
M2451 b_bla_n<1> 281 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=27883 $Y=-170 $D=636
M2452 t_bla_n<1> 282 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=27883 $Y=50503 $D=636
M2453 754 vdd vdd vdd hvtpfet l=6e-08 w=6e-07 $X=27890 $Y=18290 $D=636
M2454 755 vdd vdd vdd hvtpfet l=6e-08 w=8e-07 $X=27933 $Y=27288 $D=636
M2455 vdd vdd vdd vdd hvtpfet l=6e-08 w=6e-07 $X=27943 $Y=29008 $D=636
M2456 vdd vdd vdd vdd hvtpfet l=7e-08 w=3.2e-07 $X=28020 $Y=32628 $D=636
M2457 vdd vdd vdd vdd hvtpfet l=1e-07 w=2e-07 $X=28025 $Y=36723 $D=636
M2458 277 279 1295 vdd hvtpfet l=6e-08 w=8e-07 $X=28055 $Y=5556 $D=636
M2459 vdd b_ca<1> 279 vdd hvtpfet l=6e-08 w=4e-07 $X=28055 $Y=10611 $D=636
M2460 vdd 279 281 vdd hvtpfet l=6e-08 w=4e-07 $X=28055 $Y=12911 $D=636
M2461 vdd 280 282 vdd hvtpfet l=6e-08 w=4e-07 $X=28055 $Y=37822 $D=636
M2462 vdd t_ca<1> 280 vdd hvtpfet l=6e-08 w=4e-07 $X=28055 $Y=40122 $D=636
M2463 278 280 1296 vdd hvtpfet l=6e-08 w=8e-07 $X=28055 $Y=44777 $D=636
M2464 vdd vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=28070 $Y=35893 $D=636
M2465 325 279 b_bla<1> vdd hvtpfet l=6e-08 w=3e-07 $X=28140 $Y=1094 $D=636
M2466 b_bla<1> 279 325 vdd hvtpfet l=6e-08 w=3e-07 $X=28140 $Y=1354 $D=636
M2467 b_bla_n<1> 279 326 vdd hvtpfet l=6e-08 w=3e-07 $X=28140 $Y=1864 $D=636
M2468 326 279 b_bla_n<1> vdd hvtpfet l=6e-08 w=3e-07 $X=28140 $Y=2124 $D=636
M2469 t_bla_n<1> 280 326 vdd hvtpfet l=6e-08 w=3e-07 $X=28140 $Y=48949 $D=636
M2470 326 280 t_bla_n<1> vdd hvtpfet l=6e-08 w=3e-07 $X=28140 $Y=49209 $D=636
M2471 325 280 t_bla<1> vdd hvtpfet l=6e-08 w=3e-07 $X=28140 $Y=49719 $D=636
M2472 t_bla<1> 280 325 vdd hvtpfet l=6e-08 w=3e-07 $X=28140 $Y=49979 $D=636
M2473 b_bla<1> 281 b_bla_n<1> vdd hvtpfet l=6e-08 w=8e-07 $X=28143 $Y=-170 $D=636
M2474 t_bla<1> 282 t_bla_n<1> vdd hvtpfet l=6e-08 w=8e-07 $X=28143 $Y=50503 $D=636
M2475 vdd vdd 754 vdd hvtpfet l=6e-08 w=6e-07 $X=28150 $Y=18290 $D=636
M2476 vdd vdd 755 vdd hvtpfet l=6e-08 w=8e-07 $X=28193 $Y=27288 $D=636
M2477 vdd vdd vdd vdd hvtpfet l=6e-08 w=6e-07 $X=28203 $Y=29008 $D=636
M2478 752 vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=28275 $Y=15090 $D=636
M2479 753 vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=28275 $Y=16110 $D=636
M2480 vdd vdd vdd vdd hvtpfet l=1e-07 w=6e-07 $X=28300 $Y=32628 $D=636
M2481 vdd vdd vdd vdd hvtpfet l=1e-07 w=2e-07 $X=28325 $Y=36723 $D=636
M2482 vdd 281 b_bla<1> vdd hvtpfet l=6e-08 w=8e-07 $X=28403 $Y=-170 $D=636
M2483 vdd 282 t_bla<1> vdd hvtpfet l=6e-08 w=8e-07 $X=28403 $Y=50503 $D=636
M2484 754 vdd vdd vdd hvtpfet l=6e-08 w=6e-07 $X=28410 $Y=18290 $D=636
M2485 vdd vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=28410 $Y=35893 $D=636
M2486 755 vdd vdd vdd hvtpfet l=6e-08 w=8e-07 $X=28453 $Y=27288 $D=636
M2487 vdd vdd vdd vdd hvtpfet l=6e-08 w=6e-07 $X=28463 $Y=29008 $D=636
M2488 vdd vdd vdd vdd hvtpfet l=1e-07 w=6e-07 $X=28600 $Y=32628 $D=636
M2489 vdd vdd 752 vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=28615 $Y=15090 $D=636
M2490 vdd vdd 753 vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=28615 $Y=16110 $D=636
M2491 vdd vdd 754 vdd hvtpfet l=6e-08 w=6e-07 $X=28670 $Y=18290 $D=636
M2492 vdd vdd 755 vdd hvtpfet l=6e-08 w=8e-07 $X=28713 $Y=27288 $D=636
M2493 vdd vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=28750 $Y=35893 $D=636
M2494 b_bla<0> 285 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=28837 $Y=-170 $D=636
M2495 t_bla<0> 286 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=28837 $Y=50503 $D=636
M2496 325 283 b_bla<0> vdd hvtpfet l=6e-08 w=3e-07 $X=28860 $Y=1094 $D=636
M2497 b_bla<0> 283 325 vdd hvtpfet l=6e-08 w=3e-07 $X=28860 $Y=1354 $D=636
M2498 b_bla_n<0> 283 326 vdd hvtpfet l=6e-08 w=3e-07 $X=28860 $Y=1864 $D=636
M2499 326 283 b_bla_n<0> vdd hvtpfet l=6e-08 w=3e-07 $X=28860 $Y=2124 $D=636
M2500 t_bla_n<0> 284 326 vdd hvtpfet l=6e-08 w=3e-07 $X=28860 $Y=48949 $D=636
M2501 326 284 t_bla_n<0> vdd hvtpfet l=6e-08 w=3e-07 $X=28860 $Y=49209 $D=636
M2502 325 284 t_bla<0> vdd hvtpfet l=6e-08 w=3e-07 $X=28860 $Y=49719 $D=636
M2503 t_bla<0> 284 325 vdd hvtpfet l=6e-08 w=3e-07 $X=28860 $Y=49979 $D=636
M2504 vdd vdd vdd vdd hvtpfet l=1e-07 w=2e-07 $X=28875 $Y=36723 $D=636
M2505 vdd vdd vdd vdd hvtpfet l=1e-07 w=6e-07 $X=28900 $Y=32628 $D=636
M2506 vdd vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=29090 $Y=35893 $D=636
M2507 b_bla_n<0> 285 b_bla<0> vdd hvtpfet l=6e-08 w=8e-07 $X=29097 $Y=-170 $D=636
M2508 t_bla_n<0> 286 t_bla<0> vdd hvtpfet l=6e-08 w=8e-07 $X=29097 $Y=50503 $D=636
M2509 vdd vdd vdd vdd hvtpfet l=1e-07 w=2e-07 $X=29175 $Y=36723 $D=636
M2510 778 vdd vdd vdd hvtpfet l=6e-08 w=5e-07 $X=29180 $Y=18290 $D=636
M2511 1301 283 287 vdd hvtpfet l=6e-08 w=8e-07 $X=29185 $Y=5556 $D=636
M2512 283 b_ca<0> vdd vdd hvtpfet l=6e-08 w=4e-07 $X=29185 $Y=10611 $D=636
M2513 285 283 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=29185 $Y=12911 $D=636
M2514 286 284 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=29185 $Y=37822 $D=636
M2515 284 t_ca<0> vdd vdd hvtpfet l=6e-08 w=4e-07 $X=29185 $Y=40122 $D=636
M2516 1302 284 288 vdd hvtpfet l=6e-08 w=8e-07 $X=29185 $Y=44777 $D=636
M2517 vdd vdd vdd vdd hvtpfet l=7e-08 w=3.2e-07 $X=29210 $Y=32628 $D=636
M2518 767 vdd vdd vdd hvtpfet l=6e-08 w=6e-07 $X=29233 $Y=27488 $D=636
M2519 vdd 285 b_bla_n<0> vdd hvtpfet l=6e-08 w=8e-07 $X=29357 $Y=-170 $D=636
M2520 vdd 286 t_bla_n<0> vdd hvtpfet l=6e-08 w=8e-07 $X=29357 $Y=50503 $D=636
M2521 vdd vdd vdd vdd hvtpfet l=6e-08 w=6e-07 $X=29373 $Y=29008 $D=636
M2522 vdd vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=29430 $Y=35893 $D=636
M2523 vdd vdd 778 vdd hvtpfet l=6e-08 w=5e-07 $X=29440 $Y=18290 $D=636
M2524 vdd 20 1301 vdd hvtpfet l=6e-08 w=8e-07 $X=29445 $Y=5556 $D=636
M2525 vdd b_ma<0> 283 vdd hvtpfet l=6e-08 w=4e-07 $X=29445 $Y=10611 $D=636
M2526 vdd 22 285 vdd hvtpfet l=6e-08 w=4e-07 $X=29445 $Y=12911 $D=636
M2527 vdd 23 286 vdd hvtpfet l=6e-08 w=4e-07 $X=29445 $Y=37822 $D=636
M2528 vdd t_ma<0> 284 vdd hvtpfet l=6e-08 w=4e-07 $X=29445 $Y=40122 $D=636
M2529 vdd 20 1302 vdd hvtpfet l=6e-08 w=8e-07 $X=29445 $Y=44777 $D=636
M2530 vdd vdd vdd vdd hvtpfet l=1e-07 w=2e-07 $X=29475 $Y=36723 $D=636
M2531 vdd vdd vdd vdd hvtpfet l=7e-08 w=3.2e-07 $X=29500 $Y=32628 $D=636
M2532 vdd vdd vdd vdd hvtpfet l=6e-08 w=6e-07 $X=29633 $Y=29008 $D=636
M2533 778 vdd vdd vdd hvtpfet l=6e-08 w=5e-07 $X=29700 $Y=18290 $D=636
M2534 1303 11 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=29705 $Y=5556 $D=636
M2535 289 b_mb<0> vdd vdd hvtpfet l=6e-08 w=4e-07 $X=29705 $Y=10611 $D=636
M2536 293 13 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=29705 $Y=12911 $D=636
M2537 294 14 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=29705 $Y=37822 $D=636
M2538 290 t_mb<0> vdd vdd hvtpfet l=6e-08 w=4e-07 $X=29705 $Y=40122 $D=636
M2539 1304 11 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=29705 $Y=44777 $D=636
M2540 vdd vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=29770 $Y=35893 $D=636
M2541 vdd vdd vdd vdd hvtpfet l=1e-07 w=2e-07 $X=29775 $Y=36723 $D=636
M2542 b_blb<0> 293 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=29793 $Y=-170 $D=636
M2543 t_blb<0> 294 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=29793 $Y=50503 $D=636
M2544 768 vdd vdd vdd hvtpfet l=6e-08 w=4e-07 $X=29905 $Y=21427 $D=636
M2545 769 vdd vdd vdd hvtpfet l=6e-08 w=4e-07 $X=29905 $Y=23694 $D=636
M2546 770 vdd vdd vdd hvtpfet l=6e-08 w=4e-07 $X=29905 $Y=24394 $D=636
M2547 771 vdd vdd vdd hvtpfet l=6e-08 w=4e-07 $X=29905 $Y=24904 $D=636
M2548 vdd vdd 778 vdd hvtpfet l=6e-08 w=5e-07 $X=29960 $Y=18290 $D=636
M2549 291 289 1303 vdd hvtpfet l=6e-08 w=8e-07 $X=29965 $Y=5556 $D=636
M2550 vdd b_cb<0> 289 vdd hvtpfet l=6e-08 w=4e-07 $X=29965 $Y=10611 $D=636
M2551 vdd 289 293 vdd hvtpfet l=6e-08 w=4e-07 $X=29965 $Y=12911 $D=636
M2552 vdd 290 294 vdd hvtpfet l=6e-08 w=4e-07 $X=29965 $Y=37822 $D=636
M2553 vdd t_cb<0> 290 vdd hvtpfet l=6e-08 w=4e-07 $X=29965 $Y=40122 $D=636
M2554 292 290 1304 vdd hvtpfet l=6e-08 w=8e-07 $X=29965 $Y=44777 $D=636
M2555 296 289 b_blb<0> vdd hvtpfet l=6e-08 w=3e-07 $X=30050 $Y=1094 $D=636
M2556 b_blb<0> 289 296 vdd hvtpfet l=6e-08 w=3e-07 $X=30050 $Y=1354 $D=636
M2557 b_blb_n<0> 289 297 vdd hvtpfet l=6e-08 w=3e-07 $X=30050 $Y=1864 $D=636
M2558 297 289 b_blb_n<0> vdd hvtpfet l=6e-08 w=3e-07 $X=30050 $Y=2124 $D=636
M2559 t_blb_n<0> 290 297 vdd hvtpfet l=6e-08 w=3e-07 $X=30050 $Y=48949 $D=636
M2560 297 290 t_blb_n<0> vdd hvtpfet l=6e-08 w=3e-07 $X=30050 $Y=49209 $D=636
M2561 296 290 t_blb<0> vdd hvtpfet l=6e-08 w=3e-07 $X=30050 $Y=49719 $D=636
M2562 t_blb<0> 290 296 vdd hvtpfet l=6e-08 w=3e-07 $X=30050 $Y=49979 $D=636
M2563 b_blb_n<0> 293 b_blb<0> vdd hvtpfet l=6e-08 w=8e-07 $X=30053 $Y=-170 $D=636
M2564 t_blb_n<0> 294 t_blb<0> vdd hvtpfet l=6e-08 w=8e-07 $X=30053 $Y=50503 $D=636
M2565 vdd vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=30215 $Y=35893 $D=636
M2566 vdd 293 b_blb_n<0> vdd hvtpfet l=6e-08 w=8e-07 $X=30313 $Y=-170 $D=636
M2567 vdd 294 t_blb_n<0> vdd hvtpfet l=6e-08 w=8e-07 $X=30313 $Y=50503 $D=636
.ends

************************************************************************
* Library Name: XMC55_DPS
* Cell Name:    xmc55_dps_localc16io_dummy
************************************************************************
.SUBCKT xmc55_dps_localc16io_dummy b_dbl b_dwl b_tie_low dbl_pd_n<3> 
+ dbl_pd_n<2> dbl_pd_n<1> dbl_pd_n<0> stclk t_dbl t_dwl t_tie_low vdd vss
** N=889 EP=13 IP=0 FDC=76
M0 vss 2 17 vss hvtnfet l=6e-08 w=2e-07 $X=265 $Y=2781 $D=616
M1 vss 3 18 vss hvtnfet l=6e-08 w=2e-07 $X=265 $Y=48152 $D=616
M2 28 t_dbl vss vss hvtnfet l=6e-08 w=4e-07 $X=340 $Y=26568 $D=616
M3 vss 8 stclk vss hvtnfet l=6e-08 w=3e-07 $X=340 $Y=29928 $D=616
M4 49 b_dwl vss vss hvtnfet l=6e-08 w=4e-07 $X=535 $Y=2781 $D=616
M5 50 t_dwl vss vss hvtnfet l=6e-08 w=4e-07 $X=535 $Y=47952 $D=616
M6 b_tie_low 15 vss vss hvtnfet l=7e-08 w=3.2e-07 $X=540 $Y=4916 $D=616
M7 t_tie_low 16 vss vss hvtnfet l=7e-08 w=3.2e-07 $X=540 $Y=45897 $D=616
M8 8 b_dbl 28 vss hvtnfet l=6e-08 w=4e-07 $X=600 $Y=26568 $D=616
M9 vss dbl_pd_n<2> 12 vss hvtnfet l=6e-08 w=3e-07 $X=630 $Y=19039 $D=616
M10 vss dbl_pd_n<1> 14 vss hvtnfet l=6e-08 w=3e-07 $X=630 $Y=21399 $D=616
M11 vss dbl_pd_n<0> 13 vss hvtnfet l=6e-08 w=3e-07 $X=630 $Y=22329 $D=616
M12 vss dbl_pd_n<3> 21 vss hvtnfet l=6e-08 w=3e-07 $X=630 $Y=24794 $D=616
M13 2 21 49 vss hvtnfet l=6e-08 w=4e-07 $X=795 $Y=2781 $D=616
M14 3 21 50 vss hvtnfet l=6e-08 w=4e-07 $X=795 $Y=47952 $D=616
M15 vdd vdd vdd vdd hvtpfet l=6e-08 w=8e-07 $X=187 $Y=-170 $D=636
M16 vdd vdd vdd vdd hvtpfet l=6e-08 w=8e-07 $X=187 $Y=50503 $D=636
M17 vdd 2 17 vdd hvtpfet l=6e-08 w=4e-07 $X=265 $Y=2061 $D=636
M18 vdd 3 18 vdd hvtpfet l=6e-08 w=4e-07 $X=265 $Y=48672 $D=636
M19 8 t_dbl vdd vdd hvtpfet l=6e-08 w=4e-07 $X=340 $Y=27288 $D=636
M20 vdd 8 stclk vdd hvtpfet l=6e-08 w=6e-07 $X=340 $Y=29008 $D=636
M21 b_dbl vdd vdd vdd hvtpfet l=6e-08 w=8e-07 $X=447 $Y=-170 $D=636
M22 t_dbl vdd vdd vdd hvtpfet l=6e-08 w=8e-07 $X=447 $Y=50503 $D=636
M23 2 b_dwl vdd vdd hvtpfet l=6e-08 w=4e-07 $X=535 $Y=2061 $D=636
M24 3 t_dwl vdd vdd hvtpfet l=6e-08 w=4e-07 $X=535 $Y=48672 $D=636
M25 15 15 vdd vdd hvtpfet l=7e-08 w=6.4e-07 $X=540 $Y=5556 $D=636
M26 16 16 vdd vdd hvtpfet l=7e-08 w=6.4e-07 $X=540 $Y=44937 $D=636
M27 vdd b_dbl 8 vdd hvtpfet l=6e-08 w=4e-07 $X=600 $Y=27288 $D=636
M28 vdd dbl_pd_n<2> 12 vdd hvtpfet l=6e-08 w=5e-07 $X=630 $Y=19659 $D=636
M29 vdd dbl_pd_n<1> 14 vdd hvtpfet l=6e-08 w=5e-07 $X=630 $Y=20579 $D=636
M30 vdd dbl_pd_n<0> 13 vdd hvtpfet l=6e-08 w=5e-07 $X=630 $Y=22949 $D=636
M31 vdd dbl_pd_n<3> 21 vdd hvtpfet l=6e-08 w=5e-07 $X=630 $Y=23974 $D=636
M32 vdd b_dwl b_dbl vdd hvtpfet l=6e-08 w=8e-07 $X=707 $Y=-170 $D=636
M33 vdd t_dwl t_dbl vdd hvtpfet l=6e-08 w=8e-07 $X=707 $Y=50503 $D=636
M34 vdd 21 2 vdd hvtpfet l=6e-08 w=4e-07 $X=795 $Y=2061 $D=636
M35 vdd 21 3 vdd hvtpfet l=6e-08 w=4e-07 $X=795 $Y=48672 $D=636
M36 vss t_tie_low 29 vss srpddnfet l=6e-08 w=3.15e-07 $X=670 $Y=7281 $D=778
M37 vss t_tie_low 30 vss srpddnfet l=6e-08 w=3.15e-07 $X=670 $Y=7876 $D=778
M38 vss t_tie_low 31 vss srpddnfet l=6e-08 w=3.15e-07 $X=670 $Y=9246 $D=778
M39 vss 12 32 vss srpddnfet l=6e-08 w=3.15e-07 $X=670 $Y=10871 $D=778
M40 vss 12 33 vss srpddnfet l=6e-08 w=3.15e-07 $X=670 $Y=11466 $D=778
M41 vss 12 34 vss srpddnfet l=6e-08 w=3.15e-07 $X=670 $Y=13091 $D=778
M42 vss 12 35 vss srpddnfet l=6e-08 w=3.15e-07 $X=670 $Y=13686 $D=778
M43 vss 13 36 vss srpddnfet l=6e-08 w=3.15e-07 $X=670 $Y=15311 $D=778
M44 vss 14 37 vss srpddnfet l=6e-08 w=3.15e-07 $X=670 $Y=16681 $D=778
M45 vss 14 38 vss srpddnfet l=6e-08 w=3.15e-07 $X=670 $Y=17276 $D=778
M46 vss 14 39 vss srpddnfet l=6e-08 w=3.15e-07 $X=670 $Y=33542 $D=778
M47 vss 14 40 vss srpddnfet l=6e-08 w=3.15e-07 $X=670 $Y=34137 $D=778
M48 vss 13 41 vss srpddnfet l=6e-08 w=3.15e-07 $X=670 $Y=35507 $D=778
M49 vss 12 42 vss srpddnfet l=6e-08 w=3.15e-07 $X=670 $Y=37132 $D=778
M50 vss 12 43 vss srpddnfet l=6e-08 w=3.15e-07 $X=670 $Y=37727 $D=778
M51 vss 12 44 vss srpddnfet l=6e-08 w=3.15e-07 $X=670 $Y=39352 $D=778
M52 vss 12 45 vss srpddnfet l=6e-08 w=3.15e-07 $X=670 $Y=39947 $D=778
M53 vss t_tie_low 46 vss srpddnfet l=6e-08 w=3.15e-07 $X=670 $Y=41572 $D=778
M54 vss t_tie_low 47 vss srpddnfet l=6e-08 w=3.15e-07 $X=670 $Y=42942 $D=778
M55 vss t_tie_low 48 vss srpddnfet l=6e-08 w=3.15e-07 $X=670 $Y=43537 $D=778
M56 b_dbl 17 29 vss srpgdnfet l=7.5e-08 w=1.05e-07 $X=655 $Y=6816 $D=780
M57 b_dbl 17 30 vss srpgdnfet l=7.5e-08 w=1.05e-07 $X=655 $Y=8551 $D=780
M58 b_dbl 17 31 vss srpgdnfet l=7.5e-08 w=1.05e-07 $X=655 $Y=9921 $D=780
M59 b_dbl 17 32 vss srpgdnfet l=7.5e-08 w=1.05e-07 $X=655 $Y=10406 $D=780
M60 b_dbl 17 33 vss srpgdnfet l=7.5e-08 w=1.05e-07 $X=655 $Y=12141 $D=780
M61 b_dbl 17 34 vss srpgdnfet l=7.5e-08 w=1.05e-07 $X=655 $Y=12626 $D=780
M62 b_dbl 17 35 vss srpgdnfet l=7.5e-08 w=1.05e-07 $X=655 $Y=14361 $D=780
M63 b_dbl 17 36 vss srpgdnfet l=7.5e-08 w=1.05e-07 $X=655 $Y=14846 $D=780
M64 b_dbl 17 37 vss srpgdnfet l=7.5e-08 w=1.05e-07 $X=655 $Y=16216 $D=780
M65 b_dbl 17 38 vss srpgdnfet l=7.5e-08 w=1.05e-07 $X=655 $Y=17951 $D=780
M66 t_dbl 18 39 vss srpgdnfet l=7.5e-08 w=1.05e-07 $X=655 $Y=33077 $D=780
M67 t_dbl 18 40 vss srpgdnfet l=7.5e-08 w=1.05e-07 $X=655 $Y=34812 $D=780
M68 t_dbl 18 41 vss srpgdnfet l=7.5e-08 w=1.05e-07 $X=655 $Y=36182 $D=780
M69 t_dbl 18 42 vss srpgdnfet l=7.5e-08 w=1.05e-07 $X=655 $Y=36667 $D=780
M70 t_dbl 18 43 vss srpgdnfet l=7.5e-08 w=1.05e-07 $X=655 $Y=38402 $D=780
M71 t_dbl 18 44 vss srpgdnfet l=7.5e-08 w=1.05e-07 $X=655 $Y=38887 $D=780
M72 t_dbl 18 45 vss srpgdnfet l=7.5e-08 w=1.05e-07 $X=655 $Y=40622 $D=780
M73 t_dbl 18 46 vss srpgdnfet l=7.5e-08 w=1.05e-07 $X=655 $Y=41107 $D=780
M74 t_dbl 18 47 vss srpgdnfet l=7.5e-08 w=1.05e-07 $X=655 $Y=42477 $D=780
M75 t_dbl 18 48 vss srpgdnfet l=7.5e-08 w=1.05e-07 $X=655 $Y=44212 $D=780
.ends

************************************************************************
* Library Name: XMC55_DPS
* Cell Name:    xmc55_dps_localc16io_edge
************************************************************************
.SUBCKT xmc55_dps_localc16io_edge tie_low vdd vss
** N=1093 EP=3 IP=0 FDC=59
M0 vss vss vss vss hvtnfet l=6e-08 w=4e-07 $X=970 $Y=2941 $D=616
M1 vss vss vss vss hvtnfet l=6e-08 w=4e-07 $X=970 $Y=3201 $D=616
M2 vss vss vss vss hvtnfet l=6e-08 w=4e-07 $X=970 $Y=3881 $D=616
M3 vss vss vss vss hvtnfet l=6e-08 w=4e-07 $X=970 $Y=4141 $D=616
M4 vss vss vss vss hvtnfet l=6e-08 w=4e-07 $X=970 $Y=46932 $D=616
M5 vss vss vss vss hvtnfet l=6e-08 w=4e-07 $X=970 $Y=47192 $D=616
M6 vss vss vss vss hvtnfet l=6e-08 w=4e-07 $X=970 $Y=47872 $D=616
M7 vss vss vss vss hvtnfet l=6e-08 w=4e-07 $X=970 $Y=48132 $D=616
M8 18 tie_low vss vss hvtnfet l=6e-08 w=2.1e-07 $X=1025 $Y=14555 $D=616
M9 19 tie_low vss vss hvtnfet l=6e-08 w=2.1e-07 $X=1025 $Y=16755 $D=616
M10 20 tie_low vss vss hvtnfet l=6e-08 w=2.1e-07 $X=1025 $Y=17760 $D=616
M11 5 5 vss vss hvtnfet l=6e-08 w=3.2e-07 $X=1025 $Y=26624 $D=616
M12 vss 2 tie_low vss hvtnfet l=6e-08 w=2.1e-07 $X=1025 $Y=33548 $D=616
M13 vss tie_low 10 vss hvtnfet l=6e-08 w=4e-07 $X=1130 $Y=4836 $D=616
M14 vss tie_low 11 vss hvtnfet l=6e-08 w=4e-07 $X=1130 $Y=11331 $D=616
M15 vss tie_low 12 vss hvtnfet l=6e-08 w=4e-07 $X=1130 $Y=12191 $D=616
M16 vss tie_low 13 vss hvtnfet l=6e-08 w=4e-07 $X=1130 $Y=38542 $D=616
M17 vss tie_low 14 vss hvtnfet l=6e-08 w=4e-07 $X=1130 $Y=39402 $D=616
M18 vss tie_low 15 vss hvtnfet l=6e-08 w=4e-07 $X=1130 $Y=45897 $D=616
M19 vss 5 5 vss hvtnfet l=6e-08 w=3.2e-07 $X=1285 $Y=26624 $D=616
M20 vdd vdd vdd vdd hvtpfet l=6e-08 w=3e-07 $X=975 $Y=19812 $D=636
M21 vdd vdd vdd vdd hvtpfet l=6e-08 w=3e-07 $X=975 $Y=20072 $D=636
M22 vdd vdd vdd vdd hvtpfet l=6e-08 w=3e-07 $X=975 $Y=20902 $D=636
M23 vdd vdd vdd vdd hvtpfet l=6e-08 w=3e-07 $X=975 $Y=21162 $D=636
M24 vdd vdd vdd vdd hvtpfet l=6e-08 w=3e-07 $X=975 $Y=21422 $D=636
M25 vdd vdd vdd vdd hvtpfet l=6e-08 w=3e-07 $X=975 $Y=21682 $D=636
M26 vdd vdd vdd vdd hvtpfet l=6e-08 w=3e-07 $X=975 $Y=21942 $D=636
M27 vdd vdd vdd vdd hvtpfet l=6e-08 w=3e-07 $X=975 $Y=22762 $D=636
M28 vdd vdd vdd vdd hvtpfet l=6e-08 w=3e-07 $X=975 $Y=23729 $D=636
M29 vdd vdd vdd vdd hvtpfet l=6e-08 w=3e-07 $X=975 $Y=23989 $D=636
M30 vdd vdd vdd vdd hvtpfet l=6e-08 w=3e-07 $X=975 $Y=24249 $D=636
M31 vdd vdd vdd vdd hvtpfet l=6e-08 w=3e-07 $X=975 $Y=24509 $D=636
M32 vdd vdd vdd vdd hvtpfet l=6e-08 w=3e-07 $X=975 $Y=24769 $D=636
M33 18 tie_low vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=1025 $Y=15085 $D=636
M34 19 tie_low vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=1025 $Y=16115 $D=636
M35 20 tie_low vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=1025 $Y=18290 $D=636
M36 21 5 2 vdd hvtpfet l=6e-08 w=4.8e-07 $X=1025 $Y=27313 $D=636
M37 22 5 2 vdd hvtpfet l=6e-08 w=4.8e-07 $X=1025 $Y=29008 $D=636
M38 vdd 2 tie_low vdd hvtpfet l=6e-08 w=3.2e-07 $X=1025 $Y=32908 $D=636
M39 vdd vdd vdd vdd hvtpfet l=6e-08 w=3e-07 $X=1070 $Y=1094 $D=636
M40 vdd vdd vdd vdd hvtpfet l=6e-08 w=3e-07 $X=1070 $Y=1354 $D=636
M41 vdd vdd vdd vdd hvtpfet l=6e-08 w=3e-07 $X=1070 $Y=1864 $D=636
M42 vdd vdd vdd vdd hvtpfet l=6e-08 w=3e-07 $X=1070 $Y=2124 $D=636
M43 vdd vdd vdd vdd hvtpfet l=6e-08 w=3e-07 $X=1070 $Y=48949 $D=636
M44 vdd vdd vdd vdd hvtpfet l=6e-08 w=3e-07 $X=1070 $Y=49209 $D=636
M45 vdd vdd vdd vdd hvtpfet l=6e-08 w=3e-07 $X=1070 $Y=49719 $D=636
M46 vdd vdd vdd vdd hvtpfet l=6e-08 w=3e-07 $X=1070 $Y=49979 $D=636
M47 vdd vdd vdd vdd hvtpfet l=6e-08 w=8e-07 $X=1073 $Y=-170 $D=636
M48 vdd vdd vdd vdd hvtpfet l=6e-08 w=8e-07 $X=1073 $Y=50503 $D=636
M49 vdd tie_low 10 vdd hvtpfet l=6e-08 w=8e-07 $X=1130 $Y=5556 $D=636
M50 vdd tie_low 11 vdd hvtpfet l=6e-08 w=4e-07 $X=1130 $Y=10611 $D=636
M51 vdd tie_low 12 vdd hvtpfet l=6e-08 w=4e-07 $X=1130 $Y=12911 $D=636
M52 vdd tie_low 13 vdd hvtpfet l=6e-08 w=4e-07 $X=1130 $Y=37822 $D=636
M53 vdd tie_low 14 vdd hvtpfet l=6e-08 w=4e-07 $X=1130 $Y=40122 $D=636
M54 vdd tie_low 15 vdd hvtpfet l=6e-08 w=8e-07 $X=1130 $Y=44777 $D=636
M55 vdd 5 21 vdd hvtpfet l=6e-08 w=4.8e-07 $X=1285 $Y=27313 $D=636
M56 vdd 5 22 vdd hvtpfet l=6e-08 w=4.8e-07 $X=1285 $Y=29008 $D=636
M57 vdd vdd vdd vdd hvtpfet l=6e-08 w=8e-07 $X=1333 $Y=-170 $D=636
M58 vdd vdd vdd vdd hvtpfet l=6e-08 w=8e-07 $X=1333 $Y=50503 $D=636
.ends

************************************************************************
* Library Name: XMC55_DPS
* Cell Name:    xmc55_dps_collar_dq_16_bw
************************************************************************
.SUBCKT xmc55_dps_collar_dq_16_bw bwena bwena_int bwenb bwenb_int da da_int db 
+ db_int qa qa_int qb qb_int vdd vss
** N=1201 EP=14 IP=0 FDC=148
D0 vss bwena diodenx AREA=7.04e-14 $X=11827 $Y=130 $D=2
D1 vss da diodenx AREA=7.04e-14 $X=13732 $Y=130 $D=2
D2 vss db diodenx AREA=7.04e-14 $X=15650 $Y=130 $D=2
D3 vss bwenb diodenx AREA=7.04e-14 $X=17555 $Y=130 $D=2
M4 12 vdd vss vss hvtnfet l=6e-08 w=6e-07 $X=580 $Y=1420 $D=616
M5 13 vdd vss vss hvtnfet l=6e-08 w=9e-07 $X=1090 $Y=1120 $D=616
M6 vss vdd 13 vss hvtnfet l=6e-08 w=9e-07 $X=1350 $Y=1120 $D=616
M7 14 vdd vss vss hvtnfet l=6e-08 w=9e-07 $X=1610 $Y=1120 $D=616
M8 vss vdd 14 vss hvtnfet l=6e-08 w=9e-07 $X=1870 $Y=1120 $D=616
M9 vss vdd 15 vss hvtnfet l=6e-08 w=6e-07 $X=2380 $Y=1420 $D=616
M10 16 vdd vss vss hvtnfet l=6e-08 w=6e-07 $X=2890 $Y=1420 $D=616
M11 17 vdd vss vss hvtnfet l=6e-08 w=9e-07 $X=3400 $Y=1120 $D=616
M12 vss vdd 17 vss hvtnfet l=6e-08 w=9e-07 $X=3660 $Y=1120 $D=616
M13 18 vdd vss vss hvtnfet l=6e-08 w=6e-07 $X=4400 $Y=1420 $D=616
M14 19 vdd vss vss hvtnfet l=6e-08 w=9e-07 $X=4910 $Y=1120 $D=616
M15 vss vdd 19 vss hvtnfet l=6e-08 w=9e-07 $X=5170 $Y=1120 $D=616
M16 20 vdd vss vss hvtnfet l=6e-08 w=9e-07 $X=5430 $Y=1120 $D=616
M17 vss vdd 20 vss hvtnfet l=6e-08 w=9e-07 $X=5690 $Y=1120 $D=616
M18 vss vdd 21 vss hvtnfet l=6e-08 w=6e-07 $X=6200 $Y=1420 $D=616
M19 22 vdd vss vss hvtnfet l=6e-08 w=6e-07 $X=6710 $Y=1420 $D=616
M20 23 vdd vss vss hvtnfet l=6e-08 w=9e-07 $X=7220 $Y=1120 $D=616
M21 vss vdd 23 vss hvtnfet l=6e-08 w=9e-07 $X=7480 $Y=1120 $D=616
M22 24 vdd vss vss hvtnfet l=6e-08 w=6e-07 $X=8220 $Y=1420 $D=616
M23 25 vdd vss vss hvtnfet l=6e-08 w=9e-07 $X=8730 $Y=1120 $D=616
M24 vss vdd 25 vss hvtnfet l=6e-08 w=9e-07 $X=8990 $Y=1120 $D=616
M25 26 vdd vss vss hvtnfet l=6e-08 w=9e-07 $X=9250 $Y=1120 $D=616
M26 vss vdd 26 vss hvtnfet l=6e-08 w=9e-07 $X=9510 $Y=1120 $D=616
M27 vss vdd 27 vss hvtnfet l=6e-08 w=6e-07 $X=10020 $Y=1420 $D=616
M28 28 vdd vss vss hvtnfet l=6e-08 w=6e-07 $X=10530 $Y=1420 $D=616
M29 29 vdd vss vss hvtnfet l=6e-08 w=9e-07 $X=11040 $Y=1120 $D=616
M30 vss vdd 29 vss hvtnfet l=6e-08 w=9e-07 $X=11300 $Y=1120 $D=616
M31 3 bwena vss vss hvtnfet l=6e-08 w=6e-07 $X=12040 $Y=1420 $D=616
M32 bwena_int 3 vss vss hvtnfet l=6e-08 w=9e-07 $X=12550 $Y=1120 $D=616
M33 vss 3 bwena_int vss hvtnfet l=6e-08 w=9e-07 $X=12810 $Y=1120 $D=616
M34 qa qa_int vss vss hvtnfet l=6e-08 w=9e-07 $X=13070 $Y=1120 $D=616
M35 vss qa_int qa vss hvtnfet l=6e-08 w=9e-07 $X=13330 $Y=1120 $D=616
M36 vss vdd 32 vss hvtnfet l=6e-08 w=6e-07 $X=13840 $Y=1420 $D=616
M37 6 da vss vss hvtnfet l=6e-08 w=6e-07 $X=14350 $Y=1420 $D=616
M38 da_int 6 vss vss hvtnfet l=6e-08 w=9e-07 $X=14860 $Y=1120 $D=616
M39 vss 6 da_int vss hvtnfet l=6e-08 w=9e-07 $X=15120 $Y=1120 $D=616
M40 db_int 7 vss vss hvtnfet l=6e-08 w=9e-07 $X=15380 $Y=1120 $D=616
M41 vss 7 db_int vss hvtnfet l=6e-08 w=9e-07 $X=15640 $Y=1120 $D=616
M42 vss db 7 vss hvtnfet l=6e-08 w=6e-07 $X=16150 $Y=1420 $D=616
M43 36 vdd vss vss hvtnfet l=6e-08 w=6e-07 $X=16660 $Y=1420 $D=616
M44 qb qb_int vss vss hvtnfet l=6e-08 w=9e-07 $X=17170 $Y=1120 $D=616
M45 vss qb_int qb vss hvtnfet l=6e-08 w=9e-07 $X=17430 $Y=1120 $D=616
M46 bwenb_int 10 vss vss hvtnfet l=6e-08 w=9e-07 $X=17690 $Y=1120 $D=616
M47 vss 10 bwenb_int vss hvtnfet l=6e-08 w=9e-07 $X=17950 $Y=1120 $D=616
M48 vss bwenb 10 vss hvtnfet l=6e-08 w=6e-07 $X=18460 $Y=1420 $D=616
M49 38 vdd vss vss hvtnfet l=6e-08 w=9e-07 $X=19200 $Y=1120 $D=616
M50 vss vdd 38 vss hvtnfet l=6e-08 w=9e-07 $X=19460 $Y=1120 $D=616
M51 vss vdd 39 vss hvtnfet l=6e-08 w=6e-07 $X=19970 $Y=1420 $D=616
M52 40 vdd vss vss hvtnfet l=6e-08 w=6e-07 $X=20480 $Y=1420 $D=616
M53 41 vdd vss vss hvtnfet l=6e-08 w=9e-07 $X=20990 $Y=1120 $D=616
M54 vss vdd 41 vss hvtnfet l=6e-08 w=9e-07 $X=21250 $Y=1120 $D=616
M55 42 vdd vss vss hvtnfet l=6e-08 w=9e-07 $X=21510 $Y=1120 $D=616
M56 vss vdd 42 vss hvtnfet l=6e-08 w=9e-07 $X=21770 $Y=1120 $D=616
M57 vss vdd 43 vss hvtnfet l=6e-08 w=6e-07 $X=22280 $Y=1420 $D=616
M58 44 vdd vss vss hvtnfet l=6e-08 w=9e-07 $X=23020 $Y=1120 $D=616
M59 vss vdd 44 vss hvtnfet l=6e-08 w=9e-07 $X=23280 $Y=1120 $D=616
M60 vss vdd 45 vss hvtnfet l=6e-08 w=6e-07 $X=23790 $Y=1420 $D=616
M61 46 vdd vss vss hvtnfet l=6e-08 w=6e-07 $X=24300 $Y=1420 $D=616
M62 47 vdd vss vss hvtnfet l=6e-08 w=9e-07 $X=24810 $Y=1120 $D=616
M63 vss vdd 47 vss hvtnfet l=6e-08 w=9e-07 $X=25070 $Y=1120 $D=616
M64 48 vdd vss vss hvtnfet l=6e-08 w=9e-07 $X=25330 $Y=1120 $D=616
M65 vss vdd 48 vss hvtnfet l=6e-08 w=9e-07 $X=25590 $Y=1120 $D=616
M66 vss vdd 49 vss hvtnfet l=6e-08 w=6e-07 $X=26100 $Y=1420 $D=616
M67 50 vdd vss vss hvtnfet l=6e-08 w=9e-07 $X=26840 $Y=1120 $D=616
M68 vss vdd 50 vss hvtnfet l=6e-08 w=9e-07 $X=27100 $Y=1120 $D=616
M69 vss vdd 51 vss hvtnfet l=6e-08 w=6e-07 $X=27610 $Y=1420 $D=616
M70 52 vdd vss vss hvtnfet l=6e-08 w=6e-07 $X=28120 $Y=1420 $D=616
M71 53 vdd vss vss hvtnfet l=6e-08 w=9e-07 $X=28630 $Y=1120 $D=616
M72 vss vdd 53 vss hvtnfet l=6e-08 w=9e-07 $X=28890 $Y=1120 $D=616
M73 54 vdd vss vss hvtnfet l=6e-08 w=9e-07 $X=29150 $Y=1120 $D=616
M74 vss vdd 54 vss hvtnfet l=6e-08 w=9e-07 $X=29410 $Y=1120 $D=616
M75 vss vdd 55 vss hvtnfet l=6e-08 w=6e-07 $X=29920 $Y=1420 $D=616
M76 12 vdd vdd vdd hvtpfet l=6e-08 w=1.2e-06 $X=580 $Y=2685 $D=636
M77 13 vdd vdd vdd hvtpfet l=6e-08 w=1.8e-06 $X=1090 $Y=2340 $D=636
M78 vdd vdd 13 vdd hvtpfet l=6e-08 w=1.8e-06 $X=1350 $Y=2340 $D=636
M79 14 vdd vdd vdd hvtpfet l=6e-08 w=1.8e-06 $X=1610 $Y=2340 $D=636
M80 vdd vdd 14 vdd hvtpfet l=6e-08 w=1.8e-06 $X=1870 $Y=2340 $D=636
M81 vdd vdd 15 vdd hvtpfet l=6e-08 w=1.2e-06 $X=2380 $Y=2685 $D=636
M82 16 vdd vdd vdd hvtpfet l=6e-08 w=1.2e-06 $X=2890 $Y=2685 $D=636
M83 17 vdd vdd vdd hvtpfet l=6e-08 w=1.8e-06 $X=3400 $Y=2340 $D=636
M84 vdd vdd 17 vdd hvtpfet l=6e-08 w=1.8e-06 $X=3660 $Y=2340 $D=636
M85 18 vdd vdd vdd hvtpfet l=6e-08 w=1.2e-06 $X=4400 $Y=2685 $D=636
M86 19 vdd vdd vdd hvtpfet l=6e-08 w=1.8e-06 $X=4910 $Y=2340 $D=636
M87 vdd vdd 19 vdd hvtpfet l=6e-08 w=1.8e-06 $X=5170 $Y=2340 $D=636
M88 20 vdd vdd vdd hvtpfet l=6e-08 w=1.8e-06 $X=5430 $Y=2340 $D=636
M89 vdd vdd 20 vdd hvtpfet l=6e-08 w=1.8e-06 $X=5690 $Y=2340 $D=636
M90 vdd vdd 21 vdd hvtpfet l=6e-08 w=1.2e-06 $X=6200 $Y=2685 $D=636
M91 22 vdd vdd vdd hvtpfet l=6e-08 w=1.2e-06 $X=6710 $Y=2685 $D=636
M92 23 vdd vdd vdd hvtpfet l=6e-08 w=1.8e-06 $X=7220 $Y=2340 $D=636
M93 vdd vdd 23 vdd hvtpfet l=6e-08 w=1.8e-06 $X=7480 $Y=2340 $D=636
M94 24 vdd vdd vdd hvtpfet l=6e-08 w=1.2e-06 $X=8220 $Y=2685 $D=636
M95 25 vdd vdd vdd hvtpfet l=6e-08 w=1.8e-06 $X=8730 $Y=2340 $D=636
M96 vdd vdd 25 vdd hvtpfet l=6e-08 w=1.8e-06 $X=8990 $Y=2340 $D=636
M97 26 vdd vdd vdd hvtpfet l=6e-08 w=1.8e-06 $X=9250 $Y=2340 $D=636
M98 vdd vdd 26 vdd hvtpfet l=6e-08 w=1.8e-06 $X=9510 $Y=2340 $D=636
M99 vdd vdd 27 vdd hvtpfet l=6e-08 w=1.2e-06 $X=10020 $Y=2685 $D=636
M100 28 vdd vdd vdd hvtpfet l=6e-08 w=1.2e-06 $X=10530 $Y=2685 $D=636
M101 29 vdd vdd vdd hvtpfet l=6e-08 w=1.8e-06 $X=11040 $Y=2340 $D=636
M102 vdd vdd 29 vdd hvtpfet l=6e-08 w=1.8e-06 $X=11300 $Y=2340 $D=636
M103 3 bwena vdd vdd hvtpfet l=6e-08 w=1.2e-06 $X=12040 $Y=2685 $D=636
M104 bwena_int 3 vdd vdd hvtpfet l=6e-08 w=1.8e-06 $X=12550 $Y=2340 $D=636
M105 vdd 3 bwena_int vdd hvtpfet l=6e-08 w=1.8e-06 $X=12810 $Y=2340 $D=636
M106 qa qa_int vdd vdd hvtpfet l=6e-08 w=1.8e-06 $X=13070 $Y=2340 $D=636
M107 vdd qa_int qa vdd hvtpfet l=6e-08 w=1.8e-06 $X=13330 $Y=2340 $D=636
M108 vdd vdd 32 vdd hvtpfet l=6e-08 w=1.2e-06 $X=13840 $Y=2685 $D=636
M109 6 da vdd vdd hvtpfet l=6e-08 w=1.2e-06 $X=14350 $Y=2685 $D=636
M110 da_int 6 vdd vdd hvtpfet l=6e-08 w=1.8e-06 $X=14860 $Y=2340 $D=636
M111 vdd 6 da_int vdd hvtpfet l=6e-08 w=1.8e-06 $X=15120 $Y=2340 $D=636
M112 db_int 7 vdd vdd hvtpfet l=6e-08 w=1.8e-06 $X=15380 $Y=2340 $D=636
M113 vdd 7 db_int vdd hvtpfet l=6e-08 w=1.8e-06 $X=15640 $Y=2340 $D=636
M114 vdd db 7 vdd hvtpfet l=6e-08 w=1.2e-06 $X=16150 $Y=2685 $D=636
M115 36 vdd vdd vdd hvtpfet l=6e-08 w=1.2e-06 $X=16660 $Y=2685 $D=636
M116 qb qb_int vdd vdd hvtpfet l=6e-08 w=1.8e-06 $X=17170 $Y=2340 $D=636
M117 vdd qb_int qb vdd hvtpfet l=6e-08 w=1.8e-06 $X=17430 $Y=2340 $D=636
M118 bwenb_int 10 vdd vdd hvtpfet l=6e-08 w=1.8e-06 $X=17690 $Y=2340 $D=636
M119 vdd 10 bwenb_int vdd hvtpfet l=6e-08 w=1.8e-06 $X=17950 $Y=2340 $D=636
M120 vdd bwenb 10 vdd hvtpfet l=6e-08 w=1.2e-06 $X=18460 $Y=2685 $D=636
M121 38 vdd vdd vdd hvtpfet l=6e-08 w=1.8e-06 $X=19200 $Y=2340 $D=636
M122 vdd vdd 38 vdd hvtpfet l=6e-08 w=1.8e-06 $X=19460 $Y=2340 $D=636
M123 vdd vdd 39 vdd hvtpfet l=6e-08 w=1.2e-06 $X=19970 $Y=2685 $D=636
M124 40 vdd vdd vdd hvtpfet l=6e-08 w=1.2e-06 $X=20480 $Y=2685 $D=636
M125 41 vdd vdd vdd hvtpfet l=6e-08 w=1.8e-06 $X=20990 $Y=2340 $D=636
M126 vdd vdd 41 vdd hvtpfet l=6e-08 w=1.8e-06 $X=21250 $Y=2340 $D=636
M127 42 vdd vdd vdd hvtpfet l=6e-08 w=1.8e-06 $X=21510 $Y=2340 $D=636
M128 vdd vdd 42 vdd hvtpfet l=6e-08 w=1.8e-06 $X=21770 $Y=2340 $D=636
M129 vdd vdd 43 vdd hvtpfet l=6e-08 w=1.2e-06 $X=22280 $Y=2685 $D=636
M130 44 vdd vdd vdd hvtpfet l=6e-08 w=1.8e-06 $X=23020 $Y=2340 $D=636
M131 vdd vdd 44 vdd hvtpfet l=6e-08 w=1.8e-06 $X=23280 $Y=2340 $D=636
M132 vdd vdd 45 vdd hvtpfet l=6e-08 w=1.2e-06 $X=23790 $Y=2685 $D=636
M133 46 vdd vdd vdd hvtpfet l=6e-08 w=1.2e-06 $X=24300 $Y=2685 $D=636
M134 47 vdd vdd vdd hvtpfet l=6e-08 w=1.8e-06 $X=24810 $Y=2340 $D=636
M135 vdd vdd 47 vdd hvtpfet l=6e-08 w=1.8e-06 $X=25070 $Y=2340 $D=636
M136 48 vdd vdd vdd hvtpfet l=6e-08 w=1.8e-06 $X=25330 $Y=2340 $D=636
M137 vdd vdd 48 vdd hvtpfet l=6e-08 w=1.8e-06 $X=25590 $Y=2340 $D=636
M138 vdd vdd 49 vdd hvtpfet l=6e-08 w=1.2e-06 $X=26100 $Y=2685 $D=636
M139 50 vdd vdd vdd hvtpfet l=6e-08 w=1.8e-06 $X=26840 $Y=2340 $D=636
M140 vdd vdd 50 vdd hvtpfet l=6e-08 w=1.8e-06 $X=27100 $Y=2340 $D=636
M141 vdd vdd 51 vdd hvtpfet l=6e-08 w=1.2e-06 $X=27610 $Y=2685 $D=636
M142 52 vdd vdd vdd hvtpfet l=6e-08 w=1.2e-06 $X=28120 $Y=2685 $D=636
M143 53 vdd vdd vdd hvtpfet l=6e-08 w=1.8e-06 $X=28630 $Y=2340 $D=636
M144 vdd vdd 53 vdd hvtpfet l=6e-08 w=1.8e-06 $X=28890 $Y=2340 $D=636
M145 54 vdd vdd vdd hvtpfet l=6e-08 w=1.8e-06 $X=29150 $Y=2340 $D=636
M146 vdd vdd 54 vdd hvtpfet l=6e-08 w=1.8e-06 $X=29410 $Y=2340 $D=636
M147 vdd vdd 55 vdd hvtpfet l=6e-08 w=1.2e-06 $X=29920 $Y=2685 $D=636
.ends

************************************************************************
* Library Name: XMC55_DPS
* Cell Name:    xmc55_dps_local_ctrl8
************************************************************************
.SUBCKT xmc55_dps_local_ctrl8 aa<12> aa<11> aa<10> aa<9> aa<8> aa<7> aa<6> 
+ aa<5> aa<4> aa<3> aa<2> aa<1> aa<0> ab<12> ab<11> ab<10> ab<9> ab<8> ab<7> 
+ ab<6> ab<5> ab<4> ab<3> ab<2> ab<1> ab<0> b_pxaa<3> b_pxaa<2> b_pxaa<1> 
+ b_pxaa<0> b_pxab<3> b_pxab<2> b_pxab<1> b_pxab<0> b_pxba_n<7> b_pxba_n<6> 
+ b_pxba_n<5> b_pxba_n<4> b_pxba_n<3> b_pxba_n<2> b_pxba_n<1> b_pxba_n<0> 
+ b_pxbb_n<7> b_pxbb_n<6> b_pxbb_n<5> b_pxbb_n<4> b_pxbb_n<3> b_pxbb_n<2> 
+ b_pxbb_n<1> b_pxbb_n<0> b_pxca_n<7> b_pxca_n<6> b_pxca_n<5> b_pxca_n<4> 
+ b_pxca_n<3> b_pxca_n<2> b_pxca_n<1> b_pxca_n<0> b_pxcb_n<7> b_pxcb_n<6> 
+ b_pxcb_n<5> b_pxcb_n<4> b_pxcb_n<3> b_pxcb_n<2> b_pxcb_n<1> b_pxcb_n<0> cena 
+ cenb clka clkb dbl_pd_n<3> dbl_pd_n<2> dbl_pd_n<1> dbl_pd_n<0> ddqa ddqa_n 
+ ddqb ddqb_n dwla<1> dwla<0> dwlb<1> dwlb<0> l_clk_dqa l_clk_dqa_n l_clk_dqb 
+ l_clk_dqb_n l_lwea l_lweb l_sa_prea_n l_sa_preb_n l_saea_n l_saeb_n lb_ca<3> 
+ lb_ca<2> lb_ca<1> lb_ca<0> lb_cb<3> lb_cb<2> lb_cb<1> lb_cb<0> lb_ma<3> 
+ lb_ma<2> lb_ma<1> lb_ma<0> lb_mb<3> lb_mb<2> lb_mb<1> lb_mb<0> lb_tm_prea_n 
+ lb_tm_preb_n lt_ca<3> lt_ca<2> lt_ca<1> lt_ca<0> lt_cb<3> lt_cb<2> lt_cb<1> 
+ lt_cb<0> lt_ma<3> lt_ma<2> lt_ma<1> lt_ma<0> lt_mb<3> lt_mb<2> lt_mb<1> 
+ lt_mb<0> lt_tm_prea_n lt_tm_preb_n r_clk_dqa r_clk_dqa_n r_clk_dqb 
+ r_clk_dqb_n r_lwea r_lweb r_sa_prea_n r_sa_preb_n r_saea_n r_saeb_n rb_ca<3> 
+ rb_ca<2> rb_ca<1> rb_ca<0> rb_cb<3> rb_cb<2> rb_cb<1> rb_cb<0> rb_ma<3> 
+ rb_ma<2> rb_ma<1> rb_ma<0> rb_mb<3> rb_mb<2> rb_mb<1> rb_mb<0> rb_tm_prea_n 
+ rb_tm_preb_n rt_ca<3> rt_ca<2> rt_ca<1> rt_ca<0> rt_cb<3> rt_cb<2> rt_cb<1> 
+ rt_cb<0> rt_ma<3> rt_ma<2> rt_ma<1> rt_ma<0> rt_mb<3> rt_mb<2> rt_mb<1> 
+ rt_mb<0> rt_tm_prea_n rt_tm_preb_n stclka stclkb t_pxaa<3> t_pxaa<2> 
+ t_pxaa<1> t_pxaa<0> t_pxab<3> t_pxab<2> t_pxab<1> t_pxab<0> t_pxba_n<7> 
+ t_pxba_n<6> t_pxba_n<5> t_pxba_n<4> t_pxba_n<3> t_pxba_n<2> t_pxba_n<1> 
+ t_pxba_n<0> t_pxbb_n<7> t_pxbb_n<6> t_pxbb_n<5> t_pxbb_n<4> t_pxbb_n<3> 
+ t_pxbb_n<2> t_pxbb_n<1> t_pxbb_n<0> t_pxca_n<7> t_pxca_n<6> t_pxca_n<5> 
+ t_pxca_n<4> t_pxca_n<3> t_pxca_n<2> t_pxca_n<1> t_pxca_n<0> t_pxcb_n<7> 
+ t_pxcb_n<6> t_pxcb_n<5> t_pxcb_n<4> t_pxcb_n<3> t_pxcb_n<2> t_pxcb_n<1> 
+ t_pxcb_n<0> tm<9> tm<8> tm<7> tm<6> tm<5> tm<4> tm<3> tm<2> tm<1> tm<0> vdd 
+ vss wena wenb
** N=19585 EP=230 IP=0 FDC=3266
M0 vss 5 15 vss hvtnfet l=6e-08 w=6e-07 $X=965 $Y=37277 $D=616
M1 11 1 vss vss hvtnfet l=6e-08 w=6e-07 $X=1225 $Y=336 $D=616
M2 12 2 vss vss hvtnfet l=6e-08 w=6e-07 $X=1225 $Y=5566 $D=616
M3 13 3 vss vss hvtnfet l=6e-08 w=6e-07 $X=1225 $Y=6796 $D=616
M4 14 4 vss vss hvtnfet l=6e-08 w=6e-07 $X=1225 $Y=12026 $D=616
M5 lb_tm_preb_n 20 vss vss hvtnfet l=6e-08 w=1.287e-06 $X=1225 $Y=13280 $D=616
M6 lt_tm_preb_n 21 vss vss hvtnfet l=6e-08 w=1.287e-06 $X=1225 $Y=20124 $D=616
M7 vss 8 l_clk_dqb vss hvtnfet l=6e-08 w=1.26e-06 $X=1225 $Y=22041 $D=616
M8 vss 9 l_clk_dqb_n vss hvtnfet l=6e-08 w=1.26e-06 $X=1225 $Y=29007 $D=616
M9 l_lweb 10 vss vss hvtnfet l=6e-08 w=1.287e-06 $X=1225 $Y=30897 $D=616
M10 15 5 vss vss hvtnfet l=6e-08 w=6e-07 $X=1225 $Y=37277 $D=616
M11 16 4 vss vss hvtnfet l=6e-08 w=6e-07 $X=1225 $Y=38507 $D=616
M12 17 3 vss vss hvtnfet l=6e-08 w=6e-07 $X=1225 $Y=43737 $D=616
M13 18 6 vss vss hvtnfet l=6e-08 w=6e-07 $X=1225 $Y=44967 $D=616
M14 19 7 vss vss hvtnfet l=6e-08 w=6e-07 $X=1225 $Y=50197 $D=616
M15 vss 20 lb_tm_preb_n vss hvtnfet l=6e-08 w=1.287e-06 $X=1485 $Y=13280 $D=616
M16 vss 21 lt_tm_preb_n vss hvtnfet l=6e-08 w=1.287e-06 $X=1485 $Y=20124 $D=616
M17 l_clk_dqb 8 vss vss hvtnfet l=6e-08 w=1.26e-06 $X=1485 $Y=22041 $D=616
M18 l_clk_dqb_n 9 vss vss hvtnfet l=6e-08 w=1.26e-06 $X=1485 $Y=29007 $D=616
M19 vss 10 l_lweb vss hvtnfet l=6e-08 w=1.287e-06 $X=1485 $Y=30897 $D=616
M20 lb_cb<0> 11 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=1735 $Y=328 $D=616
M21 lb_cb<2> 12 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=1735 $Y=5316 $D=616
M22 lb_mb<0> 13 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=1735 $Y=6788 $D=616
M23 lb_mb<2> 14 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=1735 $Y=11776 $D=616
M24 l_saeb_n 15 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=1735 $Y=37027 $D=616
M25 lt_mb<2> 16 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=1735 $Y=38499 $D=616
M26 lt_mb<0> 17 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=1735 $Y=43487 $D=616
M27 lt_cb<2> 18 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=1735 $Y=44959 $D=616
M28 lt_cb<0> 19 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=1735 $Y=49947 $D=616
M29 vss 8 l_clk_dqb vss hvtnfet l=6e-08 w=1.26e-06 $X=1745 $Y=22041 $D=616
M30 vss 9 l_clk_dqb_n vss hvtnfet l=6e-08 w=1.26e-06 $X=1745 $Y=29007 $D=616
M31 vss 11 lb_cb<0> vss hvtnfet l=6e-08 w=8.58e-07 $X=1995 $Y=328 $D=616
M32 vss 12 lb_cb<2> vss hvtnfet l=6e-08 w=8.58e-07 $X=1995 $Y=5316 $D=616
M33 vss 13 lb_mb<0> vss hvtnfet l=6e-08 w=8.58e-07 $X=1995 $Y=6788 $D=616
M34 vss 14 lb_mb<2> vss hvtnfet l=6e-08 w=8.58e-07 $X=1995 $Y=11776 $D=616
M35 vss 24 20 vss hvtnfet l=6e-08 w=6e-07 $X=1995 $Y=13282 $D=616
M36 vss 25 21 vss hvtnfet l=6e-08 w=6e-07 $X=1995 $Y=20809 $D=616
M37 vss 15 l_saeb_n vss hvtnfet l=6e-08 w=8.58e-07 $X=1995 $Y=37027 $D=616
M38 vss 16 lt_mb<2> vss hvtnfet l=6e-08 w=8.58e-07 $X=1995 $Y=38499 $D=616
M39 vss 17 lt_mb<0> vss hvtnfet l=6e-08 w=8.58e-07 $X=1995 $Y=43487 $D=616
M40 vss 18 lt_cb<2> vss hvtnfet l=6e-08 w=8.58e-07 $X=1995 $Y=44959 $D=616
M41 vss 19 lt_cb<0> vss hvtnfet l=6e-08 w=8.58e-07 $X=1995 $Y=49947 $D=616
M42 8 clkb vss vss hvtnfet l=6e-08 w=1.05e-06 $X=2005 $Y=22251 $D=616
M43 9 23 vss vss hvtnfet l=6e-08 w=1.05e-06 $X=2005 $Y=29007 $D=616
M44 lb_cb<0> 11 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=2255 $Y=328 $D=616
M45 lb_cb<2> 12 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=2255 $Y=5316 $D=616
M46 lb_mb<0> 13 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=2255 $Y=6788 $D=616
M47 lb_mb<2> 14 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=2255 $Y=11776 $D=616
M48 l_saeb_n 15 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=2255 $Y=37027 $D=616
M49 lt_mb<2> 16 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=2255 $Y=38499 $D=616
M50 lt_mb<0> 17 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=2255 $Y=43487 $D=616
M51 lt_cb<2> 18 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=2255 $Y=44959 $D=616
M52 lt_cb<0> 19 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=2255 $Y=49947 $D=616
M53 vss 15 l_saeb_n vss hvtnfet l=6e-08 w=8.58e-07 $X=2515 $Y=37027 $D=616
M54 vss 34 lb_cb<1> vss hvtnfet l=6e-08 w=8.58e-07 $X=2765 $Y=328 $D=616
M55 vss 35 lb_cb<3> vss hvtnfet l=6e-08 w=8.58e-07 $X=2765 $Y=5316 $D=616
M56 vss 36 lb_mb<1> vss hvtnfet l=6e-08 w=8.58e-07 $X=2765 $Y=6788 $D=616
M57 vss 37 lb_mb<3> vss hvtnfet l=6e-08 w=8.58e-07 $X=2765 $Y=11776 $D=616
M58 vss 39 lt_mb<3> vss hvtnfet l=6e-08 w=8.58e-07 $X=2765 $Y=38499 $D=616
M59 vss 40 lt_mb<1> vss hvtnfet l=6e-08 w=8.58e-07 $X=2765 $Y=43487 $D=616
M60 vss 41 lt_cb<3> vss hvtnfet l=6e-08 w=8.58e-07 $X=2765 $Y=44959 $D=616
M61 vss 42 lt_cb<1> vss hvtnfet l=6e-08 w=8.58e-07 $X=2765 $Y=49947 $D=616
M62 l_saeb_n 15 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=2775 $Y=37027 $D=616
M63 909 26 vss vss hvtnfet l=6e-08 w=1.8e-07 $X=2821 $Y=17143 $D=616
M64 26 28 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=2821 $Y=17812 $D=616
M65 4 29 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=2821 $Y=18983 $D=616
M66 910 4 vss vss hvtnfet l=6e-08 w=1.8e-07 $X=2821 $Y=19609 $D=616
M67 911 27 vss vss hvtnfet l=6e-08 w=1.8e-07 $X=2821 $Y=24063 $D=616
M68 27 30 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=2821 $Y=24732 $D=616
M69 3 31 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=2821 $Y=25903 $D=616
M70 912 3 vss vss hvtnfet l=6e-08 w=1.8e-07 $X=2821 $Y=26529 $D=616
M71 lb_cb<1> 34 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=3025 $Y=328 $D=616
M72 lb_cb<3> 35 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=3025 $Y=5316 $D=616
M73 lb_mb<1> 36 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=3025 $Y=6788 $D=616
M74 lb_mb<3> 37 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=3025 $Y=11776 $D=616
M75 lt_mb<3> 39 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=3025 $Y=38499 $D=616
M76 lt_mb<1> 40 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=3025 $Y=43487 $D=616
M77 lt_cb<3> 41 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=3025 $Y=44959 $D=616
M78 lt_cb<1> 42 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=3025 $Y=49947 $D=616
M79 28 33 909 vss hvtnfet l=6e-08 w=1.8e-07 $X=3081 $Y=17143 $D=616
M80 vss 28 26 vss hvtnfet l=6e-08 w=1.37e-07 $X=3081 $Y=17812 $D=616
M81 vss 29 4 vss hvtnfet l=6e-08 w=1.37e-07 $X=3081 $Y=18983 $D=616
M82 29 33 910 vss hvtnfet l=6e-08 w=1.8e-07 $X=3081 $Y=19609 $D=616
M83 30 33 911 vss hvtnfet l=6e-08 w=1.8e-07 $X=3081 $Y=24063 $D=616
M84 vss 30 27 vss hvtnfet l=6e-08 w=1.37e-07 $X=3081 $Y=24732 $D=616
M85 vss 31 3 vss hvtnfet l=6e-08 w=1.37e-07 $X=3081 $Y=25903 $D=616
M86 31 33 912 vss hvtnfet l=6e-08 w=1.8e-07 $X=3081 $Y=26529 $D=616
M87 vss 34 lb_cb<1> vss hvtnfet l=6e-08 w=8.58e-07 $X=3285 $Y=328 $D=616
M88 vss 35 lb_cb<3> vss hvtnfet l=6e-08 w=8.58e-07 $X=3285 $Y=5316 $D=616
M89 vss 36 lb_mb<1> vss hvtnfet l=6e-08 w=8.58e-07 $X=3285 $Y=6788 $D=616
M90 vss 37 lb_mb<3> vss hvtnfet l=6e-08 w=8.58e-07 $X=3285 $Y=11776 $D=616
M91 vss 51 l_sa_preb_n vss hvtnfet l=6e-08 w=8.58e-07 $X=3285 $Y=37027 $D=616
M92 vss 39 lt_mb<3> vss hvtnfet l=6e-08 w=8.58e-07 $X=3285 $Y=38499 $D=616
M93 vss 40 lt_mb<1> vss hvtnfet l=6e-08 w=8.58e-07 $X=3285 $Y=43487 $D=616
M94 vss 41 lt_cb<3> vss hvtnfet l=6e-08 w=8.58e-07 $X=3285 $Y=44959 $D=616
M95 vss 42 lt_cb<1> vss hvtnfet l=6e-08 w=8.58e-07 $X=3285 $Y=49947 $D=616
M96 vss ab<2> 44 vss hvtnfet l=6e-08 w=2.74e-07 $X=3396 $Y=13476 $D=616
M97 l_sa_preb_n 51 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=3545 $Y=37027 $D=616
M98 913 43 vss vss hvtnfet l=6e-08 w=8.23e-07 $X=3591 $Y=17143 $D=616
M99 914 43 vss vss hvtnfet l=6e-08 w=8.23e-07 $X=3591 $Y=18966 $D=616
M100 915 43 vss vss hvtnfet l=6e-08 w=8.23e-07 $X=3591 $Y=24063 $D=616
M101 916 43 vss vss hvtnfet l=6e-08 w=8.23e-07 $X=3591 $Y=25886 $D=616
M102 52 stclkb vss vss hvtnfet l=6e-08 w=2.74e-07 $X=3705 $Y=30668 $D=616
M103 vss 47 34 vss hvtnfet l=6e-08 w=6e-07 $X=3795 $Y=336 $D=616
M104 vss 48 35 vss hvtnfet l=6e-08 w=6e-07 $X=3795 $Y=5566 $D=616
M105 vss 27 36 vss hvtnfet l=6e-08 w=6e-07 $X=3795 $Y=6796 $D=616
M106 vss 26 37 vss hvtnfet l=6e-08 w=6e-07 $X=3795 $Y=12026 $D=616
M107 vss 26 39 vss hvtnfet l=6e-08 w=6e-07 $X=3795 $Y=38507 $D=616
M108 vss 27 40 vss hvtnfet l=6e-08 w=6e-07 $X=3795 $Y=43737 $D=616
M109 vss 49 41 vss hvtnfet l=6e-08 w=6e-07 $X=3795 $Y=44967 $D=616
M110 vss 50 42 vss hvtnfet l=6e-08 w=6e-07 $X=3795 $Y=50197 $D=616
M111 vss 51 l_sa_preb_n vss hvtnfet l=6e-08 w=8.58e-07 $X=3805 $Y=37027 $D=616
M112 917 45 913 vss hvtnfet l=6e-08 w=5.49e-07 $X=3861 $Y=17143 $D=616
M113 918 45 914 vss hvtnfet l=6e-08 w=5.49e-07 $X=3861 $Y=19240 $D=616
M114 919 46 915 vss hvtnfet l=6e-08 w=5.49e-07 $X=3861 $Y=24063 $D=616
M115 920 46 916 vss hvtnfet l=6e-08 w=5.49e-07 $X=3861 $Y=26160 $D=616
M116 53 44 vss vss hvtnfet l=6e-08 w=2.74e-07 $X=3906 $Y=13476 $D=616
M117 vss clkb 43 vss hvtnfet l=6e-08 w=6e-07 $X=4066 $Y=32403 $D=616
M118 28 53 917 vss hvtnfet l=6e-08 w=5.49e-07 $X=4121 $Y=17143 $D=616
M119 29 44 918 vss hvtnfet l=6e-08 w=5.49e-07 $X=4121 $Y=19240 $D=616
M120 30 53 919 vss hvtnfet l=6e-08 w=5.49e-07 $X=4121 $Y=24063 $D=616
M121 31 44 920 vss hvtnfet l=6e-08 w=5.49e-07 $X=4121 $Y=26160 $D=616
M122 vss 52 59 vss hvtnfet l=6e-08 w=5.49e-07 $X=4215 $Y=30668 $D=616
M123 vss 55 51 vss hvtnfet l=6e-08 w=6e-07 $X=4315 $Y=37277 $D=616
M124 43 clkb vss vss hvtnfet l=6e-08 w=6e-07 $X=4326 $Y=32403 $D=616
M125 vss ab<3> 46 vss hvtnfet l=6e-08 w=2.74e-07 $X=4416 $Y=13476 $D=616
M126 59 56 vss vss hvtnfet l=6e-08 w=5.49e-07 $X=4475 $Y=30668 $D=616
M127 b_pxab<0> 60 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=4550 $Y=336 $D=616
M128 60 61 vss vss hvtnfet l=6e-08 w=5e-07 $X=4550 $Y=6701 $D=616
M129 61 62 vss vss hvtnfet l=6e-08 w=3e-07 $X=4550 $Y=7831 $D=616
M130 921 57 vss vss hvtnfet l=6e-08 w=4.11e-07 $X=4550 $Y=11276 $D=616
M131 922 57 vss vss hvtnfet l=6e-08 w=4.11e-07 $X=4550 $Y=39446 $D=616
M132 64 63 vss vss hvtnfet l=6e-08 w=3e-07 $X=4550 $Y=43002 $D=616
M133 65 64 vss vss hvtnfet l=6e-08 w=5e-07 $X=4550 $Y=43932 $D=616
M134 t_pxab<0> 65 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=4550 $Y=49512 $D=616
M135 vss 60 b_pxab<0> vss hvtnfet l=6e-08 w=1.285e-06 $X=4810 $Y=336 $D=616
M136 vss 61 60 vss hvtnfet l=6e-08 w=5e-07 $X=4810 $Y=6701 $D=616
M137 vss 62 61 vss hvtnfet l=6e-08 w=3e-07 $X=4810 $Y=7831 $D=616
M138 62 24 921 vss hvtnfet l=6e-08 w=4.11e-07 $X=4810 $Y=11276 $D=616
M139 63 25 922 vss hvtnfet l=6e-08 w=4.11e-07 $X=4810 $Y=39446 $D=616
M140 vss 63 64 vss hvtnfet l=6e-08 w=3e-07 $X=4810 $Y=43002 $D=616
M141 vss 64 65 vss hvtnfet l=6e-08 w=5e-07 $X=4810 $Y=43932 $D=616
M142 vss 65 t_pxab<0> vss hvtnfet l=6e-08 w=1.285e-06 $X=4810 $Y=49512 $D=616
M143 45 46 vss vss hvtnfet l=6e-08 w=2.74e-07 $X=4926 $Y=13476 $D=616
M144 vss 66 586 vss hvtnfet l=1.4e-07 w=3.2e-07 $X=4939 $Y=37127 $D=616
M145 vss 59 56 vss hvtnfet l=6e-08 w=5.49e-07 $X=4985 $Y=30668 $D=616
M146 vss 58 587 vss hvtnfet l=6e-08 w=3.2e-07 $X=5069 $Y=32828 $D=616
M147 923 67 vss vss hvtnfet l=6e-08 w=1.8e-07 $X=5141 $Y=17143 $D=616
M148 67 73 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=5141 $Y=17812 $D=616
M149 68 74 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=5141 $Y=18983 $D=616
M150 924 68 vss vss hvtnfet l=6e-08 w=1.8e-07 $X=5141 $Y=19609 $D=616
M151 925 69 vss vss hvtnfet l=6e-08 w=1.8e-07 $X=5141 $Y=24063 $D=616
M152 69 75 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=5141 $Y=24732 $D=616
M153 57 76 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=5141 $Y=25903 $D=616
M154 926 57 vss vss hvtnfet l=6e-08 w=1.8e-07 $X=5141 $Y=26529 $D=616
M155 56 70 vss vss hvtnfet l=6e-08 w=5.49e-07 $X=5245 $Y=30668 $D=616
M156 66 71 vss vss hvtnfet l=1.4e-07 w=3.2e-07 $X=5279 $Y=37127 $D=616
M157 b_pxab<1> 78 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=5320 $Y=336 $D=616
M158 78 79 vss vss hvtnfet l=6e-08 w=5e-07 $X=5320 $Y=6701 $D=616
M159 79 80 vss vss hvtnfet l=6e-08 w=3e-07 $X=5320 $Y=7831 $D=616
M160 927 24 80 vss hvtnfet l=6e-08 w=4.11e-07 $X=5320 $Y=11276 $D=616
M161 928 25 81 vss hvtnfet l=6e-08 w=4.11e-07 $X=5320 $Y=39446 $D=616
M162 82 81 vss vss hvtnfet l=6e-08 w=3e-07 $X=5320 $Y=43002 $D=616
M163 83 82 vss vss hvtnfet l=6e-08 w=5e-07 $X=5320 $Y=43932 $D=616
M164 t_pxab<1> 83 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=5320 $Y=49512 $D=616
M165 73 33 923 vss hvtnfet l=6e-08 w=1.8e-07 $X=5401 $Y=17143 $D=616
M166 vss 73 67 vss hvtnfet l=6e-08 w=1.37e-07 $X=5401 $Y=17812 $D=616
M167 vss 74 68 vss hvtnfet l=6e-08 w=1.37e-07 $X=5401 $Y=18983 $D=616
M168 74 33 924 vss hvtnfet l=6e-08 w=1.8e-07 $X=5401 $Y=19609 $D=616
M169 75 33 925 vss hvtnfet l=6e-08 w=1.8e-07 $X=5401 $Y=24063 $D=616
M170 vss 75 69 vss hvtnfet l=6e-08 w=1.37e-07 $X=5401 $Y=24732 $D=616
M171 vss 76 57 vss hvtnfet l=6e-08 w=1.37e-07 $X=5401 $Y=25903 $D=616
M172 76 33 926 vss hvtnfet l=6e-08 w=1.8e-07 $X=5401 $Y=26529 $D=616
M173 929 72 vss vss hvtnfet l=6e-08 w=6.4e-07 $X=5579 $Y=32508 $D=616
M174 vss 78 b_pxab<1> vss hvtnfet l=6e-08 w=1.285e-06 $X=5580 $Y=336 $D=616
M175 vss 79 78 vss hvtnfet l=6e-08 w=5e-07 $X=5580 $Y=6701 $D=616
M176 vss 80 79 vss hvtnfet l=6e-08 w=3e-07 $X=5580 $Y=7831 $D=616
M177 vss 69 927 vss hvtnfet l=6e-08 w=4.11e-07 $X=5580 $Y=11276 $D=616
M178 vss 69 928 vss hvtnfet l=6e-08 w=4.11e-07 $X=5580 $Y=39446 $D=616
M179 vss 81 82 vss hvtnfet l=6e-08 w=3e-07 $X=5580 $Y=43002 $D=616
M180 vss 82 83 vss hvtnfet l=6e-08 w=5e-07 $X=5580 $Y=43932 $D=616
M181 vss 83 t_pxab<1> vss hvtnfet l=6e-08 w=1.285e-06 $X=5580 $Y=49512 $D=616
M182 vss ab<5> 86 vss hvtnfet l=6e-08 w=2.74e-07 $X=5716 $Y=13476 $D=616
M183 5 85 929 vss hvtnfet l=6e-08 w=6.4e-07 $X=5839 $Y=32508 $D=616
M184 930 43 vss vss hvtnfet l=6e-08 w=8.23e-07 $X=5911 $Y=17143 $D=616
M185 931 43 vss vss hvtnfet l=6e-08 w=8.23e-07 $X=5911 $Y=18966 $D=616
M186 932 43 vss vss hvtnfet l=6e-08 w=8.23e-07 $X=5911 $Y=24063 $D=616
M187 933 43 vss vss hvtnfet l=6e-08 w=8.23e-07 $X=5911 $Y=25886 $D=616
M188 70 clkb vss vss hvtnfet l=6e-08 w=6e-07 $X=6015 $Y=30668 $D=616
M189 vss ddqb 71 vss hvtnfet l=6e-08 w=2.4e-07 $X=6079 $Y=37292 $D=616
M190 b_pxab<2> 90 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=6090 $Y=336 $D=616
M191 90 91 vss vss hvtnfet l=6e-08 w=5e-07 $X=6090 $Y=6701 $D=616
M192 91 92 vss vss hvtnfet l=6e-08 w=3e-07 $X=6090 $Y=7831 $D=616
M193 934 68 vss vss hvtnfet l=6e-08 w=4.11e-07 $X=6090 $Y=11276 $D=616
M194 935 68 vss vss hvtnfet l=6e-08 w=4.11e-07 $X=6090 $Y=39446 $D=616
M195 94 93 vss vss hvtnfet l=6e-08 w=3e-07 $X=6090 $Y=43002 $D=616
M196 95 94 vss vss hvtnfet l=6e-08 w=5e-07 $X=6090 $Y=43932 $D=616
M197 t_pxab<2> 95 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=6090 $Y=49512 $D=616
M198 936 87 930 vss hvtnfet l=6e-08 w=5.49e-07 $X=6181 $Y=17143 $D=616
M199 937 87 931 vss hvtnfet l=6e-08 w=5.49e-07 $X=6181 $Y=19240 $D=616
M200 938 88 932 vss hvtnfet l=6e-08 w=5.49e-07 $X=6181 $Y=24063 $D=616
M201 939 88 933 vss hvtnfet l=6e-08 w=5.49e-07 $X=6181 $Y=26160 $D=616
M202 97 86 vss vss hvtnfet l=6e-08 w=2.74e-07 $X=6226 $Y=13476 $D=616
M203 71 ddqb_n vss vss hvtnfet l=6e-08 w=2.4e-07 $X=6339 $Y=37292 $D=616
M204 vss 90 b_pxab<2> vss hvtnfet l=6e-08 w=1.285e-06 $X=6350 $Y=336 $D=616
M205 vss 91 90 vss hvtnfet l=6e-08 w=5e-07 $X=6350 $Y=6701 $D=616
M206 vss 92 91 vss hvtnfet l=6e-08 w=3e-07 $X=6350 $Y=7831 $D=616
M207 92 24 934 vss hvtnfet l=6e-08 w=4.11e-07 $X=6350 $Y=11276 $D=616
M208 93 25 935 vss hvtnfet l=6e-08 w=4.11e-07 $X=6350 $Y=39446 $D=616
M209 vss 93 94 vss hvtnfet l=6e-08 w=3e-07 $X=6350 $Y=43002 $D=616
M210 vss 94 95 vss hvtnfet l=6e-08 w=5e-07 $X=6350 $Y=43932 $D=616
M211 vss 95 t_pxab<2> vss hvtnfet l=6e-08 w=1.285e-06 $X=6350 $Y=49512 $D=616
M212 73 97 936 vss hvtnfet l=6e-08 w=5.49e-07 $X=6441 $Y=17143 $D=616
M213 74 86 937 vss hvtnfet l=6e-08 w=5.49e-07 $X=6441 $Y=19240 $D=616
M214 75 97 938 vss hvtnfet l=6e-08 w=5.49e-07 $X=6441 $Y=24063 $D=616
M215 76 86 939 vss hvtnfet l=6e-08 w=5.49e-07 $X=6441 $Y=26160 $D=616
M216 85 89 vss vss hvtnfet l=6e-08 w=3.2e-07 $X=6524 $Y=32828 $D=616
M217 142 clkb 595 vss hvtnfet l=6e-08 w=8e-07 $X=6525 $Y=30668 $D=616
M218 vss ab<6> 88 vss hvtnfet l=6e-08 w=2.74e-07 $X=6736 $Y=13476 $D=616
M219 595 clkb 142 vss hvtnfet l=6e-08 w=8e-07 $X=6785 $Y=30668 $D=616
M220 b_pxab<3> 99 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=6860 $Y=336 $D=616
M221 99 100 vss vss hvtnfet l=6e-08 w=5e-07 $X=6860 $Y=6701 $D=616
M222 100 101 vss vss hvtnfet l=6e-08 w=3e-07 $X=6860 $Y=7831 $D=616
M223 940 24 101 vss hvtnfet l=6e-08 w=4.11e-07 $X=6860 $Y=11276 $D=616
M224 941 25 102 vss hvtnfet l=6e-08 w=4.11e-07 $X=6860 $Y=39446 $D=616
M225 103 102 vss vss hvtnfet l=6e-08 w=3e-07 $X=6860 $Y=43002 $D=616
M226 104 103 vss vss hvtnfet l=6e-08 w=5e-07 $X=6860 $Y=43932 $D=616
M227 t_pxab<3> 104 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=6860 $Y=49512 $D=616
M228 109 85 vss vss hvtnfet l=6e-08 w=3.2e-07 $X=7034 $Y=32828 $D=616
M229 89 58 vss vss hvtnfet l=6e-08 w=3.2e-07 $X=7069 $Y=37292 $D=616
M230 vss 99 b_pxab<3> vss hvtnfet l=6e-08 w=1.285e-06 $X=7120 $Y=336 $D=616
M231 vss 100 99 vss hvtnfet l=6e-08 w=5e-07 $X=7120 $Y=6701 $D=616
M232 vss 101 100 vss hvtnfet l=6e-08 w=3e-07 $X=7120 $Y=7831 $D=616
M233 vss 67 940 vss hvtnfet l=6e-08 w=4.11e-07 $X=7120 $Y=11276 $D=616
M234 vss 67 941 vss hvtnfet l=6e-08 w=4.11e-07 $X=7120 $Y=39446 $D=616
M235 vss 102 103 vss hvtnfet l=6e-08 w=3e-07 $X=7120 $Y=43002 $D=616
M236 vss 103 104 vss hvtnfet l=6e-08 w=5e-07 $X=7120 $Y=43932 $D=616
M237 vss 104 t_pxab<3> vss hvtnfet l=6e-08 w=1.285e-06 $X=7120 $Y=49512 $D=616
M238 87 88 vss vss hvtnfet l=6e-08 w=2.74e-07 $X=7246 $Y=13476 $D=616
M239 595 59 vss vss hvtnfet l=6e-08 w=8e-07 $X=7295 $Y=30668 $D=616
M240 942 105 vss vss hvtnfet l=6e-08 w=1.8e-07 $X=7461 $Y=17143 $D=616
M241 943 106 vss vss hvtnfet l=6e-08 w=1.8e-07 $X=7461 $Y=19609 $D=616
M242 944 107 vss vss hvtnfet l=6e-08 w=1.8e-07 $X=7461 $Y=24063 $D=616
M243 945 108 vss vss hvtnfet l=6e-08 w=1.8e-07 $X=7461 $Y=26529 $D=616
M244 105 111 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=7476 $Y=17812 $D=616
M245 106 112 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=7476 $Y=18983 $D=616
M246 107 113 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=7476 $Y=24732 $D=616
M247 108 114 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=7476 $Y=25903 $D=616
M248 vss 59 595 vss hvtnfet l=6e-08 w=8e-07 $X=7555 $Y=30668 $D=616
M249 vss 110 89 vss hvtnfet l=1.2e-07 w=1.5e-07 $X=7579 $Y=37297 $D=616
M250 vss 109 119 vss hvtnfet l=2.5e-07 w=3.5e-07 $X=7604 $Y=32613 $D=616
M251 b_pxbb_n<0> 115 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=7630 $Y=336 $D=616
M252 115 116 vss vss hvtnfet l=6e-08 w=5e-07 $X=7630 $Y=6701 $D=616
M253 116 107 vss vss hvtnfet l=6e-08 w=3e-07 $X=7630 $Y=7831 $D=616
M254 117 107 vss vss hvtnfet l=6e-08 w=3e-07 $X=7630 $Y=43002 $D=616
M255 118 117 vss vss hvtnfet l=6e-08 w=5e-07 $X=7630 $Y=43932 $D=616
M256 t_pxbb_n<0> 118 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=7630 $Y=49512 $D=616
M257 111 33 942 vss hvtnfet l=6e-08 w=1.8e-07 $X=7721 $Y=17143 $D=616
M258 112 33 943 vss hvtnfet l=6e-08 w=1.8e-07 $X=7721 $Y=19609 $D=616
M259 113 33 944 vss hvtnfet l=6e-08 w=1.8e-07 $X=7721 $Y=24063 $D=616
M260 114 33 945 vss hvtnfet l=6e-08 w=1.8e-07 $X=7721 $Y=26529 $D=616
M261 vss 111 105 vss hvtnfet l=6e-08 w=1.37e-07 $X=7736 $Y=17812 $D=616
M262 vss 112 106 vss hvtnfet l=6e-08 w=1.37e-07 $X=7736 $Y=18983 $D=616
M263 vss 113 107 vss hvtnfet l=6e-08 w=1.37e-07 $X=7736 $Y=24732 $D=616
M264 vss 114 108 vss hvtnfet l=6e-08 w=1.37e-07 $X=7736 $Y=25903 $D=616
M265 vss 115 b_pxbb_n<0> vss hvtnfet l=6e-08 w=1.285e-06 $X=7890 $Y=336 $D=616
M266 vss 116 115 vss hvtnfet l=6e-08 w=5e-07 $X=7890 $Y=6701 $D=616
M267 vss 107 116 vss hvtnfet l=6e-08 w=3e-07 $X=7890 $Y=7831 $D=616
M268 vss 107 117 vss hvtnfet l=6e-08 w=3e-07 $X=7890 $Y=43002 $D=616
M269 vss 117 118 vss hvtnfet l=6e-08 w=5e-07 $X=7890 $Y=43932 $D=616
M270 vss 118 t_pxbb_n<0> vss hvtnfet l=6e-08 w=1.285e-06 $X=7890 $Y=49512 $D=616
M271 120 119 vss vss hvtnfet l=6e-08 w=3.5e-07 $X=8054 $Y=32613 $D=616
M272 110 89 vss vss hvtnfet l=6e-08 w=3e-07 $X=8149 $Y=37257 $D=616
M273 946 43 vss vss hvtnfet l=6e-08 w=8.23e-07 $X=8231 $Y=17143 $D=616
M274 947 43 vss vss hvtnfet l=6e-08 w=8.23e-07 $X=8231 $Y=18966 $D=616
M275 948 43 vss vss hvtnfet l=6e-08 w=8.23e-07 $X=8231 $Y=24063 $D=616
M276 949 43 vss vss hvtnfet l=6e-08 w=8.23e-07 $X=8231 $Y=25886 $D=616
M277 b_pxbb_n<1> 125 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=8400 $Y=336 $D=616
M278 125 126 vss vss hvtnfet l=6e-08 w=5e-07 $X=8400 $Y=6701 $D=616
M279 126 108 vss vss hvtnfet l=6e-08 w=3e-07 $X=8400 $Y=7831 $D=616
M280 127 108 vss vss hvtnfet l=6e-08 w=3e-07 $X=8400 $Y=43002 $D=616
M281 128 127 vss vss hvtnfet l=6e-08 w=5e-07 $X=8400 $Y=43932 $D=616
M282 t_pxbb_n<1> 128 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=8400 $Y=49512 $D=616
M283 vss 122 121 vss hvtnfet l=6e-08 w=2.74e-07 $X=8466 $Y=13476 $D=616
M284 950 121 946 vss hvtnfet l=6e-08 w=5.49e-07 $X=8501 $Y=17417 $D=616
M285 951 121 947 vss hvtnfet l=6e-08 w=5.49e-07 $X=8501 $Y=18966 $D=616
M286 952 122 948 vss hvtnfet l=6e-08 w=5.49e-07 $X=8501 $Y=24337 $D=616
M287 953 122 949 vss hvtnfet l=6e-08 w=5.49e-07 $X=8501 $Y=25886 $D=616
M288 123 123 vss vss hvtnfet l=6e-08 w=2e-07 $X=8594 $Y=11546 $D=616
M289 954 120 55 vss hvtnfet l=6e-08 w=6.4e-07 $X=8619 $Y=32508 $D=616
M290 dwlb<0> 124 vss vss hvtnfet l=6e-08 w=3e-07 $X=8659 $Y=31098 $D=616
M291 25 124 vss vss hvtnfet l=6e-08 w=3e-07 $X=8659 $Y=37457 $D=616
M292 vss 125 b_pxbb_n<1> vss hvtnfet l=6e-08 w=1.285e-06 $X=8660 $Y=336 $D=616
M293 vss 126 125 vss hvtnfet l=6e-08 w=5e-07 $X=8660 $Y=6701 $D=616
M294 vss 108 126 vss hvtnfet l=6e-08 w=3e-07 $X=8660 $Y=7831 $D=616
M295 vss 108 127 vss hvtnfet l=6e-08 w=3e-07 $X=8660 $Y=43002 $D=616
M296 vss 127 128 vss hvtnfet l=6e-08 w=5e-07 $X=8660 $Y=43932 $D=616
M297 vss 128 t_pxbb_n<1> vss hvtnfet l=6e-08 w=1.285e-06 $X=8660 $Y=49512 $D=616
M298 955 129 950 vss hvtnfet l=6e-08 w=5.49e-07 $X=8761 $Y=17417 $D=616
M299 956 129 951 vss hvtnfet l=6e-08 w=5.49e-07 $X=8761 $Y=18966 $D=616
M300 957 129 952 vss hvtnfet l=6e-08 w=5.49e-07 $X=8761 $Y=24337 $D=616
M301 958 129 953 vss hvtnfet l=6e-08 w=5.49e-07 $X=8761 $Y=25886 $D=616
M302 vss 131 123 vss hvtnfet l=6e-08 w=2e-07 $X=8854 $Y=11546 $D=616
M303 vss vdd 954 vss hvtnfet l=6e-08 w=6.4e-07 $X=8879 $Y=32508 $D=616
M304 vss 124 dwlb<0> vss hvtnfet l=6e-08 w=3e-07 $X=8919 $Y=31098 $D=616
M305 vss 124 25 vss hvtnfet l=6e-08 w=3e-07 $X=8919 $Y=37457 $D=616
M306 122 ab<9> vss vss hvtnfet l=6e-08 w=2.74e-07 $X=8976 $Y=13476 $D=616
M307 111 132 955 vss hvtnfet l=6e-08 w=5.49e-07 $X=9021 $Y=17417 $D=616
M308 112 133 956 vss hvtnfet l=6e-08 w=5.49e-07 $X=9021 $Y=18966 $D=616
M309 113 132 957 vss hvtnfet l=6e-08 w=5.49e-07 $X=9021 $Y=24337 $D=616
M310 114 133 958 vss hvtnfet l=6e-08 w=5.49e-07 $X=9021 $Y=25886 $D=616
M311 b_pxbb_n<2> 135 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=9170 $Y=336 $D=616
M312 135 136 vss vss hvtnfet l=6e-08 w=5e-07 $X=9170 $Y=6701 $D=616
M313 136 137 vss vss hvtnfet l=6e-08 w=3e-07 $X=9170 $Y=7831 $D=616
M314 138 137 vss vss hvtnfet l=6e-08 w=3e-07 $X=9170 $Y=43002 $D=616
M315 139 138 vss vss hvtnfet l=6e-08 w=5e-07 $X=9170 $Y=43932 $D=616
M316 t_pxbb_n<2> 139 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=9170 $Y=49512 $D=616
M317 dwlb<0> 142 vss vss hvtnfet l=6e-08 w=3e-07 $X=9429 $Y=31098 $D=616
M318 25 143 vss vss hvtnfet l=6e-08 w=3e-07 $X=9429 $Y=37457 $D=616
M319 vss 135 b_pxbb_n<2> vss hvtnfet l=6e-08 w=1.285e-06 $X=9430 $Y=336 $D=616
M320 vss 136 135 vss hvtnfet l=6e-08 w=5e-07 $X=9430 $Y=6701 $D=616
M321 vss 137 136 vss hvtnfet l=6e-08 w=3e-07 $X=9430 $Y=7831 $D=616
M322 vss 137 138 vss hvtnfet l=6e-08 w=3e-07 $X=9430 $Y=43002 $D=616
M323 vss 138 139 vss hvtnfet l=6e-08 w=5e-07 $X=9430 $Y=43932 $D=616
M324 vss 139 t_pxbb_n<2> vss hvtnfet l=6e-08 w=1.285e-06 $X=9430 $Y=49512 $D=616
M325 vss 140 1 vss hvtnfet l=6e-08 w=2e-07 $X=9586 $Y=11276 $D=616
M326 vss 141 7 vss hvtnfet l=6e-08 w=2e-07 $X=9586 $Y=39657 $D=616
M327 vss 142 dwlb<0> vss hvtnfet l=6e-08 w=3e-07 $X=9689 $Y=31098 $D=616
M328 vss 143 25 vss hvtnfet l=6e-08 w=3e-07 $X=9689 $Y=37457 $D=616
M329 b_pxbb_n<3> 146 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=9940 $Y=336 $D=616
M330 146 147 vss vss hvtnfet l=6e-08 w=5e-07 $X=9940 $Y=6701 $D=616
M331 147 148 vss vss hvtnfet l=6e-08 w=3e-07 $X=9940 $Y=7831 $D=616
M332 149 148 vss vss hvtnfet l=6e-08 w=3e-07 $X=9940 $Y=43002 $D=616
M333 150 149 vss vss hvtnfet l=6e-08 w=5e-07 $X=9940 $Y=43932 $D=616
M334 t_pxbb_n<3> 150 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=9940 $Y=49512 $D=616
M335 vss ab<8> 129 vss hvtnfet l=6e-08 w=2.74e-07 $X=9986 $Y=13476 $D=616
M336 959 145 vss vss hvtnfet l=6e-08 w=4.11e-07 $X=10096 $Y=11276 $D=616
M337 960 145 vss vss hvtnfet l=6e-08 w=4.11e-07 $X=10096 $Y=39446 $D=616
M338 dwlb<1> 142 vss vss hvtnfet l=6e-08 w=3e-07 $X=10199 $Y=31098 $D=616
M339 24 143 vss vss hvtnfet l=6e-08 w=3e-07 $X=10199 $Y=37457 $D=616
M340 vss 146 b_pxbb_n<3> vss hvtnfet l=6e-08 w=1.285e-06 $X=10200 $Y=336 $D=616
M341 vss 147 146 vss hvtnfet l=6e-08 w=5e-07 $X=10200 $Y=6701 $D=616
M342 vss 148 147 vss hvtnfet l=6e-08 w=3e-07 $X=10200 $Y=7831 $D=616
M343 vss 148 149 vss hvtnfet l=6e-08 w=3e-07 $X=10200 $Y=43002 $D=616
M344 vss 149 150 vss hvtnfet l=6e-08 w=5e-07 $X=10200 $Y=43932 $D=616
M345 vss 150 t_pxbb_n<3> vss hvtnfet l=6e-08 w=1.285e-06 $X=10200 $Y=49512 $D=616
M346 160 129 vss vss hvtnfet l=6e-08 w=2.74e-07 $X=10246 $Y=13476 $D=616
M347 140 dwlb<1> 959 vss hvtnfet l=6e-08 w=4.11e-07 $X=10356 $Y=11276 $D=616
M348 141 dwlb<0> 960 vss hvtnfet l=6e-08 w=4.11e-07 $X=10356 $Y=39446 $D=616
M349 vss 153 124 vss hvtnfet l=6e-08 w=4e-07 $X=10406 $Y=32543 $D=616
M350 vss 142 dwlb<1> vss hvtnfet l=6e-08 w=3e-07 $X=10459 $Y=31098 $D=616
M351 vss 143 24 vss hvtnfet l=6e-08 w=3e-07 $X=10459 $Y=37457 $D=616
M352 b_pxbb_n<4> 156 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=10710 $Y=336 $D=616
M353 156 157 vss vss hvtnfet l=6e-08 w=5e-07 $X=10710 $Y=6701 $D=616
M354 157 105 vss vss hvtnfet l=6e-08 w=3e-07 $X=10710 $Y=7831 $D=616
M355 158 105 vss vss hvtnfet l=6e-08 w=3e-07 $X=10710 $Y=43002 $D=616
M356 159 158 vss vss hvtnfet l=6e-08 w=5e-07 $X=10710 $Y=43932 $D=616
M357 t_pxbb_n<4> 159 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=10710 $Y=49512 $D=616
M358 vss 132 133 vss hvtnfet l=6e-08 w=2.74e-07 $X=10846 $Y=13476 $D=616
M359 961 132 168 vss hvtnfet l=6e-08 w=5.49e-07 $X=10861 $Y=17417 $D=616
M360 962 133 169 vss hvtnfet l=6e-08 w=5.49e-07 $X=10861 $Y=18966 $D=616
M361 963 132 170 vss hvtnfet l=6e-08 w=5.49e-07 $X=10861 $Y=24337 $D=616
M362 964 133 171 vss hvtnfet l=6e-08 w=5.49e-07 $X=10861 $Y=25886 $D=616
M363 965 dwlb<1> 162 vss hvtnfet l=6e-08 w=4.11e-07 $X=10866 $Y=11276 $D=616
M364 966 dwlb<0> 163 vss hvtnfet l=6e-08 w=4.11e-07 $X=10866 $Y=39446 $D=616
M365 dwlb<1> 153 vss vss hvtnfet l=6e-08 w=3e-07 $X=10969 $Y=31098 $D=616
M366 24 153 vss vss hvtnfet l=6e-08 w=3e-07 $X=10969 $Y=37457 $D=616
M367 vss 156 b_pxbb_n<4> vss hvtnfet l=6e-08 w=1.285e-06 $X=10970 $Y=336 $D=616
M368 vss 157 156 vss hvtnfet l=6e-08 w=5e-07 $X=10970 $Y=6701 $D=616
M369 vss 105 157 vss hvtnfet l=6e-08 w=3e-07 $X=10970 $Y=7831 $D=616
M370 vss 105 158 vss hvtnfet l=6e-08 w=3e-07 $X=10970 $Y=43002 $D=616
M371 vss 158 159 vss hvtnfet l=6e-08 w=5e-07 $X=10970 $Y=43932 $D=616
M372 vss 159 t_pxbb_n<4> vss hvtnfet l=6e-08 w=1.285e-06 $X=10970 $Y=49512 $D=616
M373 132 ab<7> vss vss hvtnfet l=6e-08 w=2.74e-07 $X=11106 $Y=13476 $D=616
M374 153 154 vss vss hvtnfet l=6e-08 w=5e-07 $X=11106 $Y=32443 $D=616
M375 967 160 961 vss hvtnfet l=6e-08 w=5.49e-07 $X=11121 $Y=17417 $D=616
M376 968 160 962 vss hvtnfet l=6e-08 w=5.49e-07 $X=11121 $Y=18966 $D=616
M377 969 160 963 vss hvtnfet l=6e-08 w=5.49e-07 $X=11121 $Y=24337 $D=616
M378 970 160 964 vss hvtnfet l=6e-08 w=5.49e-07 $X=11121 $Y=25886 $D=616
M379 vss 155 965 vss hvtnfet l=6e-08 w=4.11e-07 $X=11126 $Y=11276 $D=616
M380 vss 155 966 vss hvtnfet l=6e-08 w=4.11e-07 $X=11126 $Y=39446 $D=616
M381 vss 153 dwlb<1> vss hvtnfet l=6e-08 w=3e-07 $X=11229 $Y=31098 $D=616
M382 vss 153 24 vss hvtnfet l=6e-08 w=3e-07 $X=11229 $Y=37457 $D=616
M383 971 121 967 vss hvtnfet l=6e-08 w=5.49e-07 $X=11381 $Y=17417 $D=616
M384 972 121 968 vss hvtnfet l=6e-08 w=5.49e-07 $X=11381 $Y=18966 $D=616
M385 973 122 969 vss hvtnfet l=6e-08 w=5.49e-07 $X=11381 $Y=24337 $D=616
M386 974 122 970 vss hvtnfet l=6e-08 w=5.49e-07 $X=11381 $Y=25886 $D=616
M387 b_pxbb_n<5> 164 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=11480 $Y=336 $D=616
M388 164 165 vss vss hvtnfet l=6e-08 w=5e-07 $X=11480 $Y=6701 $D=616
M389 165 106 vss vss hvtnfet l=6e-08 w=3e-07 $X=11480 $Y=7831 $D=616
M390 166 106 vss vss hvtnfet l=6e-08 w=3e-07 $X=11480 $Y=43002 $D=616
M391 167 166 vss vss hvtnfet l=6e-08 w=5e-07 $X=11480 $Y=43932 $D=616
M392 t_pxbb_n<5> 167 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=11480 $Y=49512 $D=616
M393 47 162 vss vss hvtnfet l=6e-08 w=2e-07 $X=11636 $Y=11276 $D=616
M394 50 163 vss vss hvtnfet l=6e-08 w=2e-07 $X=11636 $Y=39657 $D=616
M395 vss 43 971 vss hvtnfet l=6e-08 w=8.23e-07 $X=11651 $Y=17143 $D=616
M396 vss 43 972 vss hvtnfet l=6e-08 w=8.23e-07 $X=11651 $Y=18966 $D=616
M397 vss 43 973 vss hvtnfet l=6e-08 w=8.23e-07 $X=11651 $Y=24063 $D=616
M398 vss 43 974 vss hvtnfet l=6e-08 w=8.23e-07 $X=11651 $Y=25886 $D=616
M399 172 142 vss vss hvtnfet l=6e-08 w=2e-07 $X=11739 $Y=31098 $D=616
M400 vss 164 b_pxbb_n<5> vss hvtnfet l=6e-08 w=1.285e-06 $X=11740 $Y=336 $D=616
M401 vss 165 164 vss hvtnfet l=6e-08 w=5e-07 $X=11740 $Y=6701 $D=616
M402 vss 106 165 vss hvtnfet l=6e-08 w=3e-07 $X=11740 $Y=7831 $D=616
M403 vss 106 166 vss hvtnfet l=6e-08 w=3e-07 $X=11740 $Y=43002 $D=616
M404 vss 166 167 vss hvtnfet l=6e-08 w=5e-07 $X=11740 $Y=43932 $D=616
M405 vss 167 t_pxbb_n<5> vss hvtnfet l=6e-08 w=1.285e-06 $X=11740 $Y=49512 $D=616
M406 vss tm<0> dbl_pd_n<0> vss hvtnfet l=6e-08 w=2.14e-07 $X=11746 $Y=13361 $D=616
M407 dbl_pd_n<0> tm<0> vss vss hvtnfet l=6e-08 w=2.14e-07 $X=12006 $Y=13361 $D=616
M408 179 173 vss vss hvtnfet l=6e-08 w=2e-07 $X=12086 $Y=32533 $D=616
M409 vss 174 2 vss hvtnfet l=6e-08 w=2e-07 $X=12146 $Y=11276 $D=616
M410 177 168 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=12146 $Y=17812 $D=616
M411 178 169 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=12146 $Y=18983 $D=616
M412 137 170 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=12146 $Y=24732 $D=616
M413 148 171 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=12146 $Y=25903 $D=616
M414 vss 175 6 vss hvtnfet l=6e-08 w=2e-07 $X=12146 $Y=39657 $D=616
M415 975 33 168 vss hvtnfet l=6e-08 w=1.8e-07 $X=12161 $Y=17143 $D=616
M416 976 33 169 vss hvtnfet l=6e-08 w=1.8e-07 $X=12161 $Y=19609 $D=616
M417 977 33 170 vss hvtnfet l=6e-08 w=1.8e-07 $X=12161 $Y=24063 $D=616
M418 978 33 171 vss hvtnfet l=6e-08 w=1.8e-07 $X=12161 $Y=26529 $D=616
M419 vss 172 143 vss hvtnfet l=6e-08 w=6e-07 $X=12193 $Y=37037 $D=616
M420 b_pxbb_n<6> 180 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=12250 $Y=336 $D=616
M421 180 181 vss vss hvtnfet l=6e-08 w=5e-07 $X=12250 $Y=6701 $D=616
M422 181 177 vss vss hvtnfet l=6e-08 w=3e-07 $X=12250 $Y=7831 $D=616
M423 182 177 vss vss hvtnfet l=6e-08 w=3e-07 $X=12250 $Y=43002 $D=616
M424 183 182 vss vss hvtnfet l=6e-08 w=5e-07 $X=12250 $Y=43932 $D=616
M425 t_pxbb_n<6> 183 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=12250 $Y=49512 $D=616
M426 vss tm<0> dbl_pd_n<0> vss hvtnfet l=6e-08 w=2.14e-07 $X=12266 $Y=13361 $D=616
M427 vss 142 184 vss hvtnfet l=2.5e-07 w=3.5e-07 $X=12309 $Y=30853 $D=616
M428 vss 168 177 vss hvtnfet l=6e-08 w=1.37e-07 $X=12406 $Y=17812 $D=616
M429 vss 169 178 vss hvtnfet l=6e-08 w=1.37e-07 $X=12406 $Y=18983 $D=616
M430 vss 170 137 vss hvtnfet l=6e-08 w=1.37e-07 $X=12406 $Y=24732 $D=616
M431 vss 171 148 vss hvtnfet l=6e-08 w=1.37e-07 $X=12406 $Y=25903 $D=616
M432 vss 177 975 vss hvtnfet l=6e-08 w=1.8e-07 $X=12421 $Y=17143 $D=616
M433 vss 178 976 vss hvtnfet l=6e-08 w=1.8e-07 $X=12421 $Y=19609 $D=616
M434 vss 137 977 vss hvtnfet l=6e-08 w=1.8e-07 $X=12421 $Y=24063 $D=616
M435 vss 148 978 vss hvtnfet l=6e-08 w=1.8e-07 $X=12421 $Y=26529 $D=616
M436 vss 180 b_pxbb_n<6> vss hvtnfet l=6e-08 w=1.285e-06 $X=12510 $Y=336 $D=616
M437 vss 181 180 vss hvtnfet l=6e-08 w=5e-07 $X=12510 $Y=6701 $D=616
M438 vss 177 181 vss hvtnfet l=6e-08 w=3e-07 $X=12510 $Y=7831 $D=616
M439 vss 177 182 vss hvtnfet l=6e-08 w=3e-07 $X=12510 $Y=43002 $D=616
M440 vss 182 183 vss hvtnfet l=6e-08 w=5e-07 $X=12510 $Y=43932 $D=616
M441 vss 183 t_pxbb_n<6> vss hvtnfet l=6e-08 w=1.285e-06 $X=12510 $Y=49512 $D=616
M442 vss 179 186 vss hvtnfet l=6e-08 w=2e-07 $X=12596 $Y=32533 $D=616
M443 979 185 vss vss hvtnfet l=6e-08 w=4.11e-07 $X=12656 $Y=11276 $D=616
M444 980 185 vss vss hvtnfet l=6e-08 w=4.11e-07 $X=12656 $Y=39446 $D=616
M445 191 184 vss vss hvtnfet l=6e-08 w=3.5e-07 $X=12759 $Y=30853 $D=616
M446 vss 131 dbl_pd_n<2> vss hvtnfet l=6e-08 w=2.14e-07 $X=12776 $Y=13361 $D=616
M447 186 191 vss vss hvtnfet l=6e-08 w=2e-07 $X=12856 $Y=32533 $D=616
M448 174 dwlb<1> 979 vss hvtnfet l=6e-08 w=4.11e-07 $X=12916 $Y=11276 $D=616
M449 175 dwlb<0> 980 vss hvtnfet l=6e-08 w=4.11e-07 $X=12916 $Y=39446 $D=616
M450 981 187 vss vss hvtnfet l=6e-08 w=1.8e-07 $X=12931 $Y=17143 $D=616
M451 982 188 vss vss hvtnfet l=6e-08 w=1.8e-07 $X=12931 $Y=19609 $D=616
M452 983 189 vss vss hvtnfet l=6e-08 w=1.8e-07 $X=12931 $Y=24063 $D=616
M453 984 190 vss vss hvtnfet l=6e-08 w=1.8e-07 $X=12931 $Y=26529 $D=616
M454 187 192 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=12946 $Y=17812 $D=616
M455 188 193 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=12946 $Y=18983 $D=616
M456 189 194 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=12946 $Y=24732 $D=616
M457 190 195 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=12946 $Y=25903 $D=616
M458 vss 186 143 vss hvtnfet l=6e-08 w=6e-07 $X=12973 $Y=37037 $D=616
M459 b_pxbb_n<7> 196 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=13020 $Y=336 $D=616
M460 196 197 vss vss hvtnfet l=6e-08 w=5e-07 $X=13020 $Y=6701 $D=616
M461 197 178 vss vss hvtnfet l=6e-08 w=3e-07 $X=13020 $Y=7831 $D=616
M462 198 178 vss vss hvtnfet l=6e-08 w=3e-07 $X=13020 $Y=43002 $D=616
M463 199 198 vss vss hvtnfet l=6e-08 w=5e-07 $X=13020 $Y=43932 $D=616
M464 t_pxbb_n<7> 199 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=13020 $Y=49512 $D=616
M465 dbl_pd_n<2> 131 vss vss hvtnfet l=6e-08 w=2.14e-07 $X=13036 $Y=13361 $D=616
M466 192 33 981 vss hvtnfet l=6e-08 w=1.8e-07 $X=13191 $Y=17143 $D=616
M467 193 33 982 vss hvtnfet l=6e-08 w=1.8e-07 $X=13191 $Y=19609 $D=616
M468 194 33 983 vss hvtnfet l=6e-08 w=1.8e-07 $X=13191 $Y=24063 $D=616
M469 195 33 984 vss hvtnfet l=6e-08 w=1.8e-07 $X=13191 $Y=26529 $D=616
M470 vss 192 187 vss hvtnfet l=6e-08 w=1.37e-07 $X=13206 $Y=17812 $D=616
M471 vss 193 188 vss hvtnfet l=6e-08 w=1.37e-07 $X=13206 $Y=18983 $D=616
M472 vss 194 189 vss hvtnfet l=6e-08 w=1.37e-07 $X=13206 $Y=24732 $D=616
M473 vss 195 190 vss hvtnfet l=6e-08 w=1.37e-07 $X=13206 $Y=25903 $D=616
M474 vss 196 b_pxbb_n<7> vss hvtnfet l=6e-08 w=1.285e-06 $X=13280 $Y=336 $D=616
M475 vss 197 196 vss hvtnfet l=6e-08 w=5e-07 $X=13280 $Y=6701 $D=616
M476 vss 178 197 vss hvtnfet l=6e-08 w=3e-07 $X=13280 $Y=7831 $D=616
M477 vss 178 198 vss hvtnfet l=6e-08 w=3e-07 $X=13280 $Y=43002 $D=616
M478 vss 198 199 vss hvtnfet l=6e-08 w=5e-07 $X=13280 $Y=43932 $D=616
M479 vss 199 t_pxbb_n<7> vss hvtnfet l=6e-08 w=1.285e-06 $X=13280 $Y=49512 $D=616
M480 vss 131 dbl_pd_n<2> vss hvtnfet l=6e-08 w=2.14e-07 $X=13296 $Y=13361 $D=616
M481 vss 191 202 vss hvtnfet l=2.5e-07 w=3.5e-07 $X=13429 $Y=30853 $D=616
M482 vss tm<7> 203 vss hvtnfet l=6e-08 w=2e-07 $X=13432 $Y=32533 $D=616
M483 985 43 vss vss hvtnfet l=6e-08 w=8.23e-07 $X=13701 $Y=17143 $D=616
M484 986 43 vss vss hvtnfet l=6e-08 w=8.23e-07 $X=13701 $Y=18966 $D=616
M485 987 43 vss vss hvtnfet l=6e-08 w=8.23e-07 $X=13701 $Y=24063 $D=616
M486 988 43 vss vss hvtnfet l=6e-08 w=8.23e-07 $X=13701 $Y=25886 $D=616
M487 vss 200 143 vss hvtnfet l=6e-08 w=6e-07 $X=13753 $Y=37037 $D=616
M488 b_pxcb_n<0> 206 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=13790 $Y=336 $D=616
M489 206 207 vss vss hvtnfet l=6e-08 w=5e-07 $X=13790 $Y=6701 $D=616
M490 207 189 vss vss hvtnfet l=6e-08 w=3e-07 $X=13790 $Y=7831 $D=616
M491 208 189 vss vss hvtnfet l=6e-08 w=3e-07 $X=13790 $Y=43002 $D=616
M492 209 208 vss vss hvtnfet l=6e-08 w=5e-07 $X=13790 $Y=43932 $D=616
M493 t_pxcb_n<0> 209 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=13790 $Y=49512 $D=616
M494 211 202 vss vss hvtnfet l=6e-08 w=3.5e-07 $X=13879 $Y=30853 $D=616
M495 vss 205 204 vss hvtnfet l=6e-08 w=2.74e-07 $X=13936 $Y=13476 $D=616
M496 vss 203 200 vss hvtnfet l=6e-08 w=2e-07 $X=13942 $Y=32533 $D=616
M497 989 204 985 vss hvtnfet l=6e-08 w=5.49e-07 $X=13971 $Y=17417 $D=616
M498 990 204 986 vss hvtnfet l=6e-08 w=5.49e-07 $X=13971 $Y=18966 $D=616
M499 991 205 987 vss hvtnfet l=6e-08 w=5.49e-07 $X=13971 $Y=24337 $D=616
M500 992 205 988 vss hvtnfet l=6e-08 w=5.49e-07 $X=13971 $Y=25886 $D=616
M501 vss 206 b_pxcb_n<0> vss hvtnfet l=6e-08 w=1.285e-06 $X=14050 $Y=336 $D=616
M502 vss 207 206 vss hvtnfet l=6e-08 w=5e-07 $X=14050 $Y=6701 $D=616
M503 vss 189 207 vss hvtnfet l=6e-08 w=3e-07 $X=14050 $Y=7831 $D=616
M504 vss 189 208 vss hvtnfet l=6e-08 w=3e-07 $X=14050 $Y=43002 $D=616
M505 vss 208 209 vss hvtnfet l=6e-08 w=5e-07 $X=14050 $Y=43932 $D=616
M506 vss 209 t_pxcb_n<0> vss hvtnfet l=6e-08 w=1.285e-06 $X=14050 $Y=49512 $D=616
M507 200 211 vss vss hvtnfet l=6e-08 w=2e-07 $X=14202 $Y=32533 $D=616
M508 993 dwlb<1> 216 vss hvtnfet l=6e-08 w=4.11e-07 $X=14216 $Y=11276 $D=616
M509 994 dwlb<0> 217 vss hvtnfet l=6e-08 w=4.11e-07 $X=14216 $Y=39446 $D=616
M510 995 210 989 vss hvtnfet l=6e-08 w=5.49e-07 $X=14231 $Y=17417 $D=616
M511 996 210 990 vss hvtnfet l=6e-08 w=5.49e-07 $X=14231 $Y=18966 $D=616
M512 997 210 991 vss hvtnfet l=6e-08 w=5.49e-07 $X=14231 $Y=24337 $D=616
M513 998 210 992 vss hvtnfet l=6e-08 w=5.49e-07 $X=14231 $Y=25886 $D=616
M514 205 ab<12> vss vss hvtnfet l=6e-08 w=2.74e-07 $X=14446 $Y=13476 $D=616
M515 vss 212 993 vss hvtnfet l=6e-08 w=4.11e-07 $X=14476 $Y=11276 $D=616
M516 vss 212 994 vss hvtnfet l=6e-08 w=4.11e-07 $X=14476 $Y=39446 $D=616
M517 192 213 995 vss hvtnfet l=6e-08 w=5.49e-07 $X=14491 $Y=17417 $D=616
M518 193 214 996 vss hvtnfet l=6e-08 w=5.49e-07 $X=14491 $Y=18966 $D=616
M519 194 213 997 vss hvtnfet l=6e-08 w=5.49e-07 $X=14491 $Y=24337 $D=616
M520 195 214 998 vss hvtnfet l=6e-08 w=5.49e-07 $X=14491 $Y=25886 $D=616
M521 b_pxcb_n<1> 218 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=14560 $Y=336 $D=616
M522 218 219 vss vss hvtnfet l=6e-08 w=5e-07 $X=14560 $Y=6701 $D=616
M523 219 190 vss vss hvtnfet l=6e-08 w=3e-07 $X=14560 $Y=7831 $D=616
M524 220 190 vss vss hvtnfet l=6e-08 w=3e-07 $X=14560 $Y=43002 $D=616
M525 221 220 vss vss hvtnfet l=6e-08 w=5e-07 $X=14560 $Y=43932 $D=616
M526 t_pxcb_n<1> 221 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=14560 $Y=49512 $D=616
M527 vss 123 624 vss hvtnfet l=6e-08 w=6e-07 $X=14796 $Y=30668 $D=616
M528 vss 218 b_pxcb_n<1> vss hvtnfet l=6e-08 w=1.285e-06 $X=14820 $Y=336 $D=616
M529 vss 219 218 vss hvtnfet l=6e-08 w=5e-07 $X=14820 $Y=6701 $D=616
M530 vss 190 219 vss hvtnfet l=6e-08 w=3e-07 $X=14820 $Y=7831 $D=616
M531 vss 190 220 vss hvtnfet l=6e-08 w=3e-07 $X=14820 $Y=43002 $D=616
M532 vss 220 221 vss hvtnfet l=6e-08 w=5e-07 $X=14820 $Y=43932 $D=616
M533 vss 221 t_pxcb_n<1> vss hvtnfet l=6e-08 w=1.285e-06 $X=14820 $Y=49512 $D=616
M534 vss 72 58 vss hvtnfet l=6e-08 w=2e-07 $X=14872 $Y=37045 $D=616
M535 48 216 vss vss hvtnfet l=6e-08 w=2e-07 $X=14986 $Y=11276 $D=616
M536 49 217 vss vss hvtnfet l=6e-08 w=2e-07 $X=14986 $Y=39657 $D=616
M537 vss 43 33 vss hvtnfet l=6e-08 w=7e-07 $X=15316 $Y=30668 $D=616
M538 b_pxcb_n<2> 223 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=15330 $Y=336 $D=616
M539 223 224 vss vss hvtnfet l=6e-08 w=5e-07 $X=15330 $Y=6701 $D=616
M540 224 225 vss vss hvtnfet l=6e-08 w=3e-07 $X=15330 $Y=7831 $D=616
M541 226 225 vss vss hvtnfet l=6e-08 w=3e-07 $X=15330 $Y=43002 $D=616
M542 227 226 vss vss hvtnfet l=6e-08 w=5e-07 $X=15330 $Y=43932 $D=616
M543 t_pxcb_n<2> 227 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=15330 $Y=49512 $D=616
M544 629 229 vss vss hvtnfet l=6e-08 w=4e-07 $X=15382 $Y=37045 $D=616
M545 vss ab<11> 210 vss hvtnfet l=6e-08 w=2.74e-07 $X=15456 $Y=13476 $D=616
M546 33 43 vss vss hvtnfet l=6e-08 w=7e-07 $X=15576 $Y=30668 $D=616
M547 vss 223 b_pxcb_n<2> vss hvtnfet l=6e-08 w=1.285e-06 $X=15590 $Y=336 $D=616
M548 vss 224 223 vss hvtnfet l=6e-08 w=5e-07 $X=15590 $Y=6701 $D=616
M549 vss 225 224 vss hvtnfet l=6e-08 w=3e-07 $X=15590 $Y=7831 $D=616
M550 vss 225 226 vss hvtnfet l=6e-08 w=3e-07 $X=15590 $Y=43002 $D=616
M551 vss 226 227 vss hvtnfet l=6e-08 w=5e-07 $X=15590 $Y=43932 $D=616
M552 vss 227 t_pxcb_n<2> vss hvtnfet l=6e-08 w=1.285e-06 $X=15590 $Y=49512 $D=616
M553 vss 228 231 vss hvtnfet l=6e-08 w=2.1e-07 $X=15621 $Y=32688 $D=616
M554 72 172 629 vss hvtnfet l=6e-08 w=4e-07 $X=15642 $Y=37045 $D=616
M555 240 210 vss vss hvtnfet l=6e-08 w=2.74e-07 $X=15716 $Y=13476 $D=616
M556 631 tm<0> vss vss hvtnfet l=6e-08 w=2.74e-07 $X=15880 $Y=39358 $D=616
M557 630 131 vss vss hvtnfet l=6e-08 w=2.1e-07 $X=15881 $Y=32688 $D=616
M558 vss tm<3> 242 vss hvtnfet l=7e-08 w=3.2e-07 $X=16057 $Y=11276 $D=616
M559 b_pxcb_n<3> 235 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=16100 $Y=336 $D=616
M560 235 236 vss vss hvtnfet l=6e-08 w=5e-07 $X=16100 $Y=6701 $D=616
M561 236 237 vss vss hvtnfet l=6e-08 w=3e-07 $X=16100 $Y=7831 $D=616
M562 238 237 vss vss hvtnfet l=6e-08 w=3e-07 $X=16100 $Y=43002 $D=616
M563 239 238 vss vss hvtnfet l=6e-08 w=5e-07 $X=16100 $Y=43932 $D=616
M564 t_pxcb_n<3> 239 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=16100 $Y=49512 $D=616
M565 228 231 630 vss hvtnfet l=6e-08 w=2.1e-07 $X=16141 $Y=32688 $D=616
M566 vss 213 214 vss hvtnfet l=6e-08 w=2.74e-07 $X=16316 $Y=13476 $D=616
M567 635 232 vss vss hvtnfet l=6e-08 w=3.2e-07 $X=16322 $Y=37277 $D=616
M568 243 tm<4> vss vss hvtnfet l=7e-08 w=3.2e-07 $X=16327 $Y=11276 $D=616
M569 999 213 249 vss hvtnfet l=6e-08 w=5.49e-07 $X=16331 $Y=17417 $D=616
M570 1000 214 250 vss hvtnfet l=6e-08 w=5.49e-07 $X=16331 $Y=18966 $D=616
M571 1001 213 251 vss hvtnfet l=6e-08 w=5.49e-07 $X=16331 $Y=24337 $D=616
M572 1002 214 252 vss hvtnfet l=6e-08 w=5.49e-07 $X=16331 $Y=25886 $D=616
M573 vss 123 644 vss hvtnfet l=6e-08 w=6e-07 $X=16346 $Y=30668 $D=616
M574 vss 235 b_pxcb_n<3> vss hvtnfet l=6e-08 w=1.285e-06 $X=16360 $Y=336 $D=616
M575 vss 236 235 vss hvtnfet l=6e-08 w=5e-07 $X=16360 $Y=6701 $D=616
M576 vss 237 236 vss hvtnfet l=6e-08 w=3e-07 $X=16360 $Y=7831 $D=616
M577 vss 237 238 vss hvtnfet l=6e-08 w=3e-07 $X=16360 $Y=43002 $D=616
M578 vss 238 239 vss hvtnfet l=6e-08 w=5e-07 $X=16360 $Y=43932 $D=616
M579 vss 239 t_pxcb_n<3> vss hvtnfet l=6e-08 w=1.285e-06 $X=16360 $Y=49512 $D=616
M580 636 123 228 vss hvtnfet l=6e-08 w=3.2e-07 $X=16401 $Y=32578 $D=616
M581 213 ab<10> vss vss hvtnfet l=6e-08 w=2.74e-07 $X=16576 $Y=13476 $D=616
M582 229 142 635 vss hvtnfet l=6e-08 w=3.2e-07 $X=16582 $Y=37277 $D=616
M583 1003 240 999 vss hvtnfet l=6e-08 w=5.49e-07 $X=16591 $Y=17417 $D=616
M584 1004 240 1000 vss hvtnfet l=6e-08 w=5.49e-07 $X=16591 $Y=18966 $D=616
M585 1005 240 1001 vss hvtnfet l=6e-08 w=5.49e-07 $X=16591 $Y=24337 $D=616
M586 1006 240 1002 vss hvtnfet l=6e-08 w=5.49e-07 $X=16591 $Y=25886 $D=616
M587 644 123 vss vss hvtnfet l=6e-08 w=6e-07 $X=16606 $Y=30668 $D=616
M588 vss 123 636 vss hvtnfet l=6e-08 w=3.2e-07 $X=16661 $Y=32578 $D=616
M589 637 tm<6> vss vss hvtnfet l=6e-08 w=2.74e-07 $X=16680 $Y=39358 $D=616
M590 638 244 229 vss hvtnfet l=6e-08 w=2.1e-07 $X=16842 $Y=37277 $D=616
M591 vss 243 643 vss hvtnfet l=6e-08 w=4.8e-07 $X=16847 $Y=11276 $D=616
M592 1007 204 1003 vss hvtnfet l=6e-08 w=5.49e-07 $X=16851 $Y=17417 $D=616
M593 1008 204 1004 vss hvtnfet l=6e-08 w=5.49e-07 $X=16851 $Y=18966 $D=616
M594 1009 205 1005 vss hvtnfet l=6e-08 w=5.49e-07 $X=16851 $Y=24337 $D=616
M595 1010 205 1006 vss hvtnfet l=6e-08 w=5.49e-07 $X=16851 $Y=25886 $D=616
M596 642 123 644 vss hvtnfet l=6e-08 w=6e-07 $X=16866 $Y=30668 $D=616
M597 b_pxcb_n<4> 245 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=16870 $Y=336 $D=616
M598 245 246 vss vss hvtnfet l=6e-08 w=5e-07 $X=16870 $Y=6701 $D=616
M599 246 187 vss vss hvtnfet l=6e-08 w=3e-07 $X=16870 $Y=7831 $D=616
M600 247 187 vss vss hvtnfet l=6e-08 w=3e-07 $X=16870 $Y=43002 $D=616
M601 248 247 vss vss hvtnfet l=6e-08 w=5e-07 $X=16870 $Y=43932 $D=616
M602 t_pxcb_n<4> 248 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=16870 $Y=49512 $D=616
M603 vss 172 638 vss hvtnfet l=6e-08 w=2.1e-07 $X=17102 $Y=37277 $D=616
M604 643 242 vss vss hvtnfet l=6e-08 w=4.8e-07 $X=17107 $Y=11276 $D=616
M605 vss 43 1007 vss hvtnfet l=6e-08 w=8.23e-07 $X=17121 $Y=17143 $D=616
M606 vss 43 1008 vss hvtnfet l=6e-08 w=8.23e-07 $X=17121 $Y=18966 $D=616
M607 vss 43 1009 vss hvtnfet l=6e-08 w=8.23e-07 $X=17121 $Y=24063 $D=616
M608 vss 43 1010 vss hvtnfet l=6e-08 w=8.23e-07 $X=17121 $Y=25886 $D=616
M609 644 123 642 vss hvtnfet l=6e-08 w=6e-07 $X=17126 $Y=30668 $D=616
M610 vss 245 b_pxcb_n<4> vss hvtnfet l=6e-08 w=1.285e-06 $X=17130 $Y=336 $D=616
M611 vss 246 245 vss hvtnfet l=6e-08 w=5e-07 $X=17130 $Y=6701 $D=616
M612 vss 187 246 vss hvtnfet l=6e-08 w=3e-07 $X=17130 $Y=7831 $D=616
M613 vss 187 247 vss hvtnfet l=6e-08 w=3e-07 $X=17130 $Y=43002 $D=616
M614 vss 247 248 vss hvtnfet l=6e-08 w=5e-07 $X=17130 $Y=43932 $D=616
M615 vss 248 t_pxcb_n<4> vss hvtnfet l=6e-08 w=1.285e-06 $X=17130 $Y=49512 $D=616
M616 244 229 vss vss hvtnfet l=6e-08 w=2.1e-07 $X=17362 $Y=37277 $D=616
M617 253 249 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=17616 $Y=17812 $D=616
M618 254 250 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=17616 $Y=18983 $D=616
M619 225 251 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=17616 $Y=24732 $D=616
M620 237 252 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=17616 $Y=25903 $D=616
M621 647 242 vss vss hvtnfet l=6e-08 w=4.8e-07 $X=17617 $Y=11276 $D=616
M622 1011 33 249 vss hvtnfet l=6e-08 w=1.8e-07 $X=17631 $Y=17143 $D=616
M623 1012 33 250 vss hvtnfet l=6e-08 w=1.8e-07 $X=17631 $Y=19609 $D=616
M624 1013 33 251 vss hvtnfet l=6e-08 w=1.8e-07 $X=17631 $Y=24063 $D=616
M625 1014 33 252 vss hvtnfet l=6e-08 w=1.8e-07 $X=17631 $Y=26529 $D=616
M626 b_pxcb_n<5> 255 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=17640 $Y=336 $D=616
M627 255 256 vss vss hvtnfet l=6e-08 w=5e-07 $X=17640 $Y=6701 $D=616
M628 256 188 vss vss hvtnfet l=6e-08 w=3e-07 $X=17640 $Y=7831 $D=616
M629 257 188 vss vss hvtnfet l=6e-08 w=3e-07 $X=17640 $Y=43002 $D=616
M630 258 257 vss vss hvtnfet l=6e-08 w=5e-07 $X=17640 $Y=43932 $D=616
M631 t_pxcb_n<5> 258 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=17640 $Y=49512 $D=616
M632 23 clkb vss vss hvtnfet l=6e-08 w=4.5e-07 $X=17646 $Y=30668 $D=616
M633 vss 249 253 vss hvtnfet l=6e-08 w=1.37e-07 $X=17876 $Y=17812 $D=616
M634 vss 250 254 vss hvtnfet l=6e-08 w=1.37e-07 $X=17876 $Y=18983 $D=616
M635 vss 251 225 vss hvtnfet l=6e-08 w=1.37e-07 $X=17876 $Y=24732 $D=616
M636 vss 252 237 vss hvtnfet l=6e-08 w=1.37e-07 $X=17876 $Y=25903 $D=616
M637 vss tm<4> 647 vss hvtnfet l=6e-08 w=4.8e-07 $X=17877 $Y=11276 $D=616
M638 vss 253 1011 vss hvtnfet l=6e-08 w=1.8e-07 $X=17891 $Y=17143 $D=616
M639 vss 254 1012 vss hvtnfet l=6e-08 w=1.8e-07 $X=17891 $Y=19609 $D=616
M640 vss 225 1013 vss hvtnfet l=6e-08 w=1.8e-07 $X=17891 $Y=24063 $D=616
M641 vss 237 1014 vss hvtnfet l=6e-08 w=1.8e-07 $X=17891 $Y=26529 $D=616
M642 vss 255 b_pxcb_n<5> vss hvtnfet l=6e-08 w=1.285e-06 $X=17900 $Y=336 $D=616
M643 vss 256 255 vss hvtnfet l=6e-08 w=5e-07 $X=17900 $Y=6701 $D=616
M644 vss 188 256 vss hvtnfet l=6e-08 w=3e-07 $X=17900 $Y=7831 $D=616
M645 vss 188 257 vss hvtnfet l=6e-08 w=3e-07 $X=17900 $Y=43002 $D=616
M646 vss 257 258 vss hvtnfet l=6e-08 w=5e-07 $X=17900 $Y=43932 $D=616
M647 vss 258 t_pxcb_n<5> vss hvtnfet l=6e-08 w=1.285e-06 $X=17900 $Y=49512 $D=616
M648 vss 260 273 vss hvtnfet l=6e-08 w=2.74e-07 $X=18106 $Y=13476 $D=616
M649 vss wenb 232 vss hvtnfet l=6e-08 w=2e-07 $X=18366 $Y=37147 $D=616
M650 648 tm<4> vss vss hvtnfet l=6e-08 w=4.8e-07 $X=18387 $Y=11276 $D=616
M651 b_pxcb_n<6> 265 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=18410 $Y=336 $D=616
M652 265 266 vss vss hvtnfet l=6e-08 w=5e-07 $X=18410 $Y=6701 $D=616
M653 266 253 vss vss hvtnfet l=6e-08 w=3e-07 $X=18410 $Y=7831 $D=616
M654 267 253 vss vss hvtnfet l=6e-08 w=3e-07 $X=18410 $Y=43002 $D=616
M655 268 267 vss vss hvtnfet l=6e-08 w=5e-07 $X=18410 $Y=43932 $D=616
M656 t_pxcb_n<6> 268 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=18410 $Y=49512 $D=616
M657 651 ab<4> vss vss hvtnfet l=6e-08 w=3.2e-07 $X=18460 $Y=30918 $D=616
M658 652 wenb vss vss hvtnfet l=6e-08 w=3.2e-07 $X=18460 $Y=32578 $D=616
M659 vss tm<2> 173 vss hvtnfet l=6e-08 w=2.74e-07 $X=18510 $Y=39358 $D=616
M660 260 ab<1> vss vss hvtnfet l=6e-08 w=2.74e-07 $X=18616 $Y=13476 $D=616
M661 232 264 vss vss hvtnfet l=6e-08 w=2e-07 $X=18626 $Y=37147 $D=616
M662 vss tm<3> 648 vss hvtnfet l=6e-08 w=4.8e-07 $X=18647 $Y=11276 $D=616
M663 vss 265 b_pxcb_n<6> vss hvtnfet l=6e-08 w=1.285e-06 $X=18670 $Y=336 $D=616
M664 vss 266 265 vss hvtnfet l=6e-08 w=5e-07 $X=18670 $Y=6701 $D=616
M665 vss 253 266 vss hvtnfet l=6e-08 w=3e-07 $X=18670 $Y=7831 $D=616
M666 vss 253 267 vss hvtnfet l=6e-08 w=3e-07 $X=18670 $Y=43002 $D=616
M667 vss 267 268 vss hvtnfet l=6e-08 w=5e-07 $X=18670 $Y=43932 $D=616
M668 vss 268 t_pxcb_n<6> vss hvtnfet l=6e-08 w=1.285e-06 $X=18670 $Y=49512 $D=616
M669 154 23 651 vss hvtnfet l=6e-08 w=3.2e-07 $X=18720 $Y=30918 $D=616
M670 274 23 652 vss hvtnfet l=6e-08 w=3.2e-07 $X=18720 $Y=32578 $D=616
M671 1015 269 280 vss hvtnfet l=6e-08 w=5.49e-07 $X=18911 $Y=17143 $D=616
M672 1016 270 281 vss hvtnfet l=6e-08 w=5.49e-07 $X=18911 $Y=19240 $D=616
M673 1017 269 282 vss hvtnfet l=6e-08 w=5.49e-07 $X=18911 $Y=24063 $D=616
M674 1018 270 283 vss hvtnfet l=6e-08 w=5.49e-07 $X=18911 $Y=26160 $D=616
M675 653 271 154 vss hvtnfet l=6e-08 w=2.1e-07 $X=18980 $Y=30918 $D=616
M676 654 272 274 vss hvtnfet l=6e-08 w=2.1e-07 $X=18980 $Y=32688 $D=616
M677 vss 270 269 vss hvtnfet l=6e-08 w=2.74e-07 $X=19126 $Y=13476 $D=616
M678 659 tm<3> vss vss hvtnfet l=6e-08 w=4.8e-07 $X=19157 $Y=11276 $D=616
M679 1019 273 1015 vss hvtnfet l=6e-08 w=5.49e-07 $X=19171 $Y=17143 $D=616
M680 1020 273 1016 vss hvtnfet l=6e-08 w=5.49e-07 $X=19171 $Y=19240 $D=616
M681 1021 260 1017 vss hvtnfet l=6e-08 w=5.49e-07 $X=19171 $Y=24063 $D=616
M682 1022 260 1018 vss hvtnfet l=6e-08 w=5.49e-07 $X=19171 $Y=26160 $D=616
M683 b_pxcb_n<7> 275 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=19180 $Y=336 $D=616
M684 275 276 vss vss hvtnfet l=6e-08 w=5e-07 $X=19180 $Y=6701 $D=616
M685 276 254 vss vss hvtnfet l=6e-08 w=3e-07 $X=19180 $Y=7831 $D=616
M686 277 254 vss vss hvtnfet l=6e-08 w=3e-07 $X=19180 $Y=43002 $D=616
M687 278 277 vss vss hvtnfet l=6e-08 w=5e-07 $X=19180 $Y=43932 $D=616
M688 t_pxcb_n<7> 278 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=19180 $Y=49512 $D=616
M689 vss clkb 653 vss hvtnfet l=6e-08 w=2.1e-07 $X=19240 $Y=30918 $D=616
M690 vss clkb 654 vss hvtnfet l=6e-08 w=2.1e-07 $X=19240 $Y=32688 $D=616
M691 vss 243 659 vss hvtnfet l=6e-08 w=4.8e-07 $X=19417 $Y=11276 $D=616
M692 vss 275 b_pxcb_n<7> vss hvtnfet l=6e-08 w=1.285e-06 $X=19440 $Y=336 $D=616
M693 vss 276 275 vss hvtnfet l=6e-08 w=5e-07 $X=19440 $Y=6701 $D=616
M694 vss 254 276 vss hvtnfet l=6e-08 w=3e-07 $X=19440 $Y=7831 $D=616
M695 vss 254 277 vss hvtnfet l=6e-08 w=3e-07 $X=19440 $Y=43002 $D=616
M696 vss 277 278 vss hvtnfet l=6e-08 w=5e-07 $X=19440 $Y=43932 $D=616
M697 vss 278 t_pxcb_n<7> vss hvtnfet l=6e-08 w=1.285e-06 $X=19440 $Y=49512 $D=616
M698 vss 43 1019 vss hvtnfet l=6e-08 w=8.23e-07 $X=19441 $Y=17143 $D=616
M699 vss 43 1020 vss hvtnfet l=6e-08 w=8.23e-07 $X=19441 $Y=18966 $D=616
M700 vss 43 1021 vss hvtnfet l=6e-08 w=8.23e-07 $X=19441 $Y=24063 $D=616
M701 vss 43 1022 vss hvtnfet l=6e-08 w=8.23e-07 $X=19441 $Y=25886 $D=616
M702 271 154 vss vss hvtnfet l=6e-08 w=2.1e-07 $X=19500 $Y=30918 $D=616
M703 272 274 vss vss hvtnfet l=6e-08 w=2.1e-07 $X=19500 $Y=32688 $D=616
M704 270 ab<0> vss vss hvtnfet l=6e-08 w=2.74e-07 $X=19636 $Y=13476 $D=616
M705 vss 15 r_saeb_n vss hvtnfet l=6e-08 w=8.58e-07 $X=19675 $Y=37027 $D=616
M706 r_saeb_n 15 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=19935 $Y=37027 $D=616
M707 1023 33 280 vss hvtnfet l=6e-08 w=1.8e-07 $X=19951 $Y=17143 $D=616
M708 212 280 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=19951 $Y=17812 $D=616
M709 185 281 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=19951 $Y=18983 $D=616
M710 1024 33 281 vss hvtnfet l=6e-08 w=1.8e-07 $X=19951 $Y=19609 $D=616
M711 1025 33 282 vss hvtnfet l=6e-08 w=1.8e-07 $X=19951 $Y=24063 $D=616
M712 155 282 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=19951 $Y=24732 $D=616
M713 145 283 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=19951 $Y=25903 $D=616
M714 1026 33 283 vss hvtnfet l=6e-08 w=1.8e-07 $X=19951 $Y=26529 $D=616
M715 vss 11 rb_cb<0> vss hvtnfet l=6e-08 w=8.58e-07 $X=20195 $Y=328 $D=616
M716 vss 12 rb_cb<2> vss hvtnfet l=6e-08 w=8.58e-07 $X=20195 $Y=5316 $D=616
M717 vss 13 rb_mb<0> vss hvtnfet l=6e-08 w=8.58e-07 $X=20195 $Y=6788 $D=616
M718 vss 14 rb_mb<2> vss hvtnfet l=6e-08 w=8.58e-07 $X=20195 $Y=11776 $D=616
M719 vss 15 r_saeb_n vss hvtnfet l=6e-08 w=8.58e-07 $X=20195 $Y=37027 $D=616
M720 vss 16 rt_mb<2> vss hvtnfet l=6e-08 w=8.58e-07 $X=20195 $Y=38499 $D=616
M721 vss 17 rt_mb<0> vss hvtnfet l=6e-08 w=8.58e-07 $X=20195 $Y=43487 $D=616
M722 vss 18 rt_cb<2> vss hvtnfet l=6e-08 w=8.58e-07 $X=20195 $Y=44959 $D=616
M723 vss 19 rt_cb<0> vss hvtnfet l=6e-08 w=8.58e-07 $X=20195 $Y=49947 $D=616
M724 vss 212 1023 vss hvtnfet l=6e-08 w=1.8e-07 $X=20211 $Y=17143 $D=616
M725 vss 280 212 vss hvtnfet l=6e-08 w=1.37e-07 $X=20211 $Y=17812 $D=616
M726 vss 281 185 vss hvtnfet l=6e-08 w=1.37e-07 $X=20211 $Y=18983 $D=616
M727 vss 185 1024 vss hvtnfet l=6e-08 w=1.8e-07 $X=20211 $Y=19609 $D=616
M728 vss 155 1025 vss hvtnfet l=6e-08 w=1.8e-07 $X=20211 $Y=24063 $D=616
M729 vss 282 155 vss hvtnfet l=6e-08 w=1.37e-07 $X=20211 $Y=24732 $D=616
M730 vss 283 145 vss hvtnfet l=6e-08 w=1.37e-07 $X=20211 $Y=25903 $D=616
M731 vss 145 1026 vss hvtnfet l=6e-08 w=1.8e-07 $X=20211 $Y=26529 $D=616
M732 rb_cb<0> 11 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=20455 $Y=328 $D=616
M733 rb_cb<2> 12 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=20455 $Y=5316 $D=616
M734 rb_mb<0> 13 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=20455 $Y=6788 $D=616
M735 rb_mb<2> 14 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=20455 $Y=11776 $D=616
M736 r_saeb_n 15 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=20455 $Y=37027 $D=616
M737 rt_mb<2> 16 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=20455 $Y=38499 $D=616
M738 rt_mb<0> 17 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=20455 $Y=43487 $D=616
M739 rt_cb<2> 18 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=20455 $Y=44959 $D=616
M740 rt_cb<0> 19 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=20455 $Y=49947 $D=616
M741 vss 11 rb_cb<0> vss hvtnfet l=6e-08 w=8.58e-07 $X=20715 $Y=328 $D=616
M742 vss 12 rb_cb<2> vss hvtnfet l=6e-08 w=8.58e-07 $X=20715 $Y=5316 $D=616
M743 vss 13 rb_mb<0> vss hvtnfet l=6e-08 w=8.58e-07 $X=20715 $Y=6788 $D=616
M744 vss 14 rb_mb<2> vss hvtnfet l=6e-08 w=8.58e-07 $X=20715 $Y=11776 $D=616
M745 vss 15 r_saeb_n vss hvtnfet l=6e-08 w=8.58e-07 $X=20715 $Y=37027 $D=616
M746 vss 16 rt_mb<2> vss hvtnfet l=6e-08 w=8.58e-07 $X=20715 $Y=38499 $D=616
M747 vss 17 rt_mb<0> vss hvtnfet l=6e-08 w=8.58e-07 $X=20715 $Y=43487 $D=616
M748 vss 18 rt_cb<2> vss hvtnfet l=6e-08 w=8.58e-07 $X=20715 $Y=44959 $D=616
M749 vss 19 rt_cb<0> vss hvtnfet l=6e-08 w=8.58e-07 $X=20715 $Y=49947 $D=616
M750 10 274 vss vss hvtnfet l=6e-08 w=6e-07 $X=20725 $Y=30899 $D=616
M751 rb_cb<1> 34 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=20975 $Y=328 $D=616
M752 rb_cb<3> 35 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=20975 $Y=5316 $D=616
M753 rb_mb<1> 36 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=20975 $Y=6788 $D=616
M754 rb_mb<3> 37 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=20975 $Y=11776 $D=616
M755 r_clk_dqb 8 vss vss hvtnfet l=6e-08 w=1.26e-06 $X=20975 $Y=22041 $D=616
M756 r_clk_dqb_n 9 vss vss hvtnfet l=6e-08 w=1.26e-06 $X=20975 $Y=29007 $D=616
M757 r_sa_preb_n 51 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=20975 $Y=37027 $D=616
M758 rt_mb<3> 39 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=20975 $Y=38499 $D=616
M759 rt_mb<1> 40 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=20975 $Y=43487 $D=616
M760 rt_cb<3> 41 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=20975 $Y=44959 $D=616
M761 rt_cb<1> 42 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=20975 $Y=49947 $D=616
M762 vss 34 rb_cb<1> vss hvtnfet l=6e-08 w=8.58e-07 $X=21235 $Y=328 $D=616
M763 vss 35 rb_cb<3> vss hvtnfet l=6e-08 w=8.58e-07 $X=21235 $Y=5316 $D=616
M764 vss 36 rb_mb<1> vss hvtnfet l=6e-08 w=8.58e-07 $X=21235 $Y=6788 $D=616
M765 vss 37 rb_mb<3> vss hvtnfet l=6e-08 w=8.58e-07 $X=21235 $Y=11776 $D=616
M766 rb_tm_preb_n 20 vss vss hvtnfet l=6e-08 w=1.287e-06 $X=21235 $Y=13280 $D=616
M767 rt_tm_preb_n 21 vss vss hvtnfet l=6e-08 w=1.287e-06 $X=21235 $Y=20124 $D=616
M768 vss 8 r_clk_dqb vss hvtnfet l=6e-08 w=1.26e-06 $X=21235 $Y=22041 $D=616
M769 vss 9 r_clk_dqb_n vss hvtnfet l=6e-08 w=1.26e-06 $X=21235 $Y=29007 $D=616
M770 r_lweb 10 vss vss hvtnfet l=6e-08 w=1.287e-06 $X=21235 $Y=30897 $D=616
M771 vss 51 r_sa_preb_n vss hvtnfet l=6e-08 w=8.58e-07 $X=21235 $Y=37027 $D=616
M772 vss 39 rt_mb<3> vss hvtnfet l=6e-08 w=8.58e-07 $X=21235 $Y=38499 $D=616
M773 vss 40 rt_mb<1> vss hvtnfet l=6e-08 w=8.58e-07 $X=21235 $Y=43487 $D=616
M774 vss 41 rt_cb<3> vss hvtnfet l=6e-08 w=8.58e-07 $X=21235 $Y=44959 $D=616
M775 vss 42 rt_cb<1> vss hvtnfet l=6e-08 w=8.58e-07 $X=21235 $Y=49947 $D=616
M776 rb_cb<1> 34 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=21495 $Y=328 $D=616
M777 rb_cb<3> 35 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=21495 $Y=5316 $D=616
M778 rb_mb<1> 36 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=21495 $Y=6788 $D=616
M779 rb_mb<3> 37 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=21495 $Y=11776 $D=616
M780 vss 20 rb_tm_preb_n vss hvtnfet l=6e-08 w=1.287e-06 $X=21495 $Y=13280 $D=616
M781 vss 21 rt_tm_preb_n vss hvtnfet l=6e-08 w=1.287e-06 $X=21495 $Y=20124 $D=616
M782 r_clk_dqb 8 vss vss hvtnfet l=6e-08 w=1.26e-06 $X=21495 $Y=22041 $D=616
M783 r_clk_dqb_n 9 vss vss hvtnfet l=6e-08 w=1.26e-06 $X=21495 $Y=29007 $D=616
M784 vss 10 r_lweb vss hvtnfet l=6e-08 w=1.287e-06 $X=21495 $Y=30897 $D=616
M785 r_sa_preb_n 51 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=21495 $Y=37027 $D=616
M786 rt_mb<3> 39 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=21495 $Y=38499 $D=616
M787 rt_mb<1> 40 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=21495 $Y=43487 $D=616
M788 rt_cb<3> 41 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=21495 $Y=44959 $D=616
M789 rt_cb<1> 42 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=21495 $Y=49947 $D=616
M790 vss 289 lb_ca<1> vss hvtnfet l=6e-08 w=8.58e-07 $X=22005 $Y=328 $D=616
M791 vss 290 lb_ca<3> vss hvtnfet l=6e-08 w=8.58e-07 $X=22005 $Y=5316 $D=616
M792 vss 291 lb_ma<1> vss hvtnfet l=6e-08 w=8.58e-07 $X=22005 $Y=6788 $D=616
M793 vss 292 lb_ma<3> vss hvtnfet l=6e-08 w=8.58e-07 $X=22005 $Y=11776 $D=616
M794 lb_tm_prea_n 285 vss vss hvtnfet l=6e-08 w=1.287e-06 $X=22005 $Y=13280 $D=616
M795 lt_tm_prea_n 286 vss vss hvtnfet l=6e-08 w=1.287e-06 $X=22005 $Y=20124 $D=616
M796 vss 287 l_clk_dqa vss hvtnfet l=6e-08 w=1.26e-06 $X=22005 $Y=22041 $D=616
M797 vss 288 l_clk_dqa_n vss hvtnfet l=6e-08 w=1.26e-06 $X=22005 $Y=29007 $D=616
M798 l_lwea 284 vss vss hvtnfet l=6e-08 w=1.287e-06 $X=22005 $Y=30897 $D=616
M799 vss 293 l_sa_prea_n vss hvtnfet l=6e-08 w=8.58e-07 $X=22005 $Y=37027 $D=616
M800 vss 294 lt_ma<3> vss hvtnfet l=6e-08 w=8.58e-07 $X=22005 $Y=38499 $D=616
M801 vss 295 lt_ma<1> vss hvtnfet l=6e-08 w=8.58e-07 $X=22005 $Y=43487 $D=616
M802 vss 296 lt_ca<3> vss hvtnfet l=6e-08 w=8.58e-07 $X=22005 $Y=44959 $D=616
M803 vss 297 lt_ca<1> vss hvtnfet l=6e-08 w=8.58e-07 $X=22005 $Y=49947 $D=616
M804 lb_ca<1> 289 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=22265 $Y=328 $D=616
M805 lb_ca<3> 290 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=22265 $Y=5316 $D=616
M806 lb_ma<1> 291 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=22265 $Y=6788 $D=616
M807 lb_ma<3> 292 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=22265 $Y=11776 $D=616
M808 vss 285 lb_tm_prea_n vss hvtnfet l=6e-08 w=1.287e-06 $X=22265 $Y=13280 $D=616
M809 vss 286 lt_tm_prea_n vss hvtnfet l=6e-08 w=1.287e-06 $X=22265 $Y=20124 $D=616
M810 l_clk_dqa 287 vss vss hvtnfet l=6e-08 w=1.26e-06 $X=22265 $Y=22041 $D=616
M811 l_clk_dqa_n 288 vss vss hvtnfet l=6e-08 w=1.26e-06 $X=22265 $Y=29007 $D=616
M812 vss 284 l_lwea vss hvtnfet l=6e-08 w=1.287e-06 $X=22265 $Y=30897 $D=616
M813 l_sa_prea_n 293 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=22265 $Y=37027 $D=616
M814 lt_ma<3> 294 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=22265 $Y=38499 $D=616
M815 lt_ma<1> 295 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=22265 $Y=43487 $D=616
M816 lt_ca<3> 296 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=22265 $Y=44959 $D=616
M817 lt_ca<1> 297 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=22265 $Y=49947 $D=616
M818 vss 289 lb_ca<1> vss hvtnfet l=6e-08 w=8.58e-07 $X=22525 $Y=328 $D=616
M819 vss 290 lb_ca<3> vss hvtnfet l=6e-08 w=8.58e-07 $X=22525 $Y=5316 $D=616
M820 vss 291 lb_ma<1> vss hvtnfet l=6e-08 w=8.58e-07 $X=22525 $Y=6788 $D=616
M821 vss 292 lb_ma<3> vss hvtnfet l=6e-08 w=8.58e-07 $X=22525 $Y=11776 $D=616
M822 vss 287 l_clk_dqa vss hvtnfet l=6e-08 w=1.26e-06 $X=22525 $Y=22041 $D=616
M823 vss 288 l_clk_dqa_n vss hvtnfet l=6e-08 w=1.26e-06 $X=22525 $Y=29007 $D=616
M824 vss 293 l_sa_prea_n vss hvtnfet l=6e-08 w=8.58e-07 $X=22525 $Y=37027 $D=616
M825 vss 294 lt_ma<3> vss hvtnfet l=6e-08 w=8.58e-07 $X=22525 $Y=38499 $D=616
M826 vss 295 lt_ma<1> vss hvtnfet l=6e-08 w=8.58e-07 $X=22525 $Y=43487 $D=616
M827 vss 296 lt_ca<3> vss hvtnfet l=6e-08 w=8.58e-07 $X=22525 $Y=44959 $D=616
M828 vss 297 lt_ca<1> vss hvtnfet l=6e-08 w=8.58e-07 $X=22525 $Y=49947 $D=616
M829 vss 298 284 vss hvtnfet l=6e-08 w=6e-07 $X=22775 $Y=30899 $D=616
M830 lb_ca<0> 299 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=22785 $Y=328 $D=616
M831 lb_ca<2> 300 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=22785 $Y=5316 $D=616
M832 lb_ma<0> 301 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=22785 $Y=6788 $D=616
M833 lb_ma<2> 302 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=22785 $Y=11776 $D=616
M834 l_saea_n 303 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=22785 $Y=37027 $D=616
M835 lt_ma<2> 304 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=22785 $Y=38499 $D=616
M836 lt_ma<0> 305 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=22785 $Y=43487 $D=616
M837 lt_ca<2> 306 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=22785 $Y=44959 $D=616
M838 lt_ca<0> 307 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=22785 $Y=49947 $D=616
M839 vss 299 lb_ca<0> vss hvtnfet l=6e-08 w=8.58e-07 $X=23045 $Y=328 $D=616
M840 vss 300 lb_ca<2> vss hvtnfet l=6e-08 w=8.58e-07 $X=23045 $Y=5316 $D=616
M841 vss 301 lb_ma<0> vss hvtnfet l=6e-08 w=8.58e-07 $X=23045 $Y=6788 $D=616
M842 vss 302 lb_ma<2> vss hvtnfet l=6e-08 w=8.58e-07 $X=23045 $Y=11776 $D=616
M843 vss 303 l_saea_n vss hvtnfet l=6e-08 w=8.58e-07 $X=23045 $Y=37027 $D=616
M844 vss 304 lt_ma<2> vss hvtnfet l=6e-08 w=8.58e-07 $X=23045 $Y=38499 $D=616
M845 vss 305 lt_ma<0> vss hvtnfet l=6e-08 w=8.58e-07 $X=23045 $Y=43487 $D=616
M846 vss 306 lt_ca<2> vss hvtnfet l=6e-08 w=8.58e-07 $X=23045 $Y=44959 $D=616
M847 vss 307 lt_ca<0> vss hvtnfet l=6e-08 w=8.58e-07 $X=23045 $Y=49947 $D=616
M848 1027 308 vss vss hvtnfet l=6e-08 w=1.8e-07 $X=23289 $Y=17143 $D=616
M849 308 312 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=23289 $Y=17812 $D=616
M850 309 313 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=23289 $Y=18983 $D=616
M851 1028 309 vss vss hvtnfet l=6e-08 w=1.8e-07 $X=23289 $Y=19609 $D=616
M852 1029 310 vss vss hvtnfet l=6e-08 w=1.8e-07 $X=23289 $Y=24063 $D=616
M853 310 314 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=23289 $Y=24732 $D=616
M854 311 315 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=23289 $Y=25903 $D=616
M855 1030 311 vss vss hvtnfet l=6e-08 w=1.8e-07 $X=23289 $Y=26529 $D=616
M856 lb_ca<0> 299 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=23305 $Y=328 $D=616
M857 lb_ca<2> 300 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=23305 $Y=5316 $D=616
M858 lb_ma<0> 301 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=23305 $Y=6788 $D=616
M859 lb_ma<2> 302 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=23305 $Y=11776 $D=616
M860 l_saea_n 303 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=23305 $Y=37027 $D=616
M861 lt_ma<2> 304 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=23305 $Y=38499 $D=616
M862 lt_ma<0> 305 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=23305 $Y=43487 $D=616
M863 lt_ca<2> 306 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=23305 $Y=44959 $D=616
M864 lt_ca<0> 307 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=23305 $Y=49947 $D=616
M865 312 317 1027 vss hvtnfet l=6e-08 w=1.8e-07 $X=23549 $Y=17143 $D=616
M866 vss 312 308 vss hvtnfet l=6e-08 w=1.37e-07 $X=23549 $Y=17812 $D=616
M867 vss 313 309 vss hvtnfet l=6e-08 w=1.37e-07 $X=23549 $Y=18983 $D=616
M868 313 317 1028 vss hvtnfet l=6e-08 w=1.8e-07 $X=23549 $Y=19609 $D=616
M869 314 317 1029 vss hvtnfet l=6e-08 w=1.8e-07 $X=23549 $Y=24063 $D=616
M870 vss 314 310 vss hvtnfet l=6e-08 w=1.37e-07 $X=23549 $Y=24732 $D=616
M871 vss 315 311 vss hvtnfet l=6e-08 w=1.37e-07 $X=23549 $Y=25903 $D=616
M872 315 317 1030 vss hvtnfet l=6e-08 w=1.8e-07 $X=23549 $Y=26529 $D=616
M873 vss 303 l_saea_n vss hvtnfet l=6e-08 w=8.58e-07 $X=23565 $Y=37027 $D=616
M874 l_saea_n 303 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=23825 $Y=37027 $D=616
M875 vss aa<0> 327 vss hvtnfet l=6e-08 w=2.74e-07 $X=23864 $Y=13476 $D=616
M876 vss 324 331 vss hvtnfet l=6e-08 w=2.1e-07 $X=24000 $Y=30918 $D=616
M877 vss 298 332 vss hvtnfet l=6e-08 w=2.1e-07 $X=24000 $Y=32688 $D=616
M878 1031 323 vss vss hvtnfet l=6e-08 w=8.23e-07 $X=24059 $Y=17143 $D=616
M879 1032 323 vss vss hvtnfet l=6e-08 w=8.23e-07 $X=24059 $Y=18966 $D=616
M880 1033 323 vss vss hvtnfet l=6e-08 w=8.23e-07 $X=24059 $Y=24063 $D=616
M881 1034 323 vss vss hvtnfet l=6e-08 w=8.23e-07 $X=24059 $Y=25886 $D=616
M882 b_pxca_n<7> 318 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=24060 $Y=336 $D=616
M883 318 319 vss vss hvtnfet l=6e-08 w=5e-07 $X=24060 $Y=6701 $D=616
M884 319 320 vss vss hvtnfet l=6e-08 w=3e-07 $X=24060 $Y=7831 $D=616
M885 321 320 vss vss hvtnfet l=6e-08 w=3e-07 $X=24060 $Y=43002 $D=616
M886 322 321 vss vss hvtnfet l=6e-08 w=5e-07 $X=24060 $Y=43932 $D=616
M887 t_pxca_n<7> 322 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=24060 $Y=49512 $D=616
M888 709 325 vss vss hvtnfet l=6e-08 w=4.8e-07 $X=24083 $Y=11276 $D=616
M889 710 clka vss vss hvtnfet l=6e-08 w=2.1e-07 $X=24260 $Y=30918 $D=616
M890 711 clka vss vss hvtnfet l=6e-08 w=2.1e-07 $X=24260 $Y=32688 $D=616
M891 vss 318 b_pxca_n<7> vss hvtnfet l=6e-08 w=1.285e-06 $X=24320 $Y=336 $D=616
M892 vss 319 318 vss hvtnfet l=6e-08 w=5e-07 $X=24320 $Y=6701 $D=616
M893 vss 320 319 vss hvtnfet l=6e-08 w=3e-07 $X=24320 $Y=7831 $D=616
M894 vss 320 321 vss hvtnfet l=6e-08 w=3e-07 $X=24320 $Y=43002 $D=616
M895 vss 321 322 vss hvtnfet l=6e-08 w=5e-07 $X=24320 $Y=43932 $D=616
M896 vss 322 t_pxca_n<7> vss hvtnfet l=6e-08 w=1.285e-06 $X=24320 $Y=49512 $D=616
M897 1035 328 1031 vss hvtnfet l=6e-08 w=5.49e-07 $X=24329 $Y=17143 $D=616
M898 1036 328 1032 vss hvtnfet l=6e-08 w=5.49e-07 $X=24329 $Y=19240 $D=616
M899 1037 329 1033 vss hvtnfet l=6e-08 w=5.49e-07 $X=24329 $Y=24063 $D=616
M900 1038 329 1034 vss hvtnfet l=6e-08 w=5.49e-07 $X=24329 $Y=26160 $D=616
M901 vss tm<8> 709 vss hvtnfet l=6e-08 w=4.8e-07 $X=24343 $Y=11276 $D=616
M902 334 327 vss vss hvtnfet l=6e-08 w=2.74e-07 $X=24374 $Y=13476 $D=616
M903 vss tm<5> 264 vss hvtnfet l=6e-08 w=2.74e-07 $X=24518 $Y=39358 $D=616
M904 324 331 710 vss hvtnfet l=6e-08 w=2.1e-07 $X=24520 $Y=30918 $D=616
M905 298 332 711 vss hvtnfet l=6e-08 w=2.1e-07 $X=24520 $Y=32688 $D=616
M906 312 334 1035 vss hvtnfet l=6e-08 w=5.49e-07 $X=24589 $Y=17143 $D=616
M907 313 327 1036 vss hvtnfet l=6e-08 w=5.49e-07 $X=24589 $Y=19240 $D=616
M908 314 334 1037 vss hvtnfet l=6e-08 w=5.49e-07 $X=24589 $Y=24063 $D=616
M909 315 327 1038 vss hvtnfet l=6e-08 w=5.49e-07 $X=24589 $Y=26160 $D=616
M910 714 340 324 vss hvtnfet l=6e-08 w=3.2e-07 $X=24780 $Y=30918 $D=616
M911 715 340 298 vss hvtnfet l=6e-08 w=3.2e-07 $X=24780 $Y=32578 $D=616
M912 b_pxca_n<6> 335 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=24830 $Y=336 $D=616
M913 335 336 vss vss hvtnfet l=6e-08 w=5e-07 $X=24830 $Y=6701 $D=616
M914 336 337 vss vss hvtnfet l=6e-08 w=3e-07 $X=24830 $Y=7831 $D=616
M915 338 337 vss vss hvtnfet l=6e-08 w=3e-07 $X=24830 $Y=43002 $D=616
M916 339 338 vss vss hvtnfet l=6e-08 w=5e-07 $X=24830 $Y=43932 $D=616
M917 t_pxca_n<6> 339 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=24830 $Y=49512 $D=616
M918 718 tm<8> vss vss hvtnfet l=6e-08 w=4.8e-07 $X=24853 $Y=11276 $D=616
M919 vss 264 376 vss hvtnfet l=6e-08 w=2e-07 $X=24874 $Y=37147 $D=616
M920 vss aa<1> 329 vss hvtnfet l=6e-08 w=2.74e-07 $X=24884 $Y=13476 $D=616
M921 vss aa<4> 714 vss hvtnfet l=6e-08 w=3.2e-07 $X=25040 $Y=30918 $D=616
M922 vss wena 715 vss hvtnfet l=6e-08 w=3.2e-07 $X=25040 $Y=32578 $D=616
M923 vss 335 b_pxca_n<6> vss hvtnfet l=6e-08 w=1.285e-06 $X=25090 $Y=336 $D=616
M924 vss 336 335 vss hvtnfet l=6e-08 w=5e-07 $X=25090 $Y=6701 $D=616
M925 vss 337 336 vss hvtnfet l=6e-08 w=3e-07 $X=25090 $Y=7831 $D=616
M926 vss 337 338 vss hvtnfet l=6e-08 w=3e-07 $X=25090 $Y=43002 $D=616
M927 vss 338 339 vss hvtnfet l=6e-08 w=5e-07 $X=25090 $Y=43932 $D=616
M928 vss 339 t_pxca_n<6> vss hvtnfet l=6e-08 w=1.285e-06 $X=25090 $Y=49512 $D=616
M929 vss tm<9> 718 vss hvtnfet l=6e-08 w=4.8e-07 $X=25113 $Y=11276 $D=616
M930 376 wena vss vss hvtnfet l=6e-08 w=2e-07 $X=25134 $Y=37147 $D=616
M931 328 329 vss vss hvtnfet l=6e-08 w=2.74e-07 $X=25394 $Y=13476 $D=616
M932 b_pxca_n<5> 345 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=25600 $Y=336 $D=616
M933 345 346 vss vss hvtnfet l=6e-08 w=5e-07 $X=25600 $Y=6701 $D=616
M934 346 347 vss vss hvtnfet l=6e-08 w=3e-07 $X=25600 $Y=7831 $D=616
M935 348 347 vss vss hvtnfet l=6e-08 w=3e-07 $X=25600 $Y=43002 $D=616
M936 349 348 vss vss hvtnfet l=6e-08 w=5e-07 $X=25600 $Y=43932 $D=616
M937 t_pxca_n<5> 349 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=25600 $Y=49512 $D=616
M938 1039 337 vss vss hvtnfet l=6e-08 w=1.8e-07 $X=25609 $Y=17143 $D=616
M939 1040 320 vss vss hvtnfet l=6e-08 w=1.8e-07 $X=25609 $Y=19609 $D=616
M940 1041 350 vss vss hvtnfet l=6e-08 w=1.8e-07 $X=25609 $Y=24063 $D=616
M941 1042 351 vss vss hvtnfet l=6e-08 w=1.8e-07 $X=25609 $Y=26529 $D=616
M942 721 tm<9> vss vss hvtnfet l=6e-08 w=4.8e-07 $X=25623 $Y=11276 $D=616
M943 337 352 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=25624 $Y=17812 $D=616
M944 320 353 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=25624 $Y=18983 $D=616
M945 350 354 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=25624 $Y=24732 $D=616
M946 351 355 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=25624 $Y=25903 $D=616
M947 vss clka 340 vss hvtnfet l=6e-08 w=4.5e-07 $X=25854 $Y=30668 $D=616
M948 vss 345 b_pxca_n<5> vss hvtnfet l=6e-08 w=1.285e-06 $X=25860 $Y=336 $D=616
M949 vss 346 345 vss hvtnfet l=6e-08 w=5e-07 $X=25860 $Y=6701 $D=616
M950 vss 347 346 vss hvtnfet l=6e-08 w=3e-07 $X=25860 $Y=7831 $D=616
M951 vss 347 348 vss hvtnfet l=6e-08 w=3e-07 $X=25860 $Y=43002 $D=616
M952 vss 348 349 vss hvtnfet l=6e-08 w=5e-07 $X=25860 $Y=43932 $D=616
M953 vss 349 t_pxca_n<5> vss hvtnfet l=6e-08 w=1.285e-06 $X=25860 $Y=49512 $D=616
M954 352 317 1039 vss hvtnfet l=6e-08 w=1.8e-07 $X=25869 $Y=17143 $D=616
M955 353 317 1040 vss hvtnfet l=6e-08 w=1.8e-07 $X=25869 $Y=19609 $D=616
M956 354 317 1041 vss hvtnfet l=6e-08 w=1.8e-07 $X=25869 $Y=24063 $D=616
M957 355 317 1042 vss hvtnfet l=6e-08 w=1.8e-07 $X=25869 $Y=26529 $D=616
M958 vss 366 721 vss hvtnfet l=6e-08 w=4.8e-07 $X=25883 $Y=11276 $D=616
M959 vss 352 337 vss hvtnfet l=6e-08 w=1.37e-07 $X=25884 $Y=17812 $D=616
M960 vss 353 320 vss hvtnfet l=6e-08 w=1.37e-07 $X=25884 $Y=18983 $D=616
M961 vss 354 350 vss hvtnfet l=6e-08 w=1.37e-07 $X=25884 $Y=24732 $D=616
M962 vss 355 351 vss hvtnfet l=6e-08 w=1.37e-07 $X=25884 $Y=25903 $D=616
M963 vss 356 363 vss hvtnfet l=6e-08 w=2.1e-07 $X=26138 $Y=37277 $D=616
M964 b_pxca_n<4> 357 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=26370 $Y=336 $D=616
M965 357 358 vss vss hvtnfet l=6e-08 w=5e-07 $X=26370 $Y=6701 $D=616
M966 358 359 vss vss hvtnfet l=6e-08 w=3e-07 $X=26370 $Y=7831 $D=616
M967 360 359 vss vss hvtnfet l=6e-08 w=3e-07 $X=26370 $Y=43002 $D=616
M968 361 360 vss vss hvtnfet l=6e-08 w=5e-07 $X=26370 $Y=43932 $D=616
M969 t_pxca_n<4> 361 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=26370 $Y=49512 $D=616
M970 729 123 733 vss hvtnfet l=6e-08 w=6e-07 $X=26374 $Y=30668 $D=616
M971 1043 323 vss vss hvtnfet l=6e-08 w=8.23e-07 $X=26379 $Y=17143 $D=616
M972 1044 323 vss vss hvtnfet l=6e-08 w=8.23e-07 $X=26379 $Y=18966 $D=616
M973 1045 323 vss vss hvtnfet l=6e-08 w=8.23e-07 $X=26379 $Y=24063 $D=616
M974 1046 323 vss vss hvtnfet l=6e-08 w=8.23e-07 $X=26379 $Y=25886 $D=616
M975 vss 366 727 vss hvtnfet l=6e-08 w=4.8e-07 $X=26393 $Y=11276 $D=616
M976 724 362 vss vss hvtnfet l=6e-08 w=2.1e-07 $X=26398 $Y=37277 $D=616
M977 vss 357 b_pxca_n<4> vss hvtnfet l=6e-08 w=1.285e-06 $X=26630 $Y=336 $D=616
M978 vss 358 357 vss hvtnfet l=6e-08 w=5e-07 $X=26630 $Y=6701 $D=616
M979 vss 359 358 vss hvtnfet l=6e-08 w=3e-07 $X=26630 $Y=7831 $D=616
M980 vss 359 360 vss hvtnfet l=6e-08 w=3e-07 $X=26630 $Y=43002 $D=616
M981 vss 360 361 vss hvtnfet l=6e-08 w=5e-07 $X=26630 $Y=43932 $D=616
M982 vss 361 t_pxca_n<4> vss hvtnfet l=6e-08 w=1.285e-06 $X=26630 $Y=49512 $D=616
M983 733 123 729 vss hvtnfet l=6e-08 w=6e-07 $X=26634 $Y=30668 $D=616
M984 1047 364 1043 vss hvtnfet l=6e-08 w=5.49e-07 $X=26649 $Y=17417 $D=616
M985 1048 364 1044 vss hvtnfet l=6e-08 w=5.49e-07 $X=26649 $Y=18966 $D=616
M986 1049 365 1045 vss hvtnfet l=6e-08 w=5.49e-07 $X=26649 $Y=24337 $D=616
M987 1050 365 1046 vss hvtnfet l=6e-08 w=5.49e-07 $X=26649 $Y=25886 $D=616
M988 727 325 vss vss hvtnfet l=6e-08 w=4.8e-07 $X=26653 $Y=11276 $D=616
M989 356 363 724 vss hvtnfet l=6e-08 w=2.1e-07 $X=26658 $Y=37277 $D=616
M990 vss tm<7> 726 vss hvtnfet l=6e-08 w=2.74e-07 $X=26820 $Y=39358 $D=616
M991 728 123 vss vss hvtnfet l=6e-08 w=3.2e-07 $X=26839 $Y=32578 $D=616
M992 vss 123 733 vss hvtnfet l=6e-08 w=6e-07 $X=26894 $Y=30668 $D=616
M993 1051 369 1047 vss hvtnfet l=6e-08 w=5.49e-07 $X=26909 $Y=17417 $D=616
M994 1052 369 1048 vss hvtnfet l=6e-08 w=5.49e-07 $X=26909 $Y=18966 $D=616
M995 1053 369 1049 vss hvtnfet l=6e-08 w=5.49e-07 $X=26909 $Y=24337 $D=616
M996 1054 369 1050 vss hvtnfet l=6e-08 w=5.49e-07 $X=26909 $Y=25886 $D=616
M997 730 368 356 vss hvtnfet l=6e-08 w=3.2e-07 $X=26918 $Y=37277 $D=616
M998 vss aa<10> 374 vss hvtnfet l=6e-08 w=2.74e-07 $X=26924 $Y=13476 $D=616
M999 379 123 728 vss hvtnfet l=6e-08 w=3.2e-07 $X=27099 $Y=32578 $D=616
M1000 b_pxca_n<3> 370 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=27140 $Y=336 $D=616
M1001 370 371 vss vss hvtnfet l=6e-08 w=5e-07 $X=27140 $Y=6701 $D=616
M1002 371 351 vss vss hvtnfet l=6e-08 w=3e-07 $X=27140 $Y=7831 $D=616
M1003 372 351 vss vss hvtnfet l=6e-08 w=3e-07 $X=27140 $Y=43002 $D=616
M1004 373 372 vss vss hvtnfet l=6e-08 w=5e-07 $X=27140 $Y=43932 $D=616
M1005 t_pxca_n<3> 373 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=27140 $Y=49512 $D=616
M1006 733 123 vss vss hvtnfet l=6e-08 w=6e-07 $X=27154 $Y=30668 $D=616
M1007 vss tm<9> 325 vss hvtnfet l=7e-08 w=3.2e-07 $X=27163 $Y=11276 $D=616
M1008 352 374 1051 vss hvtnfet l=6e-08 w=5.49e-07 $X=27169 $Y=17417 $D=616
M1009 353 375 1052 vss hvtnfet l=6e-08 w=5.49e-07 $X=27169 $Y=18966 $D=616
M1010 354 374 1053 vss hvtnfet l=6e-08 w=5.49e-07 $X=27169 $Y=24337 $D=616
M1011 355 375 1054 vss hvtnfet l=6e-08 w=5.49e-07 $X=27169 $Y=25886 $D=616
M1012 vss 376 730 vss hvtnfet l=6e-08 w=3.2e-07 $X=27178 $Y=37277 $D=616
M1013 375 374 vss vss hvtnfet l=6e-08 w=2.74e-07 $X=27184 $Y=13476 $D=616
M1014 734 377 379 vss hvtnfet l=6e-08 w=2.1e-07 $X=27359 $Y=32688 $D=616
M1015 vss 370 b_pxca_n<3> vss hvtnfet l=6e-08 w=1.285e-06 $X=27400 $Y=336 $D=616
M1016 vss 371 370 vss hvtnfet l=6e-08 w=5e-07 $X=27400 $Y=6701 $D=616
M1017 vss 351 371 vss hvtnfet l=6e-08 w=3e-07 $X=27400 $Y=7831 $D=616
M1018 vss 351 372 vss hvtnfet l=6e-08 w=3e-07 $X=27400 $Y=43002 $D=616
M1019 vss 372 373 vss hvtnfet l=6e-08 w=5e-07 $X=27400 $Y=43932 $D=616
M1020 vss 373 t_pxca_n<3> vss hvtnfet l=6e-08 w=1.285e-06 $X=27400 $Y=49512 $D=616
M1021 366 tm<8> vss vss hvtnfet l=7e-08 w=3.2e-07 $X=27433 $Y=11276 $D=616
M1022 vss 131 734 vss hvtnfet l=6e-08 w=2.1e-07 $X=27619 $Y=32688 $D=616
M1023 vss tm<1> 735 vss hvtnfet l=6e-08 w=2.74e-07 $X=27620 $Y=39358 $D=616
M1024 vss 380 369 vss hvtnfet l=6e-08 w=2.74e-07 $X=27784 $Y=13476 $D=616
M1025 737 362 386 vss hvtnfet l=6e-08 w=4e-07 $X=27858 $Y=37045 $D=616
M1026 377 379 vss vss hvtnfet l=6e-08 w=2.1e-07 $X=27879 $Y=32688 $D=616
M1027 b_pxca_n<2> 381 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=27910 $Y=336 $D=616
M1028 381 382 vss vss hvtnfet l=6e-08 w=5e-07 $X=27910 $Y=6701 $D=616
M1029 382 350 vss vss hvtnfet l=6e-08 w=3e-07 $X=27910 $Y=7831 $D=616
M1030 383 350 vss vss hvtnfet l=6e-08 w=3e-07 $X=27910 $Y=43002 $D=616
M1031 384 383 vss vss hvtnfet l=6e-08 w=5e-07 $X=27910 $Y=43932 $D=616
M1032 t_pxca_n<2> 384 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=27910 $Y=49512 $D=616
M1033 vss 323 317 vss hvtnfet l=6e-08 w=7e-07 $X=27924 $Y=30668 $D=616
M1034 380 aa<11> vss vss hvtnfet l=6e-08 w=2.74e-07 $X=28044 $Y=13476 $D=616
M1035 vss 356 737 vss hvtnfet l=6e-08 w=4e-07 $X=28118 $Y=37045 $D=616
M1036 vss 381 b_pxca_n<2> vss hvtnfet l=6e-08 w=1.285e-06 $X=28170 $Y=336 $D=616
M1037 vss 382 381 vss hvtnfet l=6e-08 w=5e-07 $X=28170 $Y=6701 $D=616
M1038 vss 350 382 vss hvtnfet l=6e-08 w=3e-07 $X=28170 $Y=7831 $D=616
M1039 vss 350 383 vss hvtnfet l=6e-08 w=3e-07 $X=28170 $Y=43002 $D=616
M1040 vss 383 384 vss hvtnfet l=6e-08 w=5e-07 $X=28170 $Y=43932 $D=616
M1041 vss 384 t_pxca_n<2> vss hvtnfet l=6e-08 w=1.285e-06 $X=28170 $Y=49512 $D=616
M1042 317 323 vss vss hvtnfet l=6e-08 w=7e-07 $X=28184 $Y=30668 $D=616
M1043 vss 392 541 vss hvtnfet l=6e-08 w=2e-07 $X=28514 $Y=11276 $D=616
M1044 vss 393 544 vss hvtnfet l=6e-08 w=2e-07 $X=28514 $Y=39657 $D=616
M1045 494 386 vss vss hvtnfet l=6e-08 w=2e-07 $X=28628 $Y=37045 $D=616
M1046 b_pxca_n<1> 387 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=28680 $Y=336 $D=616
M1047 387 388 vss vss hvtnfet l=6e-08 w=5e-07 $X=28680 $Y=6701 $D=616
M1048 388 389 vss vss hvtnfet l=6e-08 w=3e-07 $X=28680 $Y=7831 $D=616
M1049 390 389 vss vss hvtnfet l=6e-08 w=3e-07 $X=28680 $Y=43002 $D=616
M1050 391 390 vss vss hvtnfet l=6e-08 w=5e-07 $X=28680 $Y=43932 $D=616
M1051 t_pxca_n<1> 391 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=28680 $Y=49512 $D=616
M1052 742 123 vss vss hvtnfet l=6e-08 w=6e-07 $X=28704 $Y=30668 $D=616
M1053 vss 387 b_pxca_n<1> vss hvtnfet l=6e-08 w=1.285e-06 $X=28940 $Y=336 $D=616
M1054 vss 388 387 vss hvtnfet l=6e-08 w=5e-07 $X=28940 $Y=6701 $D=616
M1055 vss 389 388 vss hvtnfet l=6e-08 w=3e-07 $X=28940 $Y=7831 $D=616
M1056 vss 389 390 vss hvtnfet l=6e-08 w=3e-07 $X=28940 $Y=43002 $D=616
M1057 vss 390 391 vss hvtnfet l=6e-08 w=5e-07 $X=28940 $Y=43932 $D=616
M1058 vss 391 t_pxca_n<1> vss hvtnfet l=6e-08 w=1.285e-06 $X=28940 $Y=49512 $D=616
M1059 1055 374 407 vss hvtnfet l=6e-08 w=5.49e-07 $X=29009 $Y=17417 $D=616
M1060 1056 375 408 vss hvtnfet l=6e-08 w=5.49e-07 $X=29009 $Y=18966 $D=616
M1061 1057 374 409 vss hvtnfet l=6e-08 w=5.49e-07 $X=29009 $Y=24337 $D=616
M1062 1058 375 410 vss hvtnfet l=6e-08 w=5.49e-07 $X=29009 $Y=25886 $D=616
M1063 1059 308 vss vss hvtnfet l=6e-08 w=4.11e-07 $X=29024 $Y=11276 $D=616
M1064 1060 308 vss vss hvtnfet l=6e-08 w=4.11e-07 $X=29024 $Y=39446 $D=616
M1065 vss aa<12> 365 vss hvtnfet l=6e-08 w=2.74e-07 $X=29054 $Y=13476 $D=616
M1066 1061 380 1055 vss hvtnfet l=6e-08 w=5.49e-07 $X=29269 $Y=17417 $D=616
M1067 1062 380 1056 vss hvtnfet l=6e-08 w=5.49e-07 $X=29269 $Y=18966 $D=616
M1068 1063 380 1057 vss hvtnfet l=6e-08 w=5.49e-07 $X=29269 $Y=24337 $D=616
M1069 1064 380 1058 vss hvtnfet l=6e-08 w=5.49e-07 $X=29269 $Y=25886 $D=616
M1070 392 dwla<1> 1059 vss hvtnfet l=6e-08 w=4.11e-07 $X=29284 $Y=11276 $D=616
M1071 393 dwla<0> 1060 vss hvtnfet l=6e-08 w=4.11e-07 $X=29284 $Y=39446 $D=616
M1072 vss 395 403 vss hvtnfet l=6e-08 w=2e-07 $X=29298 $Y=32533 $D=616
M1073 b_pxca_n<0> 396 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=29450 $Y=336 $D=616
M1074 396 397 vss vss hvtnfet l=6e-08 w=5e-07 $X=29450 $Y=6701 $D=616
M1075 397 398 vss vss hvtnfet l=6e-08 w=3e-07 $X=29450 $Y=7831 $D=616
M1076 399 398 vss vss hvtnfet l=6e-08 w=3e-07 $X=29450 $Y=43002 $D=616
M1077 400 399 vss vss hvtnfet l=6e-08 w=5e-07 $X=29450 $Y=43932 $D=616
M1078 t_pxca_n<0> 400 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=29450 $Y=49512 $D=616
M1079 1065 364 1061 vss hvtnfet l=6e-08 w=5.49e-07 $X=29529 $Y=17417 $D=616
M1080 1066 364 1062 vss hvtnfet l=6e-08 w=5.49e-07 $X=29529 $Y=18966 $D=616
M1081 1067 365 1063 vss hvtnfet l=6e-08 w=5.49e-07 $X=29529 $Y=24337 $D=616
M1082 1068 365 1064 vss hvtnfet l=6e-08 w=5.49e-07 $X=29529 $Y=25886 $D=616
M1083 403 405 vss vss hvtnfet l=6e-08 w=2e-07 $X=29558 $Y=32533 $D=616
M1084 364 365 vss vss hvtnfet l=6e-08 w=2.74e-07 $X=29564 $Y=13476 $D=616
M1085 vss 404 395 vss hvtnfet l=6e-08 w=3.5e-07 $X=29621 $Y=30853 $D=616
M1086 vss 396 b_pxca_n<0> vss hvtnfet l=6e-08 w=1.285e-06 $X=29710 $Y=336 $D=616
M1087 vss 397 396 vss hvtnfet l=6e-08 w=5e-07 $X=29710 $Y=6701 $D=616
M1088 vss 398 397 vss hvtnfet l=6e-08 w=3e-07 $X=29710 $Y=7831 $D=616
M1089 vss 398 399 vss hvtnfet l=6e-08 w=3e-07 $X=29710 $Y=43002 $D=616
M1090 vss 399 400 vss hvtnfet l=6e-08 w=5e-07 $X=29710 $Y=43932 $D=616
M1091 vss 400 t_pxca_n<0> vss hvtnfet l=6e-08 w=1.285e-06 $X=29710 $Y=49512 $D=616
M1092 456 403 vss vss hvtnfet l=6e-08 w=6e-07 $X=29747 $Y=37037 $D=616
M1093 vss 323 1065 vss hvtnfet l=6e-08 w=8.23e-07 $X=29799 $Y=17143 $D=616
M1094 vss 323 1066 vss hvtnfet l=6e-08 w=8.23e-07 $X=29799 $Y=18966 $D=616
M1095 vss 323 1067 vss hvtnfet l=6e-08 w=8.23e-07 $X=29799 $Y=24063 $D=616
M1096 vss 323 1068 vss hvtnfet l=6e-08 w=8.23e-07 $X=29799 $Y=25886 $D=616
M1097 404 406 vss vss hvtnfet l=2.5e-07 w=3.5e-07 $X=29881 $Y=30853 $D=616
M1098 405 tm<7> vss vss hvtnfet l=6e-08 w=2e-07 $X=30068 $Y=32533 $D=616
M1099 dbl_pd_n<3> 131 vss vss hvtnfet l=6e-08 w=2.14e-07 $X=30204 $Y=13361 $D=616
M1100 b_pxba_n<7> 411 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=30220 $Y=336 $D=616
M1101 411 412 vss vss hvtnfet l=6e-08 w=5e-07 $X=30220 $Y=6701 $D=616
M1102 412 413 vss vss hvtnfet l=6e-08 w=3e-07 $X=30220 $Y=7831 $D=616
M1103 414 413 vss vss hvtnfet l=6e-08 w=3e-07 $X=30220 $Y=43002 $D=616
M1104 415 414 vss vss hvtnfet l=6e-08 w=5e-07 $X=30220 $Y=43932 $D=616
M1105 t_pxba_n<7> 415 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=30220 $Y=49512 $D=616
M1106 359 407 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=30294 $Y=17812 $D=616
M1107 347 408 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=30294 $Y=18983 $D=616
M1108 398 409 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=30294 $Y=24732 $D=616
M1109 389 410 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=30294 $Y=25903 $D=616
M1110 1069 317 407 vss hvtnfet l=6e-08 w=1.8e-07 $X=30309 $Y=17143 $D=616
M1111 1070 317 408 vss hvtnfet l=6e-08 w=1.8e-07 $X=30309 $Y=19609 $D=616
M1112 1071 317 409 vss hvtnfet l=6e-08 w=1.8e-07 $X=30309 $Y=24063 $D=616
M1113 1072 317 410 vss hvtnfet l=6e-08 w=1.8e-07 $X=30309 $Y=26529 $D=616
M1114 vss 131 dbl_pd_n<3> vss hvtnfet l=6e-08 w=2.14e-07 $X=30464 $Y=13361 $D=616
M1115 vss 411 b_pxba_n<7> vss hvtnfet l=6e-08 w=1.285e-06 $X=30480 $Y=336 $D=616
M1116 vss 412 411 vss hvtnfet l=6e-08 w=5e-07 $X=30480 $Y=6701 $D=616
M1117 vss 413 412 vss hvtnfet l=6e-08 w=3e-07 $X=30480 $Y=7831 $D=616
M1118 vss 413 414 vss hvtnfet l=6e-08 w=3e-07 $X=30480 $Y=43002 $D=616
M1119 vss 414 415 vss hvtnfet l=6e-08 w=5e-07 $X=30480 $Y=43932 $D=616
M1120 vss 415 t_pxba_n<7> vss hvtnfet l=6e-08 w=1.285e-06 $X=30480 $Y=49512 $D=616
M1121 456 416 vss vss hvtnfet l=6e-08 w=6e-07 $X=30527 $Y=37037 $D=616
M1122 vss 407 359 vss hvtnfet l=6e-08 w=1.37e-07 $X=30554 $Y=17812 $D=616
M1123 vss 408 347 vss hvtnfet l=6e-08 w=1.37e-07 $X=30554 $Y=18983 $D=616
M1124 vss 409 398 vss hvtnfet l=6e-08 w=1.37e-07 $X=30554 $Y=24732 $D=616
M1125 vss 410 389 vss hvtnfet l=6e-08 w=1.37e-07 $X=30554 $Y=25903 $D=616
M1126 vss 359 1069 vss hvtnfet l=6e-08 w=1.8e-07 $X=30569 $Y=17143 $D=616
M1127 vss 347 1070 vss hvtnfet l=6e-08 w=1.8e-07 $X=30569 $Y=19609 $D=616
M1128 vss 398 1071 vss hvtnfet l=6e-08 w=1.8e-07 $X=30569 $Y=24063 $D=616
M1129 vss 389 1072 vss hvtnfet l=6e-08 w=1.8e-07 $X=30569 $Y=26529 $D=616
M1130 1073 dwla<1> 426 vss hvtnfet l=6e-08 w=4.11e-07 $X=30584 $Y=11276 $D=616
M1131 1074 dwla<0> 427 vss hvtnfet l=6e-08 w=4.11e-07 $X=30584 $Y=39446 $D=616
M1132 vss 406 416 vss hvtnfet l=6e-08 w=2e-07 $X=30644 $Y=32533 $D=616
M1133 dbl_pd_n<3> 131 vss vss hvtnfet l=6e-08 w=2.14e-07 $X=30724 $Y=13361 $D=616
M1134 vss 417 406 vss hvtnfet l=6e-08 w=3.5e-07 $X=30741 $Y=30853 $D=616
M1135 vss 309 1073 vss hvtnfet l=6e-08 w=4.11e-07 $X=30844 $Y=11276 $D=616
M1136 vss 309 1074 vss hvtnfet l=6e-08 w=4.11e-07 $X=30844 $Y=39446 $D=616
M1137 416 423 vss vss hvtnfet l=6e-08 w=2e-07 $X=30904 $Y=32533 $D=616
M1138 b_pxba_n<6> 418 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=30990 $Y=336 $D=616
M1139 418 419 vss vss hvtnfet l=6e-08 w=5e-07 $X=30990 $Y=6701 $D=616
M1140 419 420 vss vss hvtnfet l=6e-08 w=3e-07 $X=30990 $Y=7831 $D=616
M1141 421 420 vss vss hvtnfet l=6e-08 w=3e-07 $X=30990 $Y=43002 $D=616
M1142 422 421 vss vss hvtnfet l=6e-08 w=5e-07 $X=30990 $Y=43932 $D=616
M1143 t_pxba_n<6> 422 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=30990 $Y=49512 $D=616
M1144 417 368 vss vss hvtnfet l=2.5e-07 w=3.5e-07 $X=31001 $Y=30853 $D=616
M1145 1075 420 vss vss hvtnfet l=6e-08 w=1.8e-07 $X=31079 $Y=17143 $D=616
M1146 1076 413 vss vss hvtnfet l=6e-08 w=1.8e-07 $X=31079 $Y=19609 $D=616
M1147 1077 424 vss vss hvtnfet l=6e-08 w=1.8e-07 $X=31079 $Y=24063 $D=616
M1148 1078 425 vss vss hvtnfet l=6e-08 w=1.8e-07 $X=31079 $Y=26529 $D=616
M1149 420 428 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=31094 $Y=17812 $D=616
M1150 413 429 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=31094 $Y=18983 $D=616
M1151 424 430 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=31094 $Y=24732 $D=616
M1152 425 431 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=31094 $Y=25903 $D=616
M1153 dbl_pd_n<1> tm<1> vss vss hvtnfet l=6e-08 w=2.14e-07 $X=31234 $Y=13361 $D=616
M1154 vss 418 b_pxba_n<6> vss hvtnfet l=6e-08 w=1.285e-06 $X=31250 $Y=336 $D=616
M1155 vss 419 418 vss hvtnfet l=6e-08 w=5e-07 $X=31250 $Y=6701 $D=616
M1156 vss 420 419 vss hvtnfet l=6e-08 w=3e-07 $X=31250 $Y=7831 $D=616
M1157 vss 420 421 vss hvtnfet l=6e-08 w=3e-07 $X=31250 $Y=43002 $D=616
M1158 vss 421 422 vss hvtnfet l=6e-08 w=5e-07 $X=31250 $Y=43932 $D=616
M1159 vss 422 t_pxba_n<6> vss hvtnfet l=6e-08 w=1.285e-06 $X=31250 $Y=49512 $D=616
M1160 456 362 vss vss hvtnfet l=6e-08 w=6e-07 $X=31307 $Y=37037 $D=616
M1161 428 317 1075 vss hvtnfet l=6e-08 w=1.8e-07 $X=31339 $Y=17143 $D=616
M1162 429 317 1076 vss hvtnfet l=6e-08 w=1.8e-07 $X=31339 $Y=19609 $D=616
M1163 430 317 1077 vss hvtnfet l=6e-08 w=1.8e-07 $X=31339 $Y=24063 $D=616
M1164 431 317 1078 vss hvtnfet l=6e-08 w=1.8e-07 $X=31339 $Y=26529 $D=616
M1165 556 426 vss vss hvtnfet l=6e-08 w=2e-07 $X=31354 $Y=11276 $D=616
M1166 vss 428 420 vss hvtnfet l=6e-08 w=1.37e-07 $X=31354 $Y=17812 $D=616
M1167 vss 429 413 vss hvtnfet l=6e-08 w=1.37e-07 $X=31354 $Y=18983 $D=616
M1168 vss 430 424 vss hvtnfet l=6e-08 w=1.37e-07 $X=31354 $Y=24732 $D=616
M1169 vss 431 425 vss hvtnfet l=6e-08 w=1.37e-07 $X=31354 $Y=25903 $D=616
M1170 558 427 vss vss hvtnfet l=6e-08 w=2e-07 $X=31354 $Y=39657 $D=616
M1171 vss 173 423 vss hvtnfet l=6e-08 w=2e-07 $X=31414 $Y=32533 $D=616
M1172 vss tm<1> dbl_pd_n<1> vss hvtnfet l=6e-08 w=2.14e-07 $X=31494 $Y=13361 $D=616
M1173 dbl_pd_n<1> tm<1> vss vss hvtnfet l=6e-08 w=2.14e-07 $X=31754 $Y=13361 $D=616
M1174 b_pxba_n<5> 432 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=31760 $Y=336 $D=616
M1175 432 433 vss vss hvtnfet l=6e-08 w=5e-07 $X=31760 $Y=6701 $D=616
M1176 433 434 vss vss hvtnfet l=6e-08 w=3e-07 $X=31760 $Y=7831 $D=616
M1177 435 434 vss vss hvtnfet l=6e-08 w=3e-07 $X=31760 $Y=43002 $D=616
M1178 436 435 vss vss hvtnfet l=6e-08 w=5e-07 $X=31760 $Y=43932 $D=616
M1179 t_pxba_n<5> 436 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=31760 $Y=49512 $D=616
M1180 vss 368 362 vss hvtnfet l=6e-08 w=2e-07 $X=31761 $Y=31098 $D=616
M1181 1079 323 vss vss hvtnfet l=6e-08 w=8.23e-07 $X=31849 $Y=17143 $D=616
M1182 1080 323 vss vss hvtnfet l=6e-08 w=8.23e-07 $X=31849 $Y=18966 $D=616
M1183 1081 323 vss vss hvtnfet l=6e-08 w=8.23e-07 $X=31849 $Y=24063 $D=616
M1184 1082 323 vss vss hvtnfet l=6e-08 w=8.23e-07 $X=31849 $Y=25886 $D=616
M1185 vss 437 540 vss hvtnfet l=6e-08 w=2e-07 $X=31864 $Y=11276 $D=616
M1186 vss 438 545 vss hvtnfet l=6e-08 w=2e-07 $X=31864 $Y=39657 $D=616
M1187 vss 432 b_pxba_n<5> vss hvtnfet l=6e-08 w=1.285e-06 $X=32020 $Y=336 $D=616
M1188 vss 433 432 vss hvtnfet l=6e-08 w=5e-07 $X=32020 $Y=6701 $D=616
M1189 vss 434 433 vss hvtnfet l=6e-08 w=3e-07 $X=32020 $Y=7831 $D=616
M1190 vss 434 435 vss hvtnfet l=6e-08 w=3e-07 $X=32020 $Y=43002 $D=616
M1191 vss 435 436 vss hvtnfet l=6e-08 w=5e-07 $X=32020 $Y=43932 $D=616
M1192 vss 436 t_pxba_n<5> vss hvtnfet l=6e-08 w=1.285e-06 $X=32020 $Y=49512 $D=616
M1193 1083 439 1079 vss hvtnfet l=6e-08 w=5.49e-07 $X=32119 $Y=17417 $D=616
M1194 1084 439 1080 vss hvtnfet l=6e-08 w=5.49e-07 $X=32119 $Y=18966 $D=616
M1195 1085 440 1081 vss hvtnfet l=6e-08 w=5.49e-07 $X=32119 $Y=24337 $D=616
M1196 1086 440 1082 vss hvtnfet l=6e-08 w=5.49e-07 $X=32119 $Y=25886 $D=616
M1197 dwla<1> 442 vss vss hvtnfet l=6e-08 w=3e-07 $X=32271 $Y=31098 $D=616
M1198 497 442 vss vss hvtnfet l=6e-08 w=3e-07 $X=32271 $Y=37457 $D=616
M1199 1087 310 vss vss hvtnfet l=6e-08 w=4.11e-07 $X=32374 $Y=11276 $D=616
M1200 1088 310 vss vss hvtnfet l=6e-08 w=4.11e-07 $X=32374 $Y=39446 $D=616
M1201 1089 443 1083 vss hvtnfet l=6e-08 w=5.49e-07 $X=32379 $Y=17417 $D=616
M1202 1090 443 1084 vss hvtnfet l=6e-08 w=5.49e-07 $X=32379 $Y=18966 $D=616
M1203 1091 443 1085 vss hvtnfet l=6e-08 w=5.49e-07 $X=32379 $Y=24337 $D=616
M1204 1092 443 1086 vss hvtnfet l=6e-08 w=5.49e-07 $X=32379 $Y=25886 $D=616
M1205 vss aa<7> 449 vss hvtnfet l=6e-08 w=2.74e-07 $X=32394 $Y=13476 $D=616
M1206 vss 324 442 vss hvtnfet l=6e-08 w=5e-07 $X=32394 $Y=32443 $D=616
M1207 b_pxba_n<4> 444 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=32530 $Y=336 $D=616
M1208 444 445 vss vss hvtnfet l=6e-08 w=5e-07 $X=32530 $Y=6701 $D=616
M1209 445 446 vss vss hvtnfet l=6e-08 w=3e-07 $X=32530 $Y=7831 $D=616
M1210 447 446 vss vss hvtnfet l=6e-08 w=3e-07 $X=32530 $Y=43002 $D=616
M1211 448 447 vss vss hvtnfet l=6e-08 w=5e-07 $X=32530 $Y=43932 $D=616
M1212 t_pxba_n<4> 448 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=32530 $Y=49512 $D=616
M1213 vss 442 dwla<1> vss hvtnfet l=6e-08 w=3e-07 $X=32531 $Y=31098 $D=616
M1214 vss 442 497 vss hvtnfet l=6e-08 w=3e-07 $X=32531 $Y=37457 $D=616
M1215 437 dwla<1> 1087 vss hvtnfet l=6e-08 w=4.11e-07 $X=32634 $Y=11276 $D=616
M1216 438 dwla<0> 1088 vss hvtnfet l=6e-08 w=4.11e-07 $X=32634 $Y=39446 $D=616
M1217 428 449 1089 vss hvtnfet l=6e-08 w=5.49e-07 $X=32639 $Y=17417 $D=616
M1218 429 450 1090 vss hvtnfet l=6e-08 w=5.49e-07 $X=32639 $Y=18966 $D=616
M1219 430 449 1091 vss hvtnfet l=6e-08 w=5.49e-07 $X=32639 $Y=24337 $D=616
M1220 431 450 1092 vss hvtnfet l=6e-08 w=5.49e-07 $X=32639 $Y=25886 $D=616
M1221 450 449 vss vss hvtnfet l=6e-08 w=2.74e-07 $X=32654 $Y=13476 $D=616
M1222 vss 444 b_pxba_n<4> vss hvtnfet l=6e-08 w=1.285e-06 $X=32790 $Y=336 $D=616
M1223 vss 445 444 vss hvtnfet l=6e-08 w=5e-07 $X=32790 $Y=6701 $D=616
M1224 vss 446 445 vss hvtnfet l=6e-08 w=3e-07 $X=32790 $Y=7831 $D=616
M1225 vss 446 447 vss hvtnfet l=6e-08 w=3e-07 $X=32790 $Y=43002 $D=616
M1226 vss 447 448 vss hvtnfet l=6e-08 w=5e-07 $X=32790 $Y=43932 $D=616
M1227 vss 448 t_pxba_n<4> vss hvtnfet l=6e-08 w=1.285e-06 $X=32790 $Y=49512 $D=616
M1228 dwla<1> 368 vss vss hvtnfet l=6e-08 w=3e-07 $X=33041 $Y=31098 $D=616
M1229 497 456 vss vss hvtnfet l=6e-08 w=3e-07 $X=33041 $Y=37457 $D=616
M1230 465 442 vss vss hvtnfet l=6e-08 w=4e-07 $X=33094 $Y=32543 $D=616
M1231 1093 dwla<1> 458 vss hvtnfet l=6e-08 w=4.11e-07 $X=33144 $Y=11276 $D=616
M1232 1094 dwla<0> 459 vss hvtnfet l=6e-08 w=4.11e-07 $X=33144 $Y=39446 $D=616
M1233 vss 455 443 vss hvtnfet l=6e-08 w=2.74e-07 $X=33254 $Y=13476 $D=616
M1234 b_pxba_n<3> 451 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=33300 $Y=336 $D=616
M1235 451 452 vss vss hvtnfet l=6e-08 w=5e-07 $X=33300 $Y=6701 $D=616
M1236 452 425 vss vss hvtnfet l=6e-08 w=3e-07 $X=33300 $Y=7831 $D=616
M1237 453 425 vss vss hvtnfet l=6e-08 w=3e-07 $X=33300 $Y=43002 $D=616
M1238 454 453 vss vss hvtnfet l=6e-08 w=5e-07 $X=33300 $Y=43932 $D=616
M1239 t_pxba_n<3> 454 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=33300 $Y=49512 $D=616
M1240 vss 368 dwla<1> vss hvtnfet l=6e-08 w=3e-07 $X=33301 $Y=31098 $D=616
M1241 vss 456 497 vss hvtnfet l=6e-08 w=3e-07 $X=33301 $Y=37457 $D=616
M1242 vss 311 1093 vss hvtnfet l=6e-08 w=4.11e-07 $X=33404 $Y=11276 $D=616
M1243 vss 311 1094 vss hvtnfet l=6e-08 w=4.11e-07 $X=33404 $Y=39446 $D=616
M1244 455 aa<8> vss vss hvtnfet l=6e-08 w=2.74e-07 $X=33514 $Y=13476 $D=616
M1245 vss 451 b_pxba_n<3> vss hvtnfet l=6e-08 w=1.285e-06 $X=33560 $Y=336 $D=616
M1246 vss 452 451 vss hvtnfet l=6e-08 w=5e-07 $X=33560 $Y=6701 $D=616
M1247 vss 425 452 vss hvtnfet l=6e-08 w=3e-07 $X=33560 $Y=7831 $D=616
M1248 vss 425 453 vss hvtnfet l=6e-08 w=3e-07 $X=33560 $Y=43002 $D=616
M1249 vss 453 454 vss hvtnfet l=6e-08 w=5e-07 $X=33560 $Y=43932 $D=616
M1250 vss 454 t_pxba_n<3> vss hvtnfet l=6e-08 w=1.285e-06 $X=33560 $Y=49512 $D=616
M1251 dwla<0> 368 vss vss hvtnfet l=6e-08 w=3e-07 $X=33811 $Y=31098 $D=616
M1252 498 456 vss vss hvtnfet l=6e-08 w=3e-07 $X=33811 $Y=37457 $D=616
M1253 555 458 vss vss hvtnfet l=6e-08 w=2e-07 $X=33914 $Y=11276 $D=616
M1254 559 459 vss vss hvtnfet l=6e-08 w=2e-07 $X=33914 $Y=39657 $D=616
M1255 b_pxba_n<2> 460 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=34070 $Y=336 $D=616
M1256 460 461 vss vss hvtnfet l=6e-08 w=5e-07 $X=34070 $Y=6701 $D=616
M1257 461 424 vss vss hvtnfet l=6e-08 w=3e-07 $X=34070 $Y=7831 $D=616
M1258 462 424 vss vss hvtnfet l=6e-08 w=3e-07 $X=34070 $Y=43002 $D=616
M1259 463 462 vss vss hvtnfet l=6e-08 w=5e-07 $X=34070 $Y=43932 $D=616
M1260 t_pxba_n<2> 463 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=34070 $Y=49512 $D=616
M1261 vss 368 dwla<0> vss hvtnfet l=6e-08 w=3e-07 $X=34071 $Y=31098 $D=616
M1262 vss 456 498 vss hvtnfet l=6e-08 w=3e-07 $X=34071 $Y=37457 $D=616
M1263 vss 460 b_pxba_n<2> vss hvtnfet l=6e-08 w=1.285e-06 $X=34330 $Y=336 $D=616
M1264 vss 461 460 vss hvtnfet l=6e-08 w=5e-07 $X=34330 $Y=6701 $D=616
M1265 vss 424 461 vss hvtnfet l=6e-08 w=3e-07 $X=34330 $Y=7831 $D=616
M1266 vss 424 462 vss hvtnfet l=6e-08 w=3e-07 $X=34330 $Y=43002 $D=616
M1267 vss 462 463 vss hvtnfet l=6e-08 w=5e-07 $X=34330 $Y=43932 $D=616
M1268 vss 463 t_pxba_n<2> vss hvtnfet l=6e-08 w=1.285e-06 $X=34330 $Y=49512 $D=616
M1269 1095 449 479 vss hvtnfet l=6e-08 w=5.49e-07 $X=34479 $Y=17417 $D=616
M1270 1096 450 480 vss hvtnfet l=6e-08 w=5.49e-07 $X=34479 $Y=18966 $D=616
M1271 1097 449 481 vss hvtnfet l=6e-08 w=5.49e-07 $X=34479 $Y=24337 $D=616
M1272 1098 450 482 vss hvtnfet l=6e-08 w=5.49e-07 $X=34479 $Y=25886 $D=616
M1273 vss aa<9> 440 vss hvtnfet l=6e-08 w=2.74e-07 $X=34524 $Y=13476 $D=616
M1274 dwla<0> 465 vss vss hvtnfet l=6e-08 w=3e-07 $X=34581 $Y=31098 $D=616
M1275 498 465 vss vss hvtnfet l=6e-08 w=3e-07 $X=34581 $Y=37457 $D=616
M1276 1099 vdd vss vss hvtnfet l=6e-08 w=6.4e-07 $X=34621 $Y=32508 $D=616
M1277 123 131 vss vss hvtnfet l=6e-08 w=2e-07 $X=34646 $Y=11546 $D=616
M1278 1100 455 1095 vss hvtnfet l=6e-08 w=5.49e-07 $X=34739 $Y=17417 $D=616
M1279 1101 455 1096 vss hvtnfet l=6e-08 w=5.49e-07 $X=34739 $Y=18966 $D=616
M1280 1102 455 1097 vss hvtnfet l=6e-08 w=5.49e-07 $X=34739 $Y=24337 $D=616
M1281 1103 455 1098 vss hvtnfet l=6e-08 w=5.49e-07 $X=34739 $Y=25886 $D=616
M1282 b_pxba_n<1> 466 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=34840 $Y=336 $D=616
M1283 466 467 vss vss hvtnfet l=6e-08 w=5e-07 $X=34840 $Y=6701 $D=616
M1284 467 468 vss vss hvtnfet l=6e-08 w=3e-07 $X=34840 $Y=7831 $D=616
M1285 469 468 vss vss hvtnfet l=6e-08 w=3e-07 $X=34840 $Y=43002 $D=616
M1286 470 469 vss vss hvtnfet l=6e-08 w=5e-07 $X=34840 $Y=43932 $D=616
M1287 t_pxba_n<1> 470 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=34840 $Y=49512 $D=616
M1288 vss 465 dwla<0> vss hvtnfet l=6e-08 w=3e-07 $X=34841 $Y=31098 $D=616
M1289 vss 465 498 vss hvtnfet l=6e-08 w=3e-07 $X=34841 $Y=37457 $D=616
M1290 535 471 1099 vss hvtnfet l=6e-08 w=6.4e-07 $X=34881 $Y=32508 $D=616
M1291 vss 123 123 vss hvtnfet l=6e-08 w=2e-07 $X=34906 $Y=11546 $D=616
M1292 1104 439 1100 vss hvtnfet l=6e-08 w=5.49e-07 $X=34999 $Y=17417 $D=616
M1293 1105 439 1101 vss hvtnfet l=6e-08 w=5.49e-07 $X=34999 $Y=18966 $D=616
M1294 1106 440 1102 vss hvtnfet l=6e-08 w=5.49e-07 $X=34999 $Y=24337 $D=616
M1295 1107 440 1103 vss hvtnfet l=6e-08 w=5.49e-07 $X=34999 $Y=25886 $D=616
M1296 439 440 vss vss hvtnfet l=6e-08 w=2.74e-07 $X=35034 $Y=13476 $D=616
M1297 vss 466 b_pxba_n<1> vss hvtnfet l=6e-08 w=1.285e-06 $X=35100 $Y=336 $D=616
M1298 vss 467 466 vss hvtnfet l=6e-08 w=5e-07 $X=35100 $Y=6701 $D=616
M1299 vss 468 467 vss hvtnfet l=6e-08 w=3e-07 $X=35100 $Y=7831 $D=616
M1300 vss 468 469 vss hvtnfet l=6e-08 w=3e-07 $X=35100 $Y=43002 $D=616
M1301 vss 469 470 vss hvtnfet l=6e-08 w=5e-07 $X=35100 $Y=43932 $D=616
M1302 vss 470 t_pxba_n<1> vss hvtnfet l=6e-08 w=1.285e-06 $X=35100 $Y=49512 $D=616
M1303 vss 323 1104 vss hvtnfet l=6e-08 w=8.23e-07 $X=35269 $Y=17143 $D=616
M1304 vss 323 1105 vss hvtnfet l=6e-08 w=8.23e-07 $X=35269 $Y=18966 $D=616
M1305 vss 323 1106 vss hvtnfet l=6e-08 w=8.23e-07 $X=35269 $Y=24063 $D=616
M1306 vss 323 1107 vss hvtnfet l=6e-08 w=8.23e-07 $X=35269 $Y=25886 $D=616
M1307 vss 473 484 vss hvtnfet l=6e-08 w=3e-07 $X=35351 $Y=37257 $D=616
M1308 vss 472 471 vss hvtnfet l=6e-08 w=3.5e-07 $X=35446 $Y=32613 $D=616
M1309 b_pxba_n<0> 474 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=35610 $Y=336 $D=616
M1310 474 475 vss vss hvtnfet l=6e-08 w=5e-07 $X=35610 $Y=6701 $D=616
M1311 475 476 vss vss hvtnfet l=6e-08 w=3e-07 $X=35610 $Y=7831 $D=616
M1312 477 476 vss vss hvtnfet l=6e-08 w=3e-07 $X=35610 $Y=43002 $D=616
M1313 478 477 vss vss hvtnfet l=6e-08 w=5e-07 $X=35610 $Y=43932 $D=616
M1314 t_pxba_n<0> 478 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=35610 $Y=49512 $D=616
M1315 472 483 vss vss hvtnfet l=2.5e-07 w=3.5e-07 $X=35706 $Y=32613 $D=616
M1316 446 479 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=35764 $Y=17812 $D=616
M1317 434 480 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=35764 $Y=18983 $D=616
M1318 476 481 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=35764 $Y=24732 $D=616
M1319 468 482 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=35764 $Y=25903 $D=616
M1320 1108 317 479 vss hvtnfet l=6e-08 w=1.8e-07 $X=35779 $Y=17143 $D=616
M1321 1109 317 480 vss hvtnfet l=6e-08 w=1.8e-07 $X=35779 $Y=19609 $D=616
M1322 1110 317 481 vss hvtnfet l=6e-08 w=1.8e-07 $X=35779 $Y=24063 $D=616
M1323 1111 317 482 vss hvtnfet l=6e-08 w=1.8e-07 $X=35779 $Y=26529 $D=616
M1324 473 484 vss vss hvtnfet l=1.2e-07 w=1.5e-07 $X=35861 $Y=37297 $D=616
M1325 vss 474 b_pxba_n<0> vss hvtnfet l=6e-08 w=1.285e-06 $X=35870 $Y=336 $D=616
M1326 vss 475 474 vss hvtnfet l=6e-08 w=5e-07 $X=35870 $Y=6701 $D=616
M1327 vss 476 475 vss hvtnfet l=6e-08 w=3e-07 $X=35870 $Y=7831 $D=616
M1328 vss 476 477 vss hvtnfet l=6e-08 w=3e-07 $X=35870 $Y=43002 $D=616
M1329 vss 477 478 vss hvtnfet l=6e-08 w=5e-07 $X=35870 $Y=43932 $D=616
M1330 vss 478 t_pxba_n<0> vss hvtnfet l=6e-08 w=1.285e-06 $X=35870 $Y=49512 $D=616
M1331 773 495 vss vss hvtnfet l=6e-08 w=8e-07 $X=35945 $Y=30668 $D=616
M1332 vss 479 446 vss hvtnfet l=6e-08 w=1.37e-07 $X=36024 $Y=17812 $D=616
M1333 vss 480 434 vss hvtnfet l=6e-08 w=1.37e-07 $X=36024 $Y=18983 $D=616
M1334 vss 481 476 vss hvtnfet l=6e-08 w=1.37e-07 $X=36024 $Y=24732 $D=616
M1335 vss 482 468 vss hvtnfet l=6e-08 w=1.37e-07 $X=36024 $Y=25903 $D=616
M1336 vss 446 1108 vss hvtnfet l=6e-08 w=1.8e-07 $X=36039 $Y=17143 $D=616
M1337 vss 434 1109 vss hvtnfet l=6e-08 w=1.8e-07 $X=36039 $Y=19609 $D=616
M1338 vss 476 1110 vss hvtnfet l=6e-08 w=1.8e-07 $X=36039 $Y=24063 $D=616
M1339 vss 468 1111 vss hvtnfet l=6e-08 w=1.8e-07 $X=36039 $Y=26529 $D=616
M1340 vss 495 773 vss hvtnfet l=6e-08 w=8e-07 $X=36205 $Y=30668 $D=616
M1341 vss 491 509 vss hvtnfet l=6e-08 w=2.74e-07 $X=36254 $Y=13476 $D=616
M1342 b_pxaa<3> 485 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=36380 $Y=336 $D=616
M1343 485 486 vss vss hvtnfet l=6e-08 w=5e-07 $X=36380 $Y=6701 $D=616
M1344 486 487 vss vss hvtnfet l=6e-08 w=3e-07 $X=36380 $Y=7831 $D=616
M1345 1112 492 vss vss hvtnfet l=6e-08 w=4.11e-07 $X=36380 $Y=11276 $D=616
M1346 1113 492 vss vss hvtnfet l=6e-08 w=4.11e-07 $X=36380 $Y=39446 $D=616
M1347 489 488 vss vss hvtnfet l=6e-08 w=3e-07 $X=36380 $Y=43002 $D=616
M1348 490 489 vss vss hvtnfet l=6e-08 w=5e-07 $X=36380 $Y=43932 $D=616
M1349 t_pxaa<3> 490 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=36380 $Y=49512 $D=616
M1350 vss 494 473 vss hvtnfet l=6e-08 w=3.2e-07 $X=36431 $Y=37292 $D=616
M1351 vss 496 483 vss hvtnfet l=6e-08 w=3.2e-07 $X=36466 $Y=32828 $D=616
M1352 vss 485 b_pxaa<3> vss hvtnfet l=6e-08 w=1.285e-06 $X=36640 $Y=336 $D=616
M1353 vss 486 485 vss hvtnfet l=6e-08 w=5e-07 $X=36640 $Y=6701 $D=616
M1354 vss 487 486 vss hvtnfet l=6e-08 w=3e-07 $X=36640 $Y=7831 $D=616
M1355 487 497 1112 vss hvtnfet l=6e-08 w=4.11e-07 $X=36640 $Y=11276 $D=616
M1356 488 498 1113 vss hvtnfet l=6e-08 w=4.11e-07 $X=36640 $Y=39446 $D=616
M1357 vss 488 489 vss hvtnfet l=6e-08 w=3e-07 $X=36640 $Y=43002 $D=616
M1358 vss 489 490 vss hvtnfet l=6e-08 w=5e-07 $X=36640 $Y=43932 $D=616
M1359 vss 490 t_pxaa<3> vss hvtnfet l=6e-08 w=1.285e-06 $X=36640 $Y=49512 $D=616
M1360 368 clka 773 vss hvtnfet l=6e-08 w=8e-07 $X=36715 $Y=30668 $D=616
M1361 491 aa<6> vss vss hvtnfet l=6e-08 w=2.74e-07 $X=36764 $Y=13476 $D=616
M1362 773 clka 368 vss hvtnfet l=6e-08 w=8e-07 $X=36975 $Y=30668 $D=616
M1363 vss 473 496 vss hvtnfet l=6e-08 w=3.2e-07 $X=36976 $Y=32828 $D=616
M1364 1114 501 519 vss hvtnfet l=6e-08 w=5.49e-07 $X=37059 $Y=17143 $D=616
M1365 1115 502 520 vss hvtnfet l=6e-08 w=5.49e-07 $X=37059 $Y=19240 $D=616
M1366 1116 501 521 vss hvtnfet l=6e-08 w=5.49e-07 $X=37059 $Y=24063 $D=616
M1367 1117 502 522 vss hvtnfet l=6e-08 w=5.49e-07 $X=37059 $Y=26160 $D=616
M1368 b_pxaa<2> 503 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=37150 $Y=336 $D=616
M1369 503 504 vss vss hvtnfet l=6e-08 w=5e-07 $X=37150 $Y=6701 $D=616
M1370 504 505 vss vss hvtnfet l=6e-08 w=3e-07 $X=37150 $Y=7831 $D=616
M1371 1118 497 505 vss hvtnfet l=6e-08 w=4.11e-07 $X=37150 $Y=11276 $D=616
M1372 1119 498 506 vss hvtnfet l=6e-08 w=4.11e-07 $X=37150 $Y=39446 $D=616
M1373 507 506 vss vss hvtnfet l=6e-08 w=3e-07 $X=37150 $Y=43002 $D=616
M1374 508 507 vss vss hvtnfet l=6e-08 w=5e-07 $X=37150 $Y=43932 $D=616
M1375 t_pxaa<2> 508 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=37150 $Y=49512 $D=616
M1376 vss ddqa_n 493 vss hvtnfet l=6e-08 w=2.4e-07 $X=37161 $Y=37292 $D=616
M1377 vss 502 501 vss hvtnfet l=6e-08 w=2.74e-07 $X=37274 $Y=13476 $D=616
M1378 1120 509 1114 vss hvtnfet l=6e-08 w=5.49e-07 $X=37319 $Y=17143 $D=616
M1379 1121 509 1115 vss hvtnfet l=6e-08 w=5.49e-07 $X=37319 $Y=19240 $D=616
M1380 1122 491 1116 vss hvtnfet l=6e-08 w=5.49e-07 $X=37319 $Y=24063 $D=616
M1381 1123 491 1117 vss hvtnfet l=6e-08 w=5.49e-07 $X=37319 $Y=26160 $D=616
M1382 vss 503 b_pxaa<2> vss hvtnfet l=6e-08 w=1.285e-06 $X=37410 $Y=336 $D=616
M1383 vss 504 503 vss hvtnfet l=6e-08 w=5e-07 $X=37410 $Y=6701 $D=616
M1384 vss 505 504 vss hvtnfet l=6e-08 w=3e-07 $X=37410 $Y=7831 $D=616
M1385 vss 510 1118 vss hvtnfet l=6e-08 w=4.11e-07 $X=37410 $Y=11276 $D=616
M1386 vss 510 1119 vss hvtnfet l=6e-08 w=4.11e-07 $X=37410 $Y=39446 $D=616
M1387 vss 506 507 vss hvtnfet l=6e-08 w=3e-07 $X=37410 $Y=43002 $D=616
M1388 vss 507 508 vss hvtnfet l=6e-08 w=5e-07 $X=37410 $Y=43932 $D=616
M1389 vss 508 t_pxaa<2> vss hvtnfet l=6e-08 w=1.285e-06 $X=37410 $Y=49512 $D=616
M1390 493 ddqa vss vss hvtnfet l=6e-08 w=2.4e-07 $X=37421 $Y=37292 $D=616
M1391 vss clka 524 vss hvtnfet l=6e-08 w=6e-07 $X=37485 $Y=30668 $D=616
M1392 vss 323 1120 vss hvtnfet l=6e-08 w=8.23e-07 $X=37589 $Y=17143 $D=616
M1393 vss 323 1121 vss hvtnfet l=6e-08 w=8.23e-07 $X=37589 $Y=18966 $D=616
M1394 vss 323 1122 vss hvtnfet l=6e-08 w=8.23e-07 $X=37589 $Y=24063 $D=616
M1395 vss 323 1123 vss hvtnfet l=6e-08 w=8.23e-07 $X=37589 $Y=25886 $D=616
M1396 1124 496 557 vss hvtnfet l=6e-08 w=6.4e-07 $X=37661 $Y=32508 $D=616
M1397 502 aa<5> vss vss hvtnfet l=6e-08 w=2.74e-07 $X=37784 $Y=13476 $D=616
M1398 b_pxaa<1> 512 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=37920 $Y=336 $D=616
M1399 512 513 vss vss hvtnfet l=6e-08 w=5e-07 $X=37920 $Y=6701 $D=616
M1400 513 514 vss vss hvtnfet l=6e-08 w=3e-07 $X=37920 $Y=7831 $D=616
M1401 1125 523 vss vss hvtnfet l=6e-08 w=4.11e-07 $X=37920 $Y=11276 $D=616
M1402 1126 523 vss vss hvtnfet l=6e-08 w=4.11e-07 $X=37920 $Y=39446 $D=616
M1403 516 515 vss vss hvtnfet l=6e-08 w=3e-07 $X=37920 $Y=43002 $D=616
M1404 517 516 vss vss hvtnfet l=6e-08 w=5e-07 $X=37920 $Y=43932 $D=616
M1405 t_pxaa<1> 517 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=37920 $Y=49512 $D=616
M1406 vss 386 1124 vss hvtnfet l=6e-08 w=6.4e-07 $X=37921 $Y=32508 $D=616
M1407 1127 317 519 vss hvtnfet l=6e-08 w=1.8e-07 $X=38099 $Y=17143 $D=616
M1408 492 519 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=38099 $Y=17812 $D=616
M1409 510 520 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=38099 $Y=18983 $D=616
M1410 1128 317 520 vss hvtnfet l=6e-08 w=1.8e-07 $X=38099 $Y=19609 $D=616
M1411 1129 317 521 vss hvtnfet l=6e-08 w=1.8e-07 $X=38099 $Y=24063 $D=616
M1412 523 521 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=38099 $Y=24732 $D=616
M1413 525 522 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=38099 $Y=25903 $D=616
M1414 1130 317 522 vss hvtnfet l=6e-08 w=1.8e-07 $X=38099 $Y=26529 $D=616
M1415 vss 493 526 vss hvtnfet l=1.4e-07 w=3.2e-07 $X=38141 $Y=37127 $D=616
M1416 vss 512 b_pxaa<1> vss hvtnfet l=6e-08 w=1.285e-06 $X=38180 $Y=336 $D=616
M1417 vss 513 512 vss hvtnfet l=6e-08 w=5e-07 $X=38180 $Y=6701 $D=616
M1418 vss 514 513 vss hvtnfet l=6e-08 w=3e-07 $X=38180 $Y=7831 $D=616
M1419 514 497 1125 vss hvtnfet l=6e-08 w=4.11e-07 $X=38180 $Y=11276 $D=616
M1420 515 498 1126 vss hvtnfet l=6e-08 w=4.11e-07 $X=38180 $Y=39446 $D=616
M1421 vss 515 516 vss hvtnfet l=6e-08 w=3e-07 $X=38180 $Y=43002 $D=616
M1422 vss 516 517 vss hvtnfet l=6e-08 w=5e-07 $X=38180 $Y=43932 $D=616
M1423 vss 517 t_pxaa<1> vss hvtnfet l=6e-08 w=1.285e-06 $X=38180 $Y=49512 $D=616
M1424 vss 524 534 vss hvtnfet l=6e-08 w=5.49e-07 $X=38255 $Y=30668 $D=616
M1425 vss 492 1127 vss hvtnfet l=6e-08 w=1.8e-07 $X=38359 $Y=17143 $D=616
M1426 vss 519 492 vss hvtnfet l=6e-08 w=1.37e-07 $X=38359 $Y=17812 $D=616
M1427 vss 520 510 vss hvtnfet l=6e-08 w=1.37e-07 $X=38359 $Y=18983 $D=616
M1428 vss 510 1128 vss hvtnfet l=6e-08 w=1.8e-07 $X=38359 $Y=19609 $D=616
M1429 vss 523 1129 vss hvtnfet l=6e-08 w=1.8e-07 $X=38359 $Y=24063 $D=616
M1430 vss 521 523 vss hvtnfet l=6e-08 w=1.37e-07 $X=38359 $Y=24732 $D=616
M1431 vss 522 525 vss hvtnfet l=6e-08 w=1.37e-07 $X=38359 $Y=25903 $D=616
M1432 vss 525 1130 vss hvtnfet l=6e-08 w=1.8e-07 $X=38359 $Y=26529 $D=616
M1433 779 494 vss vss hvtnfet l=6e-08 w=3.2e-07 $X=38431 $Y=32828 $D=616
M1434 780 526 vss vss hvtnfet l=1.4e-07 w=3.2e-07 $X=38481 $Y=37127 $D=616
M1435 534 495 vss vss hvtnfet l=6e-08 w=5.49e-07 $X=38515 $Y=30668 $D=616
M1436 vss 533 546 vss hvtnfet l=6e-08 w=2.74e-07 $X=38574 $Y=13476 $D=616
M1437 b_pxaa<0> 527 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=38690 $Y=336 $D=616
M1438 527 528 vss vss hvtnfet l=6e-08 w=5e-07 $X=38690 $Y=6701 $D=616
M1439 528 529 vss vss hvtnfet l=6e-08 w=3e-07 $X=38690 $Y=7831 $D=616
M1440 1131 497 529 vss hvtnfet l=6e-08 w=4.11e-07 $X=38690 $Y=11276 $D=616
M1441 1132 498 530 vss hvtnfet l=6e-08 w=4.11e-07 $X=38690 $Y=39446 $D=616
M1442 531 530 vss vss hvtnfet l=6e-08 w=3e-07 $X=38690 $Y=43002 $D=616
M1443 532 531 vss vss hvtnfet l=6e-08 w=5e-07 $X=38690 $Y=43932 $D=616
M1444 t_pxaa<0> 532 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=38690 $Y=49512 $D=616
M1445 vss 527 b_pxaa<0> vss hvtnfet l=6e-08 w=1.285e-06 $X=38950 $Y=336 $D=616
M1446 vss 528 527 vss hvtnfet l=6e-08 w=5e-07 $X=38950 $Y=6701 $D=616
M1447 vss 529 528 vss hvtnfet l=6e-08 w=3e-07 $X=38950 $Y=7831 $D=616
M1448 vss 525 1131 vss hvtnfet l=6e-08 w=4.11e-07 $X=38950 $Y=11276 $D=616
M1449 vss 525 1132 vss hvtnfet l=6e-08 w=4.11e-07 $X=38950 $Y=39446 $D=616
M1450 vss 530 531 vss hvtnfet l=6e-08 w=3e-07 $X=38950 $Y=43002 $D=616
M1451 vss 531 532 vss hvtnfet l=6e-08 w=5e-07 $X=38950 $Y=43932 $D=616
M1452 vss 532 t_pxaa<0> vss hvtnfet l=6e-08 w=1.285e-06 $X=38950 $Y=49512 $D=616
M1453 vss 534 495 vss hvtnfet l=6e-08 w=5.49e-07 $X=39025 $Y=30668 $D=616
M1454 533 aa<3> vss vss hvtnfet l=6e-08 w=2.74e-07 $X=39084 $Y=13476 $D=616
M1455 vss clka 323 vss hvtnfet l=6e-08 w=6e-07 $X=39174 $Y=32403 $D=616
M1456 293 535 vss vss hvtnfet l=6e-08 w=6e-07 $X=39185 $Y=37277 $D=616
M1457 495 539 vss vss hvtnfet l=6e-08 w=5.49e-07 $X=39285 $Y=30668 $D=616
M1458 1133 537 549 vss hvtnfet l=6e-08 w=5.49e-07 $X=39379 $Y=17143 $D=616
M1459 1134 538 550 vss hvtnfet l=6e-08 w=5.49e-07 $X=39379 $Y=19240 $D=616
M1460 1135 537 551 vss hvtnfet l=6e-08 w=5.49e-07 $X=39379 $Y=24063 $D=616
M1461 1136 538 552 vss hvtnfet l=6e-08 w=5.49e-07 $X=39379 $Y=26160 $D=616
M1462 323 clka vss vss hvtnfet l=6e-08 w=6e-07 $X=39434 $Y=32403 $D=616
M1463 vss 538 537 vss hvtnfet l=6e-08 w=2.74e-07 $X=39594 $Y=13476 $D=616
M1464 1137 546 1133 vss hvtnfet l=6e-08 w=5.49e-07 $X=39639 $Y=17143 $D=616
M1465 1138 546 1134 vss hvtnfet l=6e-08 w=5.49e-07 $X=39639 $Y=19240 $D=616
M1466 1139 533 1135 vss hvtnfet l=6e-08 w=5.49e-07 $X=39639 $Y=24063 $D=616
M1467 1140 533 1136 vss hvtnfet l=6e-08 w=5.49e-07 $X=39639 $Y=26160 $D=616
M1468 r_sa_prea_n 293 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=39695 $Y=37027 $D=616
M1469 289 540 vss vss hvtnfet l=6e-08 w=6e-07 $X=39705 $Y=336 $D=616
M1470 290 541 vss vss hvtnfet l=6e-08 w=6e-07 $X=39705 $Y=5566 $D=616
M1471 291 542 vss vss hvtnfet l=6e-08 w=6e-07 $X=39705 $Y=6796 $D=616
M1472 292 543 vss vss hvtnfet l=6e-08 w=6e-07 $X=39705 $Y=12026 $D=616
M1473 294 543 vss vss hvtnfet l=6e-08 w=6e-07 $X=39705 $Y=38507 $D=616
M1474 295 542 vss vss hvtnfet l=6e-08 w=6e-07 $X=39705 $Y=43737 $D=616
M1475 296 544 vss vss hvtnfet l=6e-08 w=6e-07 $X=39705 $Y=44967 $D=616
M1476 297 545 vss vss hvtnfet l=6e-08 w=6e-07 $X=39705 $Y=50197 $D=616
M1477 vss stclka 539 vss hvtnfet l=6e-08 w=2.74e-07 $X=39795 $Y=30668 $D=616
M1478 vss 323 1137 vss hvtnfet l=6e-08 w=8.23e-07 $X=39909 $Y=17143 $D=616
M1479 vss 323 1138 vss hvtnfet l=6e-08 w=8.23e-07 $X=39909 $Y=18966 $D=616
M1480 vss 323 1139 vss hvtnfet l=6e-08 w=8.23e-07 $X=39909 $Y=24063 $D=616
M1481 vss 323 1140 vss hvtnfet l=6e-08 w=8.23e-07 $X=39909 $Y=25886 $D=616
M1482 vss 293 r_sa_prea_n vss hvtnfet l=6e-08 w=8.58e-07 $X=39955 $Y=37027 $D=616
M1483 538 aa<2> vss vss hvtnfet l=6e-08 w=2.74e-07 $X=40104 $Y=13476 $D=616
M1484 rb_ca<1> 289 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=40215 $Y=328 $D=616
M1485 rb_ca<3> 290 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=40215 $Y=5316 $D=616
M1486 rb_ma<1> 291 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=40215 $Y=6788 $D=616
M1487 rb_ma<3> 292 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=40215 $Y=11776 $D=616
M1488 r_sa_prea_n 293 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=40215 $Y=37027 $D=616
M1489 rt_ma<3> 294 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=40215 $Y=38499 $D=616
M1490 rt_ma<1> 295 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=40215 $Y=43487 $D=616
M1491 rt_ca<3> 296 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=40215 $Y=44959 $D=616
M1492 rt_ca<1> 297 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=40215 $Y=49947 $D=616
M1493 1141 317 549 vss hvtnfet l=6e-08 w=1.8e-07 $X=40419 $Y=17143 $D=616
M1494 543 549 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=40419 $Y=17812 $D=616
M1495 553 550 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=40419 $Y=18983 $D=616
M1496 1142 317 550 vss hvtnfet l=6e-08 w=1.8e-07 $X=40419 $Y=19609 $D=616
M1497 1143 317 551 vss hvtnfet l=6e-08 w=1.8e-07 $X=40419 $Y=24063 $D=616
M1498 542 551 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=40419 $Y=24732 $D=616
M1499 554 552 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=40419 $Y=25903 $D=616
M1500 1144 317 552 vss hvtnfet l=6e-08 w=1.8e-07 $X=40419 $Y=26529 $D=616
M1501 vss 289 rb_ca<1> vss hvtnfet l=6e-08 w=8.58e-07 $X=40475 $Y=328 $D=616
M1502 vss 290 rb_ca<3> vss hvtnfet l=6e-08 w=8.58e-07 $X=40475 $Y=5316 $D=616
M1503 vss 291 rb_ma<1> vss hvtnfet l=6e-08 w=8.58e-07 $X=40475 $Y=6788 $D=616
M1504 vss 292 rb_ma<3> vss hvtnfet l=6e-08 w=8.58e-07 $X=40475 $Y=11776 $D=616
M1505 vss 294 rt_ma<3> vss hvtnfet l=6e-08 w=8.58e-07 $X=40475 $Y=38499 $D=616
M1506 vss 295 rt_ma<1> vss hvtnfet l=6e-08 w=8.58e-07 $X=40475 $Y=43487 $D=616
M1507 vss 296 rt_ca<3> vss hvtnfet l=6e-08 w=8.58e-07 $X=40475 $Y=44959 $D=616
M1508 vss 297 rt_ca<1> vss hvtnfet l=6e-08 w=8.58e-07 $X=40475 $Y=49947 $D=616
M1509 vss 543 1141 vss hvtnfet l=6e-08 w=1.8e-07 $X=40679 $Y=17143 $D=616
M1510 vss 549 543 vss hvtnfet l=6e-08 w=1.37e-07 $X=40679 $Y=17812 $D=616
M1511 vss 550 553 vss hvtnfet l=6e-08 w=1.37e-07 $X=40679 $Y=18983 $D=616
M1512 vss 553 1142 vss hvtnfet l=6e-08 w=1.8e-07 $X=40679 $Y=19609 $D=616
M1513 vss 542 1143 vss hvtnfet l=6e-08 w=1.8e-07 $X=40679 $Y=24063 $D=616
M1514 vss 551 542 vss hvtnfet l=6e-08 w=1.37e-07 $X=40679 $Y=24732 $D=616
M1515 vss 552 554 vss hvtnfet l=6e-08 w=1.37e-07 $X=40679 $Y=25903 $D=616
M1516 vss 554 1144 vss hvtnfet l=6e-08 w=1.8e-07 $X=40679 $Y=26529 $D=616
M1517 vss 303 r_saea_n vss hvtnfet l=6e-08 w=8.58e-07 $X=40725 $Y=37027 $D=616
M1518 rb_ca<1> 289 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=40735 $Y=328 $D=616
M1519 rb_ca<3> 290 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=40735 $Y=5316 $D=616
M1520 rb_ma<1> 291 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=40735 $Y=6788 $D=616
M1521 rb_ma<3> 292 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=40735 $Y=11776 $D=616
M1522 rt_ma<3> 294 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=40735 $Y=38499 $D=616
M1523 rt_ma<1> 295 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=40735 $Y=43487 $D=616
M1524 rt_ca<3> 296 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=40735 $Y=44959 $D=616
M1525 rt_ca<1> 297 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=40735 $Y=49947 $D=616
M1526 r_saea_n 303 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=40985 $Y=37027 $D=616
M1527 vss 299 rb_ca<0> vss hvtnfet l=6e-08 w=8.58e-07 $X=41245 $Y=328 $D=616
M1528 vss 300 rb_ca<2> vss hvtnfet l=6e-08 w=8.58e-07 $X=41245 $Y=5316 $D=616
M1529 vss 301 rb_ma<0> vss hvtnfet l=6e-08 w=8.58e-07 $X=41245 $Y=6788 $D=616
M1530 vss 302 rb_ma<2> vss hvtnfet l=6e-08 w=8.58e-07 $X=41245 $Y=11776 $D=616
M1531 vss 303 r_saea_n vss hvtnfet l=6e-08 w=8.58e-07 $X=41245 $Y=37027 $D=616
M1532 vss 304 rt_ma<2> vss hvtnfet l=6e-08 w=8.58e-07 $X=41245 $Y=38499 $D=616
M1533 vss 305 rt_ma<0> vss hvtnfet l=6e-08 w=8.58e-07 $X=41245 $Y=43487 $D=616
M1534 vss 306 rt_ca<2> vss hvtnfet l=6e-08 w=8.58e-07 $X=41245 $Y=44959 $D=616
M1535 vss 307 rt_ca<0> vss hvtnfet l=6e-08 w=8.58e-07 $X=41245 $Y=49947 $D=616
M1536 vss clka 287 vss hvtnfet l=6e-08 w=1.05e-06 $X=41495 $Y=22251 $D=616
M1537 vss 340 288 vss hvtnfet l=6e-08 w=1.05e-06 $X=41495 $Y=29007 $D=616
M1538 rb_ca<0> 299 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=41505 $Y=328 $D=616
M1539 rb_ca<2> 300 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=41505 $Y=5316 $D=616
M1540 rb_ma<0> 301 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=41505 $Y=6788 $D=616
M1541 rb_ma<2> 302 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=41505 $Y=11776 $D=616
M1542 285 497 vss vss hvtnfet l=6e-08 w=6e-07 $X=41505 $Y=13282 $D=616
M1543 286 498 vss vss hvtnfet l=6e-08 w=6e-07 $X=41505 $Y=20809 $D=616
M1544 r_saea_n 303 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=41505 $Y=37027 $D=616
M1545 rt_ma<2> 304 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=41505 $Y=38499 $D=616
M1546 rt_ma<0> 305 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=41505 $Y=43487 $D=616
M1547 rt_ca<2> 306 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=41505 $Y=44959 $D=616
M1548 rt_ca<0> 307 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=41505 $Y=49947 $D=616
M1549 r_clk_dqa 287 vss vss hvtnfet l=6e-08 w=1.26e-06 $X=41755 $Y=22041 $D=616
M1550 r_clk_dqa_n 288 vss vss hvtnfet l=6e-08 w=1.26e-06 $X=41755 $Y=29007 $D=616
M1551 vss 299 rb_ca<0> vss hvtnfet l=6e-08 w=8.58e-07 $X=41765 $Y=328 $D=616
M1552 vss 300 rb_ca<2> vss hvtnfet l=6e-08 w=8.58e-07 $X=41765 $Y=5316 $D=616
M1553 vss 301 rb_ma<0> vss hvtnfet l=6e-08 w=8.58e-07 $X=41765 $Y=6788 $D=616
M1554 vss 302 rb_ma<2> vss hvtnfet l=6e-08 w=8.58e-07 $X=41765 $Y=11776 $D=616
M1555 vss 303 r_saea_n vss hvtnfet l=6e-08 w=8.58e-07 $X=41765 $Y=37027 $D=616
M1556 vss 304 rt_ma<2> vss hvtnfet l=6e-08 w=8.58e-07 $X=41765 $Y=38499 $D=616
M1557 vss 305 rt_ma<0> vss hvtnfet l=6e-08 w=8.58e-07 $X=41765 $Y=43487 $D=616
M1558 vss 306 rt_ca<2> vss hvtnfet l=6e-08 w=8.58e-07 $X=41765 $Y=44959 $D=616
M1559 vss 307 rt_ca<0> vss hvtnfet l=6e-08 w=8.58e-07 $X=41765 $Y=49947 $D=616
M1560 rb_tm_prea_n 285 vss vss hvtnfet l=6e-08 w=1.287e-06 $X=42015 $Y=13280 $D=616
M1561 rt_tm_prea_n 286 vss vss hvtnfet l=6e-08 w=1.287e-06 $X=42015 $Y=20124 $D=616
M1562 vss 287 r_clk_dqa vss hvtnfet l=6e-08 w=1.26e-06 $X=42015 $Y=22041 $D=616
M1563 vss 288 r_clk_dqa_n vss hvtnfet l=6e-08 w=1.26e-06 $X=42015 $Y=29007 $D=616
M1564 r_lwea 284 vss vss hvtnfet l=6e-08 w=1.287e-06 $X=42015 $Y=30897 $D=616
M1565 vss 555 299 vss hvtnfet l=6e-08 w=6e-07 $X=42275 $Y=336 $D=616
M1566 vss 556 300 vss hvtnfet l=6e-08 w=6e-07 $X=42275 $Y=5566 $D=616
M1567 vss 554 301 vss hvtnfet l=6e-08 w=6e-07 $X=42275 $Y=6796 $D=616
M1568 vss 553 302 vss hvtnfet l=6e-08 w=6e-07 $X=42275 $Y=12026 $D=616
M1569 vss 285 rb_tm_prea_n vss hvtnfet l=6e-08 w=1.287e-06 $X=42275 $Y=13280 $D=616
M1570 vss 286 rt_tm_prea_n vss hvtnfet l=6e-08 w=1.287e-06 $X=42275 $Y=20124 $D=616
M1571 r_clk_dqa 287 vss vss hvtnfet l=6e-08 w=1.26e-06 $X=42275 $Y=22041 $D=616
M1572 r_clk_dqa_n 288 vss vss hvtnfet l=6e-08 w=1.26e-06 $X=42275 $Y=29007 $D=616
M1573 vss 284 r_lwea vss hvtnfet l=6e-08 w=1.287e-06 $X=42275 $Y=30897 $D=616
M1574 vss 557 303 vss hvtnfet l=6e-08 w=6e-07 $X=42275 $Y=37277 $D=616
M1575 vss 553 304 vss hvtnfet l=6e-08 w=6e-07 $X=42275 $Y=38507 $D=616
M1576 vss 554 305 vss hvtnfet l=6e-08 w=6e-07 $X=42275 $Y=43737 $D=616
M1577 vss 558 306 vss hvtnfet l=6e-08 w=6e-07 $X=42275 $Y=44967 $D=616
M1578 vss 559 307 vss hvtnfet l=6e-08 w=6e-07 $X=42275 $Y=50197 $D=616
M1579 303 557 vss vss hvtnfet l=6e-08 w=6e-07 $X=42535 $Y=37277 $D=616
M1580 vdd 5 15 vdd hvtpfet l=6e-08 w=1.2e-06 $X=965 $Y=35277 $D=636
M1581 11 1 vdd vdd hvtpfet l=6e-08 w=1.2e-06 $X=1225 $Y=1736 $D=636
M1582 12 2 vdd vdd hvtpfet l=6e-08 w=1.2e-06 $X=1225 $Y=3566 $D=636
M1583 13 3 vdd vdd hvtpfet l=6e-08 w=1.2e-06 $X=1225 $Y=8196 $D=636
M1584 14 4 vdd vdd hvtpfet l=6e-08 w=1.2e-06 $X=1225 $Y=10026 $D=636
M1585 lb_tm_preb_n 20 vdd vdd hvtpfet l=6e-08 w=2.145e-06 $X=1225 $Y=14887 $D=636
M1586 lt_tm_preb_n 21 vdd vdd hvtpfet l=6e-08 w=2.145e-06 $X=1225 $Y=17659 $D=636
M1587 vdd 8 l_clk_dqb vdd hvtpfet l=6e-08 w=2.1e-06 $X=1225 $Y=23621 $D=636
M1588 vdd 9 l_clk_dqb_n vdd hvtpfet l=6e-08 w=2.1e-06 $X=1225 $Y=26587 $D=636
M1589 l_lweb 10 vdd vdd hvtpfet l=6e-08 w=2.145e-06 $X=1225 $Y=32504 $D=636
M1590 15 5 vdd vdd hvtpfet l=6e-08 w=1.2e-06 $X=1225 $Y=35277 $D=636
M1591 16 4 vdd vdd hvtpfet l=6e-08 w=1.2e-06 $X=1225 $Y=39907 $D=636
M1592 17 3 vdd vdd hvtpfet l=6e-08 w=1.2e-06 $X=1225 $Y=41737 $D=636
M1593 18 6 vdd vdd hvtpfet l=6e-08 w=1.2e-06 $X=1225 $Y=46367 $D=636
M1594 19 7 vdd vdd hvtpfet l=6e-08 w=1.2e-06 $X=1225 $Y=48197 $D=636
M1595 vdd 20 lb_tm_preb_n vdd hvtpfet l=6e-08 w=2.145e-06 $X=1485 $Y=14887 $D=636
M1596 vdd 21 lt_tm_preb_n vdd hvtpfet l=6e-08 w=2.145e-06 $X=1485 $Y=17659 $D=636
M1597 l_clk_dqb 8 vdd vdd hvtpfet l=6e-08 w=2.1e-06 $X=1485 $Y=23621 $D=636
M1598 l_clk_dqb_n 9 vdd vdd hvtpfet l=6e-08 w=2.1e-06 $X=1485 $Y=26587 $D=636
M1599 vdd 10 l_lweb vdd hvtpfet l=6e-08 w=2.145e-06 $X=1485 $Y=32504 $D=636
M1600 lb_cb<0> 11 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=1735 $Y=1506 $D=636
M1601 lb_cb<2> 12 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=1735 $Y=3566 $D=636
M1602 lb_mb<0> 13 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=1735 $Y=7966 $D=636
M1603 lb_mb<2> 14 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=1735 $Y=10026 $D=636
M1604 l_saeb_n 15 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=1735 $Y=35277 $D=636
M1605 lt_mb<2> 16 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=1735 $Y=39677 $D=636
M1606 lt_mb<0> 17 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=1735 $Y=41737 $D=636
M1607 lt_cb<2> 18 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=1735 $Y=46137 $D=636
M1608 lt_cb<0> 19 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=1735 $Y=48197 $D=636
M1609 vdd 8 l_clk_dqb vdd hvtpfet l=6e-08 w=2.1e-06 $X=1745 $Y=23621 $D=636
M1610 vdd 9 l_clk_dqb_n vdd hvtpfet l=6e-08 w=2.1e-06 $X=1745 $Y=26587 $D=636
M1611 vdd 11 lb_cb<0> vdd hvtpfet l=6e-08 w=1.43e-06 $X=1995 $Y=1506 $D=636
M1612 vdd 12 lb_cb<2> vdd hvtpfet l=6e-08 w=1.43e-06 $X=1995 $Y=3566 $D=636
M1613 vdd 13 lb_mb<0> vdd hvtpfet l=6e-08 w=1.43e-06 $X=1995 $Y=7966 $D=636
M1614 vdd 14 lb_mb<2> vdd hvtpfet l=6e-08 w=1.43e-06 $X=1995 $Y=10026 $D=636
M1615 vdd 24 20 vdd hvtpfet l=6e-08 w=1.2e-06 $X=1995 $Y=15067 $D=636
M1616 vdd 25 21 vdd hvtpfet l=6e-08 w=1.2e-06 $X=1995 $Y=18424 $D=636
M1617 vdd 15 l_saeb_n vdd hvtpfet l=6e-08 w=1.43e-06 $X=1995 $Y=35277 $D=636
M1618 vdd 16 lt_mb<2> vdd hvtpfet l=6e-08 w=1.43e-06 $X=1995 $Y=39677 $D=636
M1619 vdd 17 lt_mb<0> vdd hvtpfet l=6e-08 w=1.43e-06 $X=1995 $Y=41737 $D=636
M1620 vdd 18 lt_cb<2> vdd hvtpfet l=6e-08 w=1.43e-06 $X=1995 $Y=46137 $D=636
M1621 vdd 19 lt_cb<0> vdd hvtpfet l=6e-08 w=1.43e-06 $X=1995 $Y=48197 $D=636
M1622 8 clkb vdd vdd hvtpfet l=6e-08 w=2.1e-06 $X=2005 $Y=23621 $D=636
M1623 9 23 vdd vdd hvtpfet l=6e-08 w=2.1e-06 $X=2005 $Y=26587 $D=636
M1624 lb_cb<0> 11 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=2255 $Y=1506 $D=636
M1625 lb_cb<2> 12 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=2255 $Y=3566 $D=636
M1626 lb_mb<0> 13 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=2255 $Y=7966 $D=636
M1627 lb_mb<2> 14 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=2255 $Y=10026 $D=636
M1628 l_saeb_n 15 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=2255 $Y=35277 $D=636
M1629 lt_mb<2> 16 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=2255 $Y=39677 $D=636
M1630 lt_mb<0> 17 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=2255 $Y=41737 $D=636
M1631 lt_cb<2> 18 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=2255 $Y=46137 $D=636
M1632 lt_cb<0> 19 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=2255 $Y=48197 $D=636
M1633 vdd 15 l_saeb_n vdd hvtpfet l=6e-08 w=1.43e-06 $X=2515 $Y=35277 $D=636
M1634 vdd 34 lb_cb<1> vdd hvtpfet l=6e-08 w=1.43e-06 $X=2765 $Y=1506 $D=636
M1635 vdd 35 lb_cb<3> vdd hvtpfet l=6e-08 w=1.43e-06 $X=2765 $Y=3566 $D=636
M1636 vdd 36 lb_mb<1> vdd hvtpfet l=6e-08 w=1.43e-06 $X=2765 $Y=7966 $D=636
M1637 vdd 37 lb_mb<3> vdd hvtpfet l=6e-08 w=1.43e-06 $X=2765 $Y=10026 $D=636
M1638 vdd 39 lt_mb<3> vdd hvtpfet l=6e-08 w=1.43e-06 $X=2765 $Y=39677 $D=636
M1639 vdd 40 lt_mb<1> vdd hvtpfet l=6e-08 w=1.43e-06 $X=2765 $Y=41737 $D=636
M1640 vdd 41 lt_cb<3> vdd hvtpfet l=6e-08 w=1.43e-06 $X=2765 $Y=46137 $D=636
M1641 vdd 42 lt_cb<1> vdd hvtpfet l=6e-08 w=1.43e-06 $X=2765 $Y=48197 $D=636
M1642 l_saeb_n 15 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=2775 $Y=35277 $D=636
M1643 26 28 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=2821 $Y=15321 $D=636
M1644 1145 26 vdd vdd hvtpfet l=6e-08 w=2.74e-07 $X=2821 $Y=16069 $D=636
M1645 1146 4 vdd vdd hvtpfet l=6e-08 w=2.74e-07 $X=2821 $Y=20589 $D=636
M1646 4 29 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=2821 $Y=21405 $D=636
M1647 27 30 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=2821 $Y=22241 $D=636
M1648 1147 27 vdd vdd hvtpfet l=6e-08 w=2.74e-07 $X=2821 $Y=22989 $D=636
M1649 1148 3 vdd vdd hvtpfet l=6e-08 w=2.74e-07 $X=2821 $Y=27509 $D=636
M1650 3 31 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=2821 $Y=28325 $D=636
M1651 lb_cb<1> 34 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=3025 $Y=1506 $D=636
M1652 lb_cb<3> 35 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=3025 $Y=3566 $D=636
M1653 lb_mb<1> 36 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=3025 $Y=7966 $D=636
M1654 lb_mb<3> 37 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=3025 $Y=10026 $D=636
M1655 lt_mb<3> 39 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=3025 $Y=39677 $D=636
M1656 lt_mb<1> 40 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=3025 $Y=41737 $D=636
M1657 lt_cb<3> 41 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=3025 $Y=46137 $D=636
M1658 lt_cb<1> 42 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=3025 $Y=48197 $D=636
M1659 vdd 28 26 vdd hvtpfet l=6e-08 w=2.06e-07 $X=3081 $Y=15321 $D=636
M1660 28 43 1145 vdd hvtpfet l=6e-08 w=2.74e-07 $X=3081 $Y=16069 $D=636
M1661 29 43 1146 vdd hvtpfet l=6e-08 w=2.74e-07 $X=3081 $Y=20589 $D=636
M1662 vdd 29 4 vdd hvtpfet l=6e-08 w=2.06e-07 $X=3081 $Y=21405 $D=636
M1663 vdd 30 27 vdd hvtpfet l=6e-08 w=2.06e-07 $X=3081 $Y=22241 $D=636
M1664 30 43 1147 vdd hvtpfet l=6e-08 w=2.74e-07 $X=3081 $Y=22989 $D=636
M1665 31 43 1148 vdd hvtpfet l=6e-08 w=2.74e-07 $X=3081 $Y=27509 $D=636
M1666 vdd 31 3 vdd hvtpfet l=6e-08 w=2.06e-07 $X=3081 $Y=28325 $D=636
M1667 vdd 34 lb_cb<1> vdd hvtpfet l=6e-08 w=1.43e-06 $X=3285 $Y=1506 $D=636
M1668 vdd 35 lb_cb<3> vdd hvtpfet l=6e-08 w=1.43e-06 $X=3285 $Y=3566 $D=636
M1669 vdd 36 lb_mb<1> vdd hvtpfet l=6e-08 w=1.43e-06 $X=3285 $Y=7966 $D=636
M1670 vdd 37 lb_mb<3> vdd hvtpfet l=6e-08 w=1.43e-06 $X=3285 $Y=10026 $D=636
M1671 vdd 51 l_sa_preb_n vdd hvtpfet l=6e-08 w=1.43e-06 $X=3285 $Y=35277 $D=636
M1672 vdd 39 lt_mb<3> vdd hvtpfet l=6e-08 w=1.43e-06 $X=3285 $Y=39677 $D=636
M1673 vdd 40 lt_mb<1> vdd hvtpfet l=6e-08 w=1.43e-06 $X=3285 $Y=41737 $D=636
M1674 vdd 41 lt_cb<3> vdd hvtpfet l=6e-08 w=1.43e-06 $X=3285 $Y=46137 $D=636
M1675 vdd 42 lt_cb<1> vdd hvtpfet l=6e-08 w=1.43e-06 $X=3285 $Y=48197 $D=636
M1676 vdd ab<2> 44 vdd hvtpfet l=6e-08 w=4.11e-07 $X=3396 $Y=14280 $D=636
M1677 l_sa_preb_n 51 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=3545 $Y=35277 $D=636
M1678 vdd clkb 43 vdd hvtpfet l=6e-08 w=6e-07 $X=3546 $Y=33747 $D=636
M1679 1149 33 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=3591 $Y=15520 $D=636
M1680 1150 33 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=3591 $Y=20589 $D=636
M1681 1151 33 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=3591 $Y=22440 $D=636
M1682 1152 33 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=3591 $Y=27509 $D=636
M1683 52 stclkb vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=3705 $Y=29937 $D=636
M1684 vdd 47 34 vdd hvtpfet l=6e-08 w=1.2e-06 $X=3795 $Y=1736 $D=636
M1685 vdd 48 35 vdd hvtpfet l=6e-08 w=1.2e-06 $X=3795 $Y=3566 $D=636
M1686 vdd 27 36 vdd hvtpfet l=6e-08 w=1.2e-06 $X=3795 $Y=8196 $D=636
M1687 vdd 26 37 vdd hvtpfet l=6e-08 w=1.2e-06 $X=3795 $Y=10026 $D=636
M1688 vdd 26 39 vdd hvtpfet l=6e-08 w=1.2e-06 $X=3795 $Y=39907 $D=636
M1689 vdd 27 40 vdd hvtpfet l=6e-08 w=1.2e-06 $X=3795 $Y=41737 $D=636
M1690 vdd 49 41 vdd hvtpfet l=6e-08 w=1.2e-06 $X=3795 $Y=46367 $D=636
M1691 vdd 50 42 vdd hvtpfet l=6e-08 w=1.2e-06 $X=3795 $Y=48197 $D=636
M1692 vdd 51 l_sa_preb_n vdd hvtpfet l=6e-08 w=1.43e-06 $X=3805 $Y=35277 $D=636
M1693 43 clkb vdd vdd hvtpfet l=6e-08 w=6e-07 $X=3806 $Y=33747 $D=636
M1694 28 45 1149 vdd hvtpfet l=6e-08 w=4.11e-07 $X=3861 $Y=15932 $D=636
M1695 29 45 1150 vdd hvtpfet l=6e-08 w=4.11e-07 $X=3861 $Y=20589 $D=636
M1696 30 46 1151 vdd hvtpfet l=6e-08 w=4.11e-07 $X=3861 $Y=22852 $D=636
M1697 31 46 1152 vdd hvtpfet l=6e-08 w=4.11e-07 $X=3861 $Y=27509 $D=636
M1698 53 44 vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=3906 $Y=14280 $D=636
M1699 vdd clkb 43 vdd hvtpfet l=6e-08 w=6e-07 $X=4066 $Y=33747 $D=636
M1700 1153 53 28 vdd hvtpfet l=6e-08 w=4.11e-07 $X=4121 $Y=15932 $D=636
M1701 1154 44 29 vdd hvtpfet l=6e-08 w=4.11e-07 $X=4121 $Y=20589 $D=636
M1702 1155 53 30 vdd hvtpfet l=6e-08 w=4.11e-07 $X=4121 $Y=22852 $D=636
M1703 1156 44 31 vdd hvtpfet l=6e-08 w=4.11e-07 $X=4121 $Y=27509 $D=636
M1704 1157 52 59 vdd hvtpfet l=6e-08 w=8.23e-07 $X=4215 $Y=29525 $D=636
M1705 vdd 55 51 vdd hvtpfet l=6e-08 w=1.2e-06 $X=4315 $Y=35277 $D=636
M1706 43 clkb vdd vdd hvtpfet l=6e-08 w=6e-07 $X=4326 $Y=33747 $D=636
M1707 vdd 33 1153 vdd hvtpfet l=6e-08 w=8.23e-07 $X=4391 $Y=15520 $D=636
M1708 vdd 33 1154 vdd hvtpfet l=6e-08 w=8.23e-07 $X=4391 $Y=20589 $D=636
M1709 vdd 33 1155 vdd hvtpfet l=6e-08 w=8.23e-07 $X=4391 $Y=22440 $D=636
M1710 vdd 33 1156 vdd hvtpfet l=6e-08 w=8.23e-07 $X=4391 $Y=27509 $D=636
M1711 vdd ab<3> 46 vdd hvtpfet l=6e-08 w=4.11e-07 $X=4416 $Y=14280 $D=636
M1712 vdd 56 1157 vdd hvtpfet l=6e-08 w=8.23e-07 $X=4475 $Y=29525 $D=636
M1713 b_pxab<0> 60 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=4550 $Y=1941 $D=636
M1714 60 61 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=4550 $Y=5141 $D=636
M1715 61 62 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=4550 $Y=8691 $D=636
M1716 vdd 57 62 vdd hvtpfet l=6e-08 w=4.11e-07 $X=4550 $Y=10156 $D=636
M1717 vdd 57 63 vdd hvtpfet l=6e-08 w=4.11e-07 $X=4550 $Y=40566 $D=636
M1718 64 63 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=4550 $Y=41842 $D=636
M1719 65 64 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=4550 $Y=44992 $D=636
M1720 t_pxab<0> 65 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=4550 $Y=46622 $D=636
M1721 vdd 60 b_pxab<0> vdd hvtpfet l=6e-08 w=2.57e-06 $X=4810 $Y=1941 $D=636
M1722 vdd 61 60 vdd hvtpfet l=6e-08 w=1e-06 $X=4810 $Y=5141 $D=636
M1723 vdd 62 61 vdd hvtpfet l=6e-08 w=6e-07 $X=4810 $Y=8691 $D=636
M1724 62 24 vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=4810 $Y=10156 $D=636
M1725 63 25 vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=4810 $Y=40566 $D=636
M1726 vdd 63 64 vdd hvtpfet l=6e-08 w=6e-07 $X=4810 $Y=41842 $D=636
M1727 vdd 64 65 vdd hvtpfet l=6e-08 w=1e-06 $X=4810 $Y=44992 $D=636
M1728 vdd 65 t_pxab<0> vdd hvtpfet l=6e-08 w=2.57e-06 $X=4810 $Y=46622 $D=636
M1729 45 46 vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=4926 $Y=14280 $D=636
M1730 vdd 66 586 vdd hvtpfet l=1.4e-07 w=6.4e-07 $X=4939 $Y=36067 $D=636
M1731 1158 59 56 vdd hvtpfet l=6e-08 w=8.23e-07 $X=4985 $Y=29525 $D=636
M1732 vdd 58 587 vdd hvtpfet l=6e-08 w=6.4e-07 $X=5069 $Y=33468 $D=636
M1733 67 73 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=5141 $Y=15321 $D=636
M1734 1159 67 vdd vdd hvtpfet l=6e-08 w=2.74e-07 $X=5141 $Y=16069 $D=636
M1735 1160 68 vdd vdd hvtpfet l=6e-08 w=2.74e-07 $X=5141 $Y=20589 $D=636
M1736 68 74 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=5141 $Y=21405 $D=636
M1737 69 75 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=5141 $Y=22241 $D=636
M1738 1161 69 vdd vdd hvtpfet l=6e-08 w=2.74e-07 $X=5141 $Y=22989 $D=636
M1739 1162 57 vdd vdd hvtpfet l=6e-08 w=2.74e-07 $X=5141 $Y=27509 $D=636
M1740 57 76 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=5141 $Y=28325 $D=636
M1741 vdd 70 1158 vdd hvtpfet l=6e-08 w=8.23e-07 $X=5245 $Y=29525 $D=636
M1742 66 71 vdd vdd hvtpfet l=1.4e-07 w=6.4e-07 $X=5279 $Y=36067 $D=636
M1743 b_pxab<1> 78 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=5320 $Y=1941 $D=636
M1744 78 79 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=5320 $Y=5141 $D=636
M1745 79 80 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=5320 $Y=8691 $D=636
M1746 vdd 24 80 vdd hvtpfet l=6e-08 w=4.11e-07 $X=5320 $Y=10156 $D=636
M1747 vdd 25 81 vdd hvtpfet l=6e-08 w=4.11e-07 $X=5320 $Y=40566 $D=636
M1748 82 81 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=5320 $Y=41842 $D=636
M1749 83 82 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=5320 $Y=44992 $D=636
M1750 t_pxab<1> 83 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=5320 $Y=46622 $D=636
M1751 vdd 73 67 vdd hvtpfet l=6e-08 w=2.06e-07 $X=5401 $Y=15321 $D=636
M1752 73 43 1159 vdd hvtpfet l=6e-08 w=2.74e-07 $X=5401 $Y=16069 $D=636
M1753 74 43 1160 vdd hvtpfet l=6e-08 w=2.74e-07 $X=5401 $Y=20589 $D=636
M1754 vdd 74 68 vdd hvtpfet l=6e-08 w=2.06e-07 $X=5401 $Y=21405 $D=636
M1755 vdd 75 69 vdd hvtpfet l=6e-08 w=2.06e-07 $X=5401 $Y=22241 $D=636
M1756 75 43 1161 vdd hvtpfet l=6e-08 w=2.74e-07 $X=5401 $Y=22989 $D=636
M1757 76 43 1162 vdd hvtpfet l=6e-08 w=2.74e-07 $X=5401 $Y=27509 $D=636
M1758 vdd 76 57 vdd hvtpfet l=6e-08 w=2.06e-07 $X=5401 $Y=28325 $D=636
M1759 vdd 72 5 vdd hvtpfet l=6e-08 w=6.4e-07 $X=5579 $Y=33693 $D=636
M1760 vdd 78 b_pxab<1> vdd hvtpfet l=6e-08 w=2.57e-06 $X=5580 $Y=1941 $D=636
M1761 vdd 79 78 vdd hvtpfet l=6e-08 w=1e-06 $X=5580 $Y=5141 $D=636
M1762 vdd 80 79 vdd hvtpfet l=6e-08 w=6e-07 $X=5580 $Y=8691 $D=636
M1763 80 69 vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=5580 $Y=10156 $D=636
M1764 81 69 vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=5580 $Y=40566 $D=636
M1765 vdd 81 82 vdd hvtpfet l=6e-08 w=6e-07 $X=5580 $Y=41842 $D=636
M1766 vdd 82 83 vdd hvtpfet l=6e-08 w=1e-06 $X=5580 $Y=44992 $D=636
M1767 vdd 83 t_pxab<1> vdd hvtpfet l=6e-08 w=2.57e-06 $X=5580 $Y=46622 $D=636
M1768 vdd ab<5> 86 vdd hvtpfet l=6e-08 w=4.11e-07 $X=5716 $Y=14280 $D=636
M1769 5 85 vdd vdd hvtpfet l=6e-08 w=6.4e-07 $X=5839 $Y=33693 $D=636
M1770 1163 33 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=5911 $Y=15520 $D=636
M1771 1164 33 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=5911 $Y=20589 $D=636
M1772 1165 33 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=5911 $Y=22440 $D=636
M1773 1166 33 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=5911 $Y=27509 $D=636
M1774 70 clkb vdd vdd hvtpfet l=6e-08 w=1.2e-06 $X=6015 $Y=29148 $D=636
M1775 592 ddqb 71 vdd hvtpfet l=6e-08 w=6.4e-07 $X=6079 $Y=35802 $D=636
M1776 b_pxab<2> 90 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=6090 $Y=1941 $D=636
M1777 90 91 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=6090 $Y=5141 $D=636
M1778 91 92 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=6090 $Y=8691 $D=636
M1779 vdd 68 92 vdd hvtpfet l=6e-08 w=4.11e-07 $X=6090 $Y=10156 $D=636
M1780 vdd 68 93 vdd hvtpfet l=6e-08 w=4.11e-07 $X=6090 $Y=40566 $D=636
M1781 94 93 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=6090 $Y=41842 $D=636
M1782 95 94 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=6090 $Y=44992 $D=636
M1783 t_pxab<2> 95 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=6090 $Y=46622 $D=636
M1784 73 87 1163 vdd hvtpfet l=6e-08 w=4.11e-07 $X=6181 $Y=15932 $D=636
M1785 74 87 1164 vdd hvtpfet l=6e-08 w=4.11e-07 $X=6181 $Y=20589 $D=636
M1786 75 88 1165 vdd hvtpfet l=6e-08 w=4.11e-07 $X=6181 $Y=22852 $D=636
M1787 76 88 1166 vdd hvtpfet l=6e-08 w=4.11e-07 $X=6181 $Y=27509 $D=636
M1788 97 86 vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=6226 $Y=14280 $D=636
M1789 vdd ddqb_n 592 vdd hvtpfet l=6e-08 w=6.4e-07 $X=6339 $Y=35802 $D=636
M1790 vdd 90 b_pxab<2> vdd hvtpfet l=6e-08 w=2.57e-06 $X=6350 $Y=1941 $D=636
M1791 vdd 91 90 vdd hvtpfet l=6e-08 w=1e-06 $X=6350 $Y=5141 $D=636
M1792 vdd 92 91 vdd hvtpfet l=6e-08 w=6e-07 $X=6350 $Y=8691 $D=636
M1793 92 24 vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=6350 $Y=10156 $D=636
M1794 93 25 vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=6350 $Y=40566 $D=636
M1795 vdd 93 94 vdd hvtpfet l=6e-08 w=6e-07 $X=6350 $Y=41842 $D=636
M1796 vdd 94 95 vdd hvtpfet l=6e-08 w=1e-06 $X=6350 $Y=44992 $D=636
M1797 vdd 95 t_pxab<2> vdd hvtpfet l=6e-08 w=2.57e-06 $X=6350 $Y=46622 $D=636
M1798 1167 97 73 vdd hvtpfet l=6e-08 w=4.11e-07 $X=6441 $Y=15932 $D=636
M1799 1168 86 74 vdd hvtpfet l=6e-08 w=4.11e-07 $X=6441 $Y=20589 $D=636
M1800 1169 97 75 vdd hvtpfet l=6e-08 w=4.11e-07 $X=6441 $Y=22852 $D=636
M1801 1170 86 76 vdd hvtpfet l=6e-08 w=4.11e-07 $X=6441 $Y=27509 $D=636
M1802 85 89 vdd vdd hvtpfet l=6e-08 w=6.4e-07 $X=6524 $Y=33693 $D=636
M1803 142 clkb vdd vdd hvtpfet l=6e-08 w=8e-07 $X=6525 $Y=29548 $D=636
M1804 vdd 33 1167 vdd hvtpfet l=6e-08 w=8.23e-07 $X=6711 $Y=15520 $D=636
M1805 vdd 33 1168 vdd hvtpfet l=6e-08 w=8.23e-07 $X=6711 $Y=20589 $D=636
M1806 vdd 33 1169 vdd hvtpfet l=6e-08 w=8.23e-07 $X=6711 $Y=22440 $D=636
M1807 vdd 33 1170 vdd hvtpfet l=6e-08 w=8.23e-07 $X=6711 $Y=27509 $D=636
M1808 vdd ab<6> 88 vdd hvtpfet l=6e-08 w=4.11e-07 $X=6736 $Y=14280 $D=636
M1809 vdd clkb 142 vdd hvtpfet l=6e-08 w=8e-07 $X=6785 $Y=29548 $D=636
M1810 b_pxab<3> 99 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=6860 $Y=1941 $D=636
M1811 99 100 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=6860 $Y=5141 $D=636
M1812 100 101 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=6860 $Y=8691 $D=636
M1813 vdd 24 101 vdd hvtpfet l=6e-08 w=4.11e-07 $X=6860 $Y=10156 $D=636
M1814 vdd 25 102 vdd hvtpfet l=6e-08 w=4.11e-07 $X=6860 $Y=40566 $D=636
M1815 103 102 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=6860 $Y=41842 $D=636
M1816 104 103 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=6860 $Y=44992 $D=636
M1817 t_pxab<3> 104 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=6860 $Y=46622 $D=636
M1818 109 85 vdd vdd hvtpfet l=6e-08 w=6.4e-07 $X=7034 $Y=33468 $D=636
M1819 89 71 vdd vdd hvtpfet l=6e-08 w=6.4e-07 $X=7069 $Y=35802 $D=636
M1820 vdd 99 b_pxab<3> vdd hvtpfet l=6e-08 w=2.57e-06 $X=7120 $Y=1941 $D=636
M1821 vdd 100 99 vdd hvtpfet l=6e-08 w=1e-06 $X=7120 $Y=5141 $D=636
M1822 vdd 101 100 vdd hvtpfet l=6e-08 w=6e-07 $X=7120 $Y=8691 $D=636
M1823 101 67 vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=7120 $Y=10156 $D=636
M1824 102 67 vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=7120 $Y=40566 $D=636
M1825 vdd 102 103 vdd hvtpfet l=6e-08 w=6e-07 $X=7120 $Y=41842 $D=636
M1826 vdd 103 104 vdd hvtpfet l=6e-08 w=1e-06 $X=7120 $Y=44992 $D=636
M1827 vdd 104 t_pxab<3> vdd hvtpfet l=6e-08 w=2.57e-06 $X=7120 $Y=46622 $D=636
M1828 87 88 vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=7246 $Y=14280 $D=636
M1829 142 59 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=7295 $Y=29548 $D=636
M1830 105 111 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=7461 $Y=15321 $D=636
M1831 1171 105 vdd vdd hvtpfet l=6e-08 w=2.74e-07 $X=7461 $Y=16069 $D=636
M1832 1172 106 vdd vdd hvtpfet l=6e-08 w=2.74e-07 $X=7461 $Y=20589 $D=636
M1833 106 112 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=7461 $Y=21405 $D=636
M1834 107 113 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=7461 $Y=22241 $D=636
M1835 1173 107 vdd vdd hvtpfet l=6e-08 w=2.74e-07 $X=7461 $Y=22989 $D=636
M1836 1174 108 vdd vdd hvtpfet l=6e-08 w=2.74e-07 $X=7461 $Y=27509 $D=636
M1837 108 114 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=7461 $Y=28325 $D=636
M1838 vdd 59 142 vdd hvtpfet l=6e-08 w=8e-07 $X=7555 $Y=29548 $D=636
M1839 vdd 110 89 vdd hvtpfet l=1.2e-07 w=3e-07 $X=7579 $Y=36382 $D=636
M1840 b_pxbb_n<0> 115 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=7630 $Y=1941 $D=636
M1841 115 116 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=7630 $Y=5141 $D=636
M1842 116 107 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=7630 $Y=8691 $D=636
M1843 117 107 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=7630 $Y=41842 $D=636
M1844 118 117 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=7630 $Y=44992 $D=636
M1845 t_pxbb_n<0> 118 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=7630 $Y=46622 $D=636
M1846 vdd 109 119 vdd hvtpfet l=6e-08 w=5e-07 $X=7634 $Y=33503 $D=636
M1847 vdd 111 105 vdd hvtpfet l=6e-08 w=2.06e-07 $X=7721 $Y=15321 $D=636
M1848 111 43 1171 vdd hvtpfet l=6e-08 w=2.74e-07 $X=7721 $Y=16069 $D=636
M1849 112 43 1172 vdd hvtpfet l=6e-08 w=2.74e-07 $X=7721 $Y=20589 $D=636
M1850 vdd 112 106 vdd hvtpfet l=6e-08 w=2.06e-07 $X=7721 $Y=21405 $D=636
M1851 vdd 113 107 vdd hvtpfet l=6e-08 w=2.06e-07 $X=7721 $Y=22241 $D=636
M1852 113 43 1173 vdd hvtpfet l=6e-08 w=2.74e-07 $X=7721 $Y=22989 $D=636
M1853 114 43 1174 vdd hvtpfet l=6e-08 w=2.74e-07 $X=7721 $Y=27509 $D=636
M1854 vdd 114 108 vdd hvtpfet l=6e-08 w=2.06e-07 $X=7721 $Y=28325 $D=636
M1855 vdd 115 b_pxbb_n<0> vdd hvtpfet l=6e-08 w=2.57e-06 $X=7890 $Y=1941 $D=636
M1856 vdd 116 115 vdd hvtpfet l=6e-08 w=1e-06 $X=7890 $Y=5141 $D=636
M1857 vdd 107 116 vdd hvtpfet l=6e-08 w=6e-07 $X=7890 $Y=8691 $D=636
M1858 vdd 107 117 vdd hvtpfet l=6e-08 w=6e-07 $X=7890 $Y=41842 $D=636
M1859 vdd 117 118 vdd hvtpfet l=6e-08 w=1e-06 $X=7890 $Y=44992 $D=636
M1860 vdd 118 t_pxbb_n<0> vdd hvtpfet l=6e-08 w=2.57e-06 $X=7890 $Y=46622 $D=636
M1861 120 119 vdd vdd hvtpfet l=2.5e-07 w=5e-07 $X=7894 $Y=33503 $D=636
M1862 110 89 vdd vdd hvtpfet l=6e-08 w=3e-07 $X=8149 $Y=36377 $D=636
M1863 1175 33 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=8231 $Y=15520 $D=636
M1864 1176 33 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=8231 $Y=20589 $D=636
M1865 1177 33 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=8231 $Y=22440 $D=636
M1866 1178 33 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=8231 $Y=27509 $D=636
M1867 b_pxbb_n<1> 125 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=8400 $Y=1941 $D=636
M1868 125 126 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=8400 $Y=5141 $D=636
M1869 126 108 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=8400 $Y=8691 $D=636
M1870 127 108 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=8400 $Y=41842 $D=636
M1871 128 127 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=8400 $Y=44992 $D=636
M1872 t_pxbb_n<1> 128 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=8400 $Y=46622 $D=636
M1873 vdd 122 121 vdd hvtpfet l=6e-08 w=4.11e-07 $X=8466 $Y=14280 $D=636
M1874 111 121 1175 vdd hvtpfet l=6e-08 w=4.11e-07 $X=8501 $Y=15932 $D=636
M1875 112 121 1176 vdd hvtpfet l=6e-08 w=4.11e-07 $X=8501 $Y=20589 $D=636
M1876 113 122 1177 vdd hvtpfet l=6e-08 w=4.11e-07 $X=8501 $Y=22852 $D=636
M1877 114 122 1178 vdd hvtpfet l=6e-08 w=4.11e-07 $X=8501 $Y=27509 $D=636
M1878 131 123 vdd vdd hvtpfet l=6e-08 w=2e-07 $X=8594 $Y=10756 $D=636
M1879 vdd 120 55 vdd hvtpfet l=6e-08 w=6.4e-07 $X=8619 $Y=33468 $D=636
M1880 602 124 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=8659 $Y=29348 $D=636
M1881 603 124 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=8659 $Y=35707 $D=636
M1882 vdd 125 b_pxbb_n<1> vdd hvtpfet l=6e-08 w=2.57e-06 $X=8660 $Y=1941 $D=636
M1883 vdd 126 125 vdd hvtpfet l=6e-08 w=1e-06 $X=8660 $Y=5141 $D=636
M1884 vdd 108 126 vdd hvtpfet l=6e-08 w=6e-07 $X=8660 $Y=8691 $D=636
M1885 vdd 108 127 vdd hvtpfet l=6e-08 w=6e-07 $X=8660 $Y=41842 $D=636
M1886 vdd 127 128 vdd hvtpfet l=6e-08 w=1e-06 $X=8660 $Y=44992 $D=636
M1887 vdd 128 t_pxbb_n<1> vdd hvtpfet l=6e-08 w=2.57e-06 $X=8660 $Y=46622 $D=636
M1888 1179 129 111 vdd hvtpfet l=6e-08 w=4.11e-07 $X=8761 $Y=15932 $D=636
M1889 1180 129 112 vdd hvtpfet l=6e-08 w=4.11e-07 $X=8761 $Y=20589 $D=636
M1890 1181 129 113 vdd hvtpfet l=6e-08 w=4.11e-07 $X=8761 $Y=22852 $D=636
M1891 1182 129 114 vdd hvtpfet l=6e-08 w=4.11e-07 $X=8761 $Y=27509 $D=636
M1892 55 vdd vdd vdd hvtpfet l=6e-08 w=6.4e-07 $X=8879 $Y=33468 $D=636
M1893 vdd 124 602 vdd hvtpfet l=6e-08 w=1e-06 $X=8919 $Y=29348 $D=636
M1894 vdd 124 603 vdd hvtpfet l=6e-08 w=1e-06 $X=8919 $Y=35707 $D=636
M1895 122 ab<9> vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=8976 $Y=14280 $D=636
M1896 vdd 33 1179 vdd hvtpfet l=6e-08 w=8.23e-07 $X=9031 $Y=15520 $D=636
M1897 vdd 33 1180 vdd hvtpfet l=6e-08 w=8.23e-07 $X=9031 $Y=20589 $D=636
M1898 vdd 33 1181 vdd hvtpfet l=6e-08 w=8.23e-07 $X=9031 $Y=22440 $D=636
M1899 vdd 33 1182 vdd hvtpfet l=6e-08 w=8.23e-07 $X=9031 $Y=27509 $D=636
M1900 b_pxbb_n<2> 135 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=9170 $Y=1941 $D=636
M1901 135 136 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=9170 $Y=5141 $D=636
M1902 136 137 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=9170 $Y=8691 $D=636
M1903 138 137 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=9170 $Y=41842 $D=636
M1904 139 138 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=9170 $Y=44992 $D=636
M1905 t_pxbb_n<2> 139 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=9170 $Y=46622 $D=636
M1906 dwlb<0> 142 602 vdd hvtpfet l=6e-08 w=1e-06 $X=9429 $Y=29348 $D=636
M1907 25 143 603 vdd hvtpfet l=6e-08 w=1e-06 $X=9429 $Y=35707 $D=636
M1908 vdd 135 b_pxbb_n<2> vdd hvtpfet l=6e-08 w=2.57e-06 $X=9430 $Y=1941 $D=636
M1909 vdd 136 135 vdd hvtpfet l=6e-08 w=1e-06 $X=9430 $Y=5141 $D=636
M1910 vdd 137 136 vdd hvtpfet l=6e-08 w=6e-07 $X=9430 $Y=8691 $D=636
M1911 vdd 137 138 vdd hvtpfet l=6e-08 w=6e-07 $X=9430 $Y=41842 $D=636
M1912 vdd 138 139 vdd hvtpfet l=6e-08 w=1e-06 $X=9430 $Y=44992 $D=636
M1913 vdd 139 t_pxbb_n<2> vdd hvtpfet l=6e-08 w=2.57e-06 $X=9430 $Y=46622 $D=636
M1914 1183 132 111 vdd hvtpfet l=6e-08 w=4.11e-07 $X=9541 $Y=15932 $D=636
M1915 1184 133 112 vdd hvtpfet l=6e-08 w=4.11e-07 $X=9541 $Y=20589 $D=636
M1916 1185 132 113 vdd hvtpfet l=6e-08 w=4.11e-07 $X=9541 $Y=22852 $D=636
M1917 1186 133 114 vdd hvtpfet l=6e-08 w=4.11e-07 $X=9541 $Y=27509 $D=636
M1918 vdd 140 1 vdd hvtpfet l=6e-08 w=4e-07 $X=9586 $Y=10167 $D=636
M1919 vdd 141 7 vdd hvtpfet l=6e-08 w=4e-07 $X=9586 $Y=40566 $D=636
M1920 602 142 dwlb<0> vdd hvtpfet l=6e-08 w=1e-06 $X=9689 $Y=29348 $D=636
M1921 603 143 25 vdd hvtpfet l=6e-08 w=1e-06 $X=9689 $Y=35707 $D=636
M1922 vdd 33 1183 vdd hvtpfet l=6e-08 w=8.23e-07 $X=9811 $Y=15520 $D=636
M1923 vdd 33 1184 vdd hvtpfet l=6e-08 w=8.23e-07 $X=9811 $Y=20589 $D=636
M1924 vdd 33 1185 vdd hvtpfet l=6e-08 w=8.23e-07 $X=9811 $Y=22440 $D=636
M1925 vdd 33 1186 vdd hvtpfet l=6e-08 w=8.23e-07 $X=9811 $Y=27509 $D=636
M1926 b_pxbb_n<3> 146 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=9940 $Y=1941 $D=636
M1927 146 147 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=9940 $Y=5141 $D=636
M1928 147 148 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=9940 $Y=8691 $D=636
M1929 149 148 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=9940 $Y=41842 $D=636
M1930 150 149 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=9940 $Y=44992 $D=636
M1931 t_pxbb_n<3> 150 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=9940 $Y=46622 $D=636
M1932 vdd ab<8> 129 vdd hvtpfet l=6e-08 w=4.11e-07 $X=9986 $Y=14280 $D=636
M1933 1187 33 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=10071 $Y=15520 $D=636
M1934 1188 33 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=10071 $Y=20589 $D=636
M1935 1189 33 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=10071 $Y=22440 $D=636
M1936 1190 33 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=10071 $Y=27509 $D=636
M1937 vdd 145 140 vdd hvtpfet l=6e-08 w=4.11e-07 $X=10096 $Y=10156 $D=636
M1938 vdd 145 141 vdd hvtpfet l=6e-08 w=4.11e-07 $X=10096 $Y=40566 $D=636
M1939 dwlb<1> 142 608 vdd hvtpfet l=6e-08 w=1e-06 $X=10199 $Y=29348 $D=636
M1940 24 143 609 vdd hvtpfet l=6e-08 w=1e-06 $X=10199 $Y=35707 $D=636
M1941 vdd 146 b_pxbb_n<3> vdd hvtpfet l=6e-08 w=2.57e-06 $X=10200 $Y=1941 $D=636
M1942 vdd 147 146 vdd hvtpfet l=6e-08 w=1e-06 $X=10200 $Y=5141 $D=636
M1943 vdd 148 147 vdd hvtpfet l=6e-08 w=6e-07 $X=10200 $Y=8691 $D=636
M1944 vdd 148 149 vdd hvtpfet l=6e-08 w=6e-07 $X=10200 $Y=41842 $D=636
M1945 vdd 149 150 vdd hvtpfet l=6e-08 w=1e-06 $X=10200 $Y=44992 $D=636
M1946 vdd 150 t_pxbb_n<3> vdd hvtpfet l=6e-08 w=2.57e-06 $X=10200 $Y=46622 $D=636
M1947 160 129 vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=10246 $Y=14280 $D=636
M1948 168 132 1187 vdd hvtpfet l=6e-08 w=4.11e-07 $X=10341 $Y=15932 $D=636
M1949 169 133 1188 vdd hvtpfet l=6e-08 w=4.11e-07 $X=10341 $Y=20589 $D=636
M1950 170 132 1189 vdd hvtpfet l=6e-08 w=4.11e-07 $X=10341 $Y=22852 $D=636
M1951 171 133 1190 vdd hvtpfet l=6e-08 w=4.11e-07 $X=10341 $Y=27509 $D=636
M1952 140 dwlb<1> vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=10356 $Y=10156 $D=636
M1953 141 dwlb<0> vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=10356 $Y=40566 $D=636
M1954 vdd 153 124 vdd hvtpfet l=6e-08 w=8e-07 $X=10406 $Y=33493 $D=636
M1955 608 142 dwlb<1> vdd hvtpfet l=6e-08 w=1e-06 $X=10459 $Y=29348 $D=636
M1956 609 143 24 vdd hvtpfet l=6e-08 w=1e-06 $X=10459 $Y=35707 $D=636
M1957 b_pxbb_n<4> 156 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=10710 $Y=1941 $D=636
M1958 156 157 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=10710 $Y=5141 $D=636
M1959 157 105 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=10710 $Y=8691 $D=636
M1960 158 105 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=10710 $Y=41842 $D=636
M1961 159 158 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=10710 $Y=44992 $D=636
M1962 t_pxbb_n<4> 159 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=10710 $Y=46622 $D=636
M1963 vdd 132 133 vdd hvtpfet l=6e-08 w=4.11e-07 $X=10846 $Y=14280 $D=636
M1964 1191 33 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=10851 $Y=15520 $D=636
M1965 1192 33 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=10851 $Y=20589 $D=636
M1966 1193 33 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=10851 $Y=22440 $D=636
M1967 1194 33 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=10851 $Y=27509 $D=636
M1968 vdd dwlb<1> 162 vdd hvtpfet l=6e-08 w=4.11e-07 $X=10866 $Y=10156 $D=636
M1969 vdd dwlb<0> 163 vdd hvtpfet l=6e-08 w=4.11e-07 $X=10866 $Y=40566 $D=636
M1970 608 153 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=10969 $Y=29348 $D=636
M1971 609 153 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=10969 $Y=35707 $D=636
M1972 vdd 156 b_pxbb_n<4> vdd hvtpfet l=6e-08 w=2.57e-06 $X=10970 $Y=1941 $D=636
M1973 vdd 157 156 vdd hvtpfet l=6e-08 w=1e-06 $X=10970 $Y=5141 $D=636
M1974 vdd 105 157 vdd hvtpfet l=6e-08 w=6e-07 $X=10970 $Y=8691 $D=636
M1975 vdd 105 158 vdd hvtpfet l=6e-08 w=6e-07 $X=10970 $Y=41842 $D=636
M1976 vdd 158 159 vdd hvtpfet l=6e-08 w=1e-06 $X=10970 $Y=44992 $D=636
M1977 vdd 159 t_pxbb_n<4> vdd hvtpfet l=6e-08 w=2.57e-06 $X=10970 $Y=46622 $D=636
M1978 132 ab<7> vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=11106 $Y=14280 $D=636
M1979 153 154 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=11106 $Y=33493 $D=636
M1980 168 160 1191 vdd hvtpfet l=6e-08 w=4.11e-07 $X=11121 $Y=15932 $D=636
M1981 169 160 1192 vdd hvtpfet l=6e-08 w=4.11e-07 $X=11121 $Y=20589 $D=636
M1982 170 160 1193 vdd hvtpfet l=6e-08 w=4.11e-07 $X=11121 $Y=22852 $D=636
M1983 171 160 1194 vdd hvtpfet l=6e-08 w=4.11e-07 $X=11121 $Y=27509 $D=636
M1984 162 155 vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=11126 $Y=10156 $D=636
M1985 163 155 vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=11126 $Y=40566 $D=636
M1986 vdd 153 608 vdd hvtpfet l=6e-08 w=1e-06 $X=11229 $Y=29348 $D=636
M1987 vdd 153 609 vdd hvtpfet l=6e-08 w=1e-06 $X=11229 $Y=35707 $D=636
M1988 1195 121 168 vdd hvtpfet l=6e-08 w=4.11e-07 $X=11381 $Y=15932 $D=636
M1989 1196 121 169 vdd hvtpfet l=6e-08 w=4.11e-07 $X=11381 $Y=20589 $D=636
M1990 1197 122 170 vdd hvtpfet l=6e-08 w=4.11e-07 $X=11381 $Y=22852 $D=636
M1991 1198 122 171 vdd hvtpfet l=6e-08 w=4.11e-07 $X=11381 $Y=27509 $D=636
M1992 b_pxbb_n<5> 164 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=11480 $Y=1941 $D=636
M1993 164 165 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=11480 $Y=5141 $D=636
M1994 165 106 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=11480 $Y=8691 $D=636
M1995 166 106 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=11480 $Y=41842 $D=636
M1996 167 166 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=11480 $Y=44992 $D=636
M1997 t_pxbb_n<5> 167 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=11480 $Y=46622 $D=636
M1998 47 162 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=11636 $Y=10167 $D=636
M1999 50 163 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=11636 $Y=40566 $D=636
M2000 vdd 33 1195 vdd hvtpfet l=6e-08 w=8.23e-07 $X=11651 $Y=15520 $D=636
M2001 vdd 33 1196 vdd hvtpfet l=6e-08 w=8.23e-07 $X=11651 $Y=20589 $D=636
M2002 vdd 33 1197 vdd hvtpfet l=6e-08 w=8.23e-07 $X=11651 $Y=22440 $D=636
M2003 vdd 33 1198 vdd hvtpfet l=6e-08 w=8.23e-07 $X=11651 $Y=27509 $D=636
M2004 172 142 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=11739 $Y=29948 $D=636
M2005 vdd 164 b_pxbb_n<5> vdd hvtpfet l=6e-08 w=2.57e-06 $X=11740 $Y=1941 $D=636
M2006 vdd 165 164 vdd hvtpfet l=6e-08 w=1e-06 $X=11740 $Y=5141 $D=636
M2007 vdd 106 165 vdd hvtpfet l=6e-08 w=6e-07 $X=11740 $Y=8691 $D=636
M2008 vdd 106 166 vdd hvtpfet l=6e-08 w=6e-07 $X=11740 $Y=41842 $D=636
M2009 vdd 166 167 vdd hvtpfet l=6e-08 w=1e-06 $X=11740 $Y=44992 $D=636
M2010 vdd 167 t_pxbb_n<5> vdd hvtpfet l=6e-08 w=2.57e-06 $X=11740 $Y=46622 $D=636
M2011 vdd tm<0> dbl_pd_n<0> vdd hvtpfet l=6e-08 w=4.28e-07 $X=11746 $Y=14263 $D=636
M2012 616 172 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=11933 $Y=35707 $D=636
M2013 dbl_pd_n<0> tm<0> vdd vdd hvtpfet l=6e-08 w=4.28e-07 $X=12006 $Y=14263 $D=636
M2014 179 173 vdd vdd hvtpfet l=6e-08 w=3e-07 $X=12086 $Y=33468 $D=636
M2015 vdd 174 2 vdd hvtpfet l=6e-08 w=4e-07 $X=12146 $Y=10167 $D=636
M2016 vdd 175 6 vdd hvtpfet l=6e-08 w=4e-07 $X=12146 $Y=40566 $D=636
M2017 177 168 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=12161 $Y=15321 $D=636
M2018 1199 43 168 vdd hvtpfet l=6e-08 w=2.74e-07 $X=12161 $Y=16069 $D=636
M2019 1200 43 169 vdd hvtpfet l=6e-08 w=2.74e-07 $X=12161 $Y=20589 $D=636
M2020 178 169 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=12161 $Y=21405 $D=636
M2021 137 170 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=12161 $Y=22241 $D=636
M2022 1201 43 170 vdd hvtpfet l=6e-08 w=2.74e-07 $X=12161 $Y=22989 $D=636
M2023 1202 43 171 vdd hvtpfet l=6e-08 w=2.74e-07 $X=12161 $Y=27509 $D=636
M2024 148 171 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=12161 $Y=28325 $D=636
M2025 vdd 172 616 vdd hvtpfet l=6e-08 w=1e-06 $X=12193 $Y=35707 $D=636
M2026 b_pxbb_n<6> 180 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=12250 $Y=1941 $D=636
M2027 180 181 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=12250 $Y=5141 $D=636
M2028 181 177 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=12250 $Y=8691 $D=636
M2029 182 177 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=12250 $Y=41842 $D=636
M2030 183 182 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=12250 $Y=44992 $D=636
M2031 t_pxbb_n<6> 183 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=12250 $Y=46622 $D=636
M2032 vdd tm<0> dbl_pd_n<0> vdd hvtpfet l=6e-08 w=4.28e-07 $X=12266 $Y=14263 $D=636
M2033 vdd 142 184 vdd hvtpfet l=6e-08 w=5e-07 $X=12339 $Y=29813 $D=636
M2034 vdd 168 177 vdd hvtpfet l=6e-08 w=2.06e-07 $X=12421 $Y=15321 $D=636
M2035 vdd 177 1199 vdd hvtpfet l=6e-08 w=2.74e-07 $X=12421 $Y=16069 $D=636
M2036 vdd 178 1200 vdd hvtpfet l=6e-08 w=2.74e-07 $X=12421 $Y=20589 $D=636
M2037 vdd 169 178 vdd hvtpfet l=6e-08 w=2.06e-07 $X=12421 $Y=21405 $D=636
M2038 vdd 170 137 vdd hvtpfet l=6e-08 w=2.06e-07 $X=12421 $Y=22241 $D=636
M2039 vdd 137 1201 vdd hvtpfet l=6e-08 w=2.74e-07 $X=12421 $Y=22989 $D=636
M2040 vdd 148 1202 vdd hvtpfet l=6e-08 w=2.74e-07 $X=12421 $Y=27509 $D=636
M2041 vdd 171 148 vdd hvtpfet l=6e-08 w=2.06e-07 $X=12421 $Y=28325 $D=636
M2042 616 172 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=12453 $Y=35707 $D=636
M2043 vdd 180 b_pxbb_n<6> vdd hvtpfet l=6e-08 w=2.57e-06 $X=12510 $Y=1941 $D=636
M2044 vdd 181 180 vdd hvtpfet l=6e-08 w=1e-06 $X=12510 $Y=5141 $D=636
M2045 vdd 177 181 vdd hvtpfet l=6e-08 w=6e-07 $X=12510 $Y=8691 $D=636
M2046 vdd 177 182 vdd hvtpfet l=6e-08 w=6e-07 $X=12510 $Y=41842 $D=636
M2047 vdd 182 183 vdd hvtpfet l=6e-08 w=1e-06 $X=12510 $Y=44992 $D=636
M2048 vdd 183 t_pxbb_n<6> vdd hvtpfet l=6e-08 w=2.57e-06 $X=12510 $Y=46622 $D=636
M2049 615 179 186 vdd hvtpfet l=6e-08 w=6e-07 $X=12596 $Y=33468 $D=636
M2050 191 184 vdd vdd hvtpfet l=2.5e-07 w=5e-07 $X=12599 $Y=29813 $D=636
M2051 vdd 185 174 vdd hvtpfet l=6e-08 w=4.11e-07 $X=12656 $Y=10156 $D=636
M2052 vdd 185 175 vdd hvtpfet l=6e-08 w=4.11e-07 $X=12656 $Y=40566 $D=636
M2053 620 186 616 vdd hvtpfet l=6e-08 w=1e-06 $X=12713 $Y=35707 $D=636
M2054 vdd 131 dbl_pd_n<2> vdd hvtpfet l=6e-08 w=4.28e-07 $X=12776 $Y=14263 $D=636
M2055 vdd 191 615 vdd hvtpfet l=6e-08 w=6e-07 $X=12856 $Y=33468 $D=636
M2056 174 dwlb<1> vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=12916 $Y=10156 $D=636
M2057 175 dwlb<0> vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=12916 $Y=40566 $D=636
M2058 187 192 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=12931 $Y=15321 $D=636
M2059 1203 187 vdd vdd hvtpfet l=6e-08 w=2.74e-07 $X=12931 $Y=16069 $D=636
M2060 1204 188 vdd vdd hvtpfet l=6e-08 w=2.74e-07 $X=12931 $Y=20589 $D=636
M2061 188 193 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=12931 $Y=21405 $D=636
M2062 189 194 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=12931 $Y=22241 $D=636
M2063 1205 189 vdd vdd hvtpfet l=6e-08 w=2.74e-07 $X=12931 $Y=22989 $D=636
M2064 1206 190 vdd vdd hvtpfet l=6e-08 w=2.74e-07 $X=12931 $Y=27509 $D=636
M2065 190 195 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=12931 $Y=28325 $D=636
M2066 616 186 620 vdd hvtpfet l=6e-08 w=1e-06 $X=12973 $Y=35707 $D=636
M2067 b_pxbb_n<7> 196 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=13020 $Y=1941 $D=636
M2068 196 197 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=13020 $Y=5141 $D=636
M2069 197 178 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=13020 $Y=8691 $D=636
M2070 198 178 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=13020 $Y=41842 $D=636
M2071 199 198 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=13020 $Y=44992 $D=636
M2072 t_pxbb_n<7> 199 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=13020 $Y=46622 $D=636
M2073 dbl_pd_n<2> 131 vdd vdd hvtpfet l=6e-08 w=4.28e-07 $X=13036 $Y=14263 $D=636
M2074 vdd 192 187 vdd hvtpfet l=6e-08 w=2.06e-07 $X=13191 $Y=15321 $D=636
M2075 192 43 1203 vdd hvtpfet l=6e-08 w=2.74e-07 $X=13191 $Y=16069 $D=636
M2076 193 43 1204 vdd hvtpfet l=6e-08 w=2.74e-07 $X=13191 $Y=20589 $D=636
M2077 vdd 193 188 vdd hvtpfet l=6e-08 w=2.06e-07 $X=13191 $Y=21405 $D=636
M2078 vdd 194 189 vdd hvtpfet l=6e-08 w=2.06e-07 $X=13191 $Y=22241 $D=636
M2079 194 43 1205 vdd hvtpfet l=6e-08 w=2.74e-07 $X=13191 $Y=22989 $D=636
M2080 195 43 1206 vdd hvtpfet l=6e-08 w=2.74e-07 $X=13191 $Y=27509 $D=636
M2081 vdd 195 190 vdd hvtpfet l=6e-08 w=2.06e-07 $X=13191 $Y=28325 $D=636
M2082 620 186 616 vdd hvtpfet l=6e-08 w=1e-06 $X=13233 $Y=35707 $D=636
M2083 vdd 196 b_pxbb_n<7> vdd hvtpfet l=6e-08 w=2.57e-06 $X=13280 $Y=1941 $D=636
M2084 vdd 197 196 vdd hvtpfet l=6e-08 w=1e-06 $X=13280 $Y=5141 $D=636
M2085 vdd 178 197 vdd hvtpfet l=6e-08 w=6e-07 $X=13280 $Y=8691 $D=636
M2086 vdd 178 198 vdd hvtpfet l=6e-08 w=6e-07 $X=13280 $Y=41842 $D=636
M2087 vdd 198 199 vdd hvtpfet l=6e-08 w=1e-06 $X=13280 $Y=44992 $D=636
M2088 vdd 199 t_pxbb_n<7> vdd hvtpfet l=6e-08 w=2.57e-06 $X=13280 $Y=46622 $D=636
M2089 vdd 131 dbl_pd_n<2> vdd hvtpfet l=6e-08 w=4.28e-07 $X=13296 $Y=14263 $D=636
M2090 vdd tm<7> 203 vdd hvtpfet l=6e-08 w=3e-07 $X=13432 $Y=33468 $D=636
M2091 vdd 191 202 vdd hvtpfet l=6e-08 w=5e-07 $X=13459 $Y=29813 $D=636
M2092 143 200 620 vdd hvtpfet l=6e-08 w=1e-06 $X=13493 $Y=35707 $D=636
M2093 1207 33 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=13701 $Y=15520 $D=636
M2094 1208 33 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=13701 $Y=20589 $D=636
M2095 1209 33 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=13701 $Y=22440 $D=636
M2096 1210 33 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=13701 $Y=27509 $D=636
M2097 211 202 vdd vdd hvtpfet l=2.5e-07 w=5e-07 $X=13719 $Y=29813 $D=636
M2098 620 200 143 vdd hvtpfet l=6e-08 w=1e-06 $X=13753 $Y=35707 $D=636
M2099 b_pxcb_n<0> 206 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=13790 $Y=1941 $D=636
M2100 206 207 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=13790 $Y=5141 $D=636
M2101 207 189 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=13790 $Y=8691 $D=636
M2102 208 189 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=13790 $Y=41842 $D=636
M2103 209 208 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=13790 $Y=44992 $D=636
M2104 t_pxcb_n<0> 209 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=13790 $Y=46622 $D=636
M2105 vdd 205 204 vdd hvtpfet l=6e-08 w=4.11e-07 $X=13936 $Y=14280 $D=636
M2106 623 203 200 vdd hvtpfet l=6e-08 w=6e-07 $X=13942 $Y=33468 $D=636
M2107 192 204 1207 vdd hvtpfet l=6e-08 w=4.11e-07 $X=13971 $Y=15932 $D=636
M2108 193 204 1208 vdd hvtpfet l=6e-08 w=4.11e-07 $X=13971 $Y=20589 $D=636
M2109 194 205 1209 vdd hvtpfet l=6e-08 w=4.11e-07 $X=13971 $Y=22852 $D=636
M2110 195 205 1210 vdd hvtpfet l=6e-08 w=4.11e-07 $X=13971 $Y=27509 $D=636
M2111 143 200 620 vdd hvtpfet l=6e-08 w=1e-06 $X=14013 $Y=35707 $D=636
M2112 vdd 206 b_pxcb_n<0> vdd hvtpfet l=6e-08 w=2.57e-06 $X=14050 $Y=1941 $D=636
M2113 vdd 207 206 vdd hvtpfet l=6e-08 w=1e-06 $X=14050 $Y=5141 $D=636
M2114 vdd 189 207 vdd hvtpfet l=6e-08 w=6e-07 $X=14050 $Y=8691 $D=636
M2115 vdd 189 208 vdd hvtpfet l=6e-08 w=6e-07 $X=14050 $Y=41842 $D=636
M2116 vdd 208 209 vdd hvtpfet l=6e-08 w=1e-06 $X=14050 $Y=44992 $D=636
M2117 vdd 209 t_pxcb_n<0> vdd hvtpfet l=6e-08 w=2.57e-06 $X=14050 $Y=46622 $D=636
M2118 vdd 211 623 vdd hvtpfet l=6e-08 w=6e-07 $X=14202 $Y=33468 $D=636
M2119 vdd dwlb<1> 216 vdd hvtpfet l=6e-08 w=4.11e-07 $X=14216 $Y=10156 $D=636
M2120 vdd dwlb<0> 217 vdd hvtpfet l=6e-08 w=4.11e-07 $X=14216 $Y=40566 $D=636
M2121 1211 210 192 vdd hvtpfet l=6e-08 w=4.11e-07 $X=14231 $Y=15932 $D=636
M2122 1212 210 193 vdd hvtpfet l=6e-08 w=4.11e-07 $X=14231 $Y=20589 $D=636
M2123 1213 210 194 vdd hvtpfet l=6e-08 w=4.11e-07 $X=14231 $Y=22852 $D=636
M2124 1214 210 195 vdd hvtpfet l=6e-08 w=4.11e-07 $X=14231 $Y=27509 $D=636
M2125 205 ab<12> vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=14446 $Y=14280 $D=636
M2126 216 212 vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=14476 $Y=10156 $D=636
M2127 217 212 vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=14476 $Y=40566 $D=636
M2128 vdd 33 1211 vdd hvtpfet l=6e-08 w=8.23e-07 $X=14501 $Y=15520 $D=636
M2129 vdd 33 1212 vdd hvtpfet l=6e-08 w=8.23e-07 $X=14501 $Y=20589 $D=636
M2130 vdd 33 1213 vdd hvtpfet l=6e-08 w=8.23e-07 $X=14501 $Y=22440 $D=636
M2131 vdd 33 1214 vdd hvtpfet l=6e-08 w=8.23e-07 $X=14501 $Y=27509 $D=636
M2132 b_pxcb_n<1> 218 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=14560 $Y=1941 $D=636
M2133 218 219 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=14560 $Y=5141 $D=636
M2134 219 190 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=14560 $Y=8691 $D=636
M2135 220 190 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=14560 $Y=41842 $D=636
M2136 221 220 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=14560 $Y=44992 $D=636
M2137 t_pxcb_n<1> 221 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=14560 $Y=46622 $D=636
M2138 vdd 123 624 vdd hvtpfet l=6e-08 w=1.2e-06 $X=14796 $Y=29148 $D=636
M2139 vdd 218 b_pxcb_n<1> vdd hvtpfet l=6e-08 w=2.57e-06 $X=14820 $Y=1941 $D=636
M2140 vdd 219 218 vdd hvtpfet l=6e-08 w=1e-06 $X=14820 $Y=5141 $D=636
M2141 vdd 190 219 vdd hvtpfet l=6e-08 w=6e-07 $X=14820 $Y=8691 $D=636
M2142 vdd 190 220 vdd hvtpfet l=6e-08 w=6e-07 $X=14820 $Y=41842 $D=636
M2143 vdd 220 221 vdd hvtpfet l=6e-08 w=1e-06 $X=14820 $Y=44992 $D=636
M2144 vdd 221 t_pxcb_n<1> vdd hvtpfet l=6e-08 w=2.57e-06 $X=14820 $Y=46622 $D=636
M2145 vdd 72 58 vdd hvtpfet l=6e-08 w=4e-07 $X=14872 $Y=35682 $D=636
M2146 48 216 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=14986 $Y=10167 $D=636
M2147 49 217 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=14986 $Y=40566 $D=636
M2148 1215 213 192 vdd hvtpfet l=6e-08 w=4.11e-07 $X=15011 $Y=15932 $D=636
M2149 1216 214 193 vdd hvtpfet l=6e-08 w=4.11e-07 $X=15011 $Y=20589 $D=636
M2150 1217 213 194 vdd hvtpfet l=6e-08 w=4.11e-07 $X=15011 $Y=22852 $D=636
M2151 1218 214 195 vdd hvtpfet l=6e-08 w=4.11e-07 $X=15011 $Y=27509 $D=636
M2152 33 43 vdd vdd hvtpfet l=6e-08 w=7e-07 $X=15056 $Y=29648 $D=636
M2153 vdd 33 1215 vdd hvtpfet l=6e-08 w=8.23e-07 $X=15281 $Y=15520 $D=636
M2154 vdd 33 1216 vdd hvtpfet l=6e-08 w=8.23e-07 $X=15281 $Y=20589 $D=636
M2155 vdd 33 1217 vdd hvtpfet l=6e-08 w=8.23e-07 $X=15281 $Y=22440 $D=636
M2156 vdd 33 1218 vdd hvtpfet l=6e-08 w=8.23e-07 $X=15281 $Y=27509 $D=636
M2157 vdd 43 33 vdd hvtpfet l=6e-08 w=7e-07 $X=15316 $Y=29648 $D=636
M2158 b_pxcb_n<2> 223 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=15330 $Y=1941 $D=636
M2159 223 224 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=15330 $Y=5141 $D=636
M2160 224 225 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=15330 $Y=8691 $D=636
M2161 226 225 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=15330 $Y=41842 $D=636
M2162 227 226 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=15330 $Y=44992 $D=636
M2163 t_pxcb_n<2> 227 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=15330 $Y=46622 $D=636
M2164 vdd 229 72 vdd hvtpfet l=6e-08 w=4e-07 $X=15382 $Y=35682 $D=636
M2165 vdd ab<11> 210 vdd hvtpfet l=6e-08 w=4.11e-07 $X=15456 $Y=14280 $D=636
M2166 1219 33 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=15541 $Y=15520 $D=636
M2167 1220 33 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=15541 $Y=20589 $D=636
M2168 1221 33 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=15541 $Y=22440 $D=636
M2169 1222 33 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=15541 $Y=27509 $D=636
M2170 33 43 vdd vdd hvtpfet l=6e-08 w=7e-07 $X=15576 $Y=29648 $D=636
M2171 vdd 223 b_pxcb_n<2> vdd hvtpfet l=6e-08 w=2.57e-06 $X=15590 $Y=1941 $D=636
M2172 vdd 224 223 vdd hvtpfet l=6e-08 w=1e-06 $X=15590 $Y=5141 $D=636
M2173 vdd 225 224 vdd hvtpfet l=6e-08 w=6e-07 $X=15590 $Y=8691 $D=636
M2174 vdd 225 226 vdd hvtpfet l=6e-08 w=6e-07 $X=15590 $Y=41842 $D=636
M2175 vdd 226 227 vdd hvtpfet l=6e-08 w=1e-06 $X=15590 $Y=44992 $D=636
M2176 vdd 227 t_pxcb_n<2> vdd hvtpfet l=6e-08 w=2.57e-06 $X=15590 $Y=46622 $D=636
M2177 vdd 228 231 vdd hvtpfet l=6e-08 w=3.2e-07 $X=15621 $Y=33942 $D=636
M2178 72 172 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=15642 $Y=35682 $D=636
M2179 240 210 vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=15716 $Y=14280 $D=636
M2180 249 213 1219 vdd hvtpfet l=6e-08 w=4.11e-07 $X=15811 $Y=15932 $D=636
M2181 250 214 1220 vdd hvtpfet l=6e-08 w=4.11e-07 $X=15811 $Y=20589 $D=636
M2182 251 213 1221 vdd hvtpfet l=6e-08 w=4.11e-07 $X=15811 $Y=22852 $D=636
M2183 252 214 1222 vdd hvtpfet l=6e-08 w=4.11e-07 $X=15811 $Y=27509 $D=636
M2184 vdd 43 33 vdd hvtpfet l=6e-08 w=7e-07 $X=15836 $Y=29648 $D=636
M2185 631 tm<0> vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=15880 $Y=40177 $D=636
M2186 632 123 vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=15881 $Y=33942 $D=636
M2187 vdd tm<3> 242 vdd hvtpfet l=7e-08 w=4.8e-07 $X=16057 $Y=10476 $D=636
M2188 b_pxcb_n<3> 235 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=16100 $Y=1941 $D=636
M2189 235 236 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=16100 $Y=5141 $D=636
M2190 236 237 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=16100 $Y=8691 $D=636
M2191 238 237 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=16100 $Y=41842 $D=636
M2192 239 238 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=16100 $Y=44992 $D=636
M2193 t_pxcb_n<3> 239 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=16100 $Y=46622 $D=636
M2194 228 231 632 vdd hvtpfet l=6e-08 w=3.2e-07 $X=16141 $Y=33942 $D=636
M2195 vdd 213 214 vdd hvtpfet l=6e-08 w=4.11e-07 $X=16316 $Y=14280 $D=636
M2196 1225 33 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=16321 $Y=15520 $D=636
M2197 1226 33 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=16321 $Y=20589 $D=636
M2198 1227 33 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=16321 $Y=22440 $D=636
M2199 1228 33 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=16321 $Y=27509 $D=636
M2200 1223 232 vdd vdd hvtpfet l=6e-08 w=4.8e-07 $X=16322 $Y=35753 $D=636
M2201 243 tm<4> vdd vdd hvtpfet l=7e-08 w=4.8e-07 $X=16327 $Y=10476 $D=636
M2202 642 123 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=16346 $Y=29274 $D=636
M2203 vdd 235 b_pxcb_n<3> vdd hvtpfet l=6e-08 w=2.57e-06 $X=16360 $Y=1941 $D=636
M2204 vdd 236 235 vdd hvtpfet l=6e-08 w=1e-06 $X=16360 $Y=5141 $D=636
M2205 vdd 237 236 vdd hvtpfet l=6e-08 w=6e-07 $X=16360 $Y=8691 $D=636
M2206 vdd 237 238 vdd hvtpfet l=6e-08 w=6e-07 $X=16360 $Y=41842 $D=636
M2207 vdd 238 239 vdd hvtpfet l=6e-08 w=1e-06 $X=16360 $Y=44992 $D=636
M2208 vdd 239 t_pxcb_n<3> vdd hvtpfet l=6e-08 w=2.57e-06 $X=16360 $Y=46622 $D=636
M2209 1224 131 228 vdd hvtpfet l=6e-08 w=4.8e-07 $X=16401 $Y=33942 $D=636
M2210 213 ab<10> vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=16576 $Y=14280 $D=636
M2211 229 172 1223 vdd hvtpfet l=6e-08 w=4.8e-07 $X=16582 $Y=35753 $D=636
M2212 249 240 1225 vdd hvtpfet l=6e-08 w=4.11e-07 $X=16591 $Y=15932 $D=636
M2213 250 240 1226 vdd hvtpfet l=6e-08 w=4.11e-07 $X=16591 $Y=20589 $D=636
M2214 251 240 1227 vdd hvtpfet l=6e-08 w=4.11e-07 $X=16591 $Y=22852 $D=636
M2215 252 240 1228 vdd hvtpfet l=6e-08 w=4.11e-07 $X=16591 $Y=27509 $D=636
M2216 vdd 123 642 vdd hvtpfet l=6e-08 w=6e-07 $X=16606 $Y=29274 $D=636
M2217 vdd 123 1224 vdd hvtpfet l=6e-08 w=4.8e-07 $X=16661 $Y=33942 $D=636
M2218 637 tm<6> vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=16680 $Y=40177 $D=636
M2219 639 244 229 vdd hvtpfet l=6e-08 w=3.2e-07 $X=16842 $Y=35913 $D=636
M2220 1229 243 643 vdd hvtpfet l=6e-08 w=4.8e-07 $X=16847 $Y=10476 $D=636
M2221 1230 204 249 vdd hvtpfet l=6e-08 w=4.11e-07 $X=16851 $Y=15932 $D=636
M2222 1231 204 250 vdd hvtpfet l=6e-08 w=4.11e-07 $X=16851 $Y=20589 $D=636
M2223 1232 205 251 vdd hvtpfet l=6e-08 w=4.11e-07 $X=16851 $Y=22852 $D=636
M2224 1233 205 252 vdd hvtpfet l=6e-08 w=4.11e-07 $X=16851 $Y=27509 $D=636
M2225 642 123 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=16866 $Y=29274 $D=636
M2226 b_pxcb_n<4> 245 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=16870 $Y=1941 $D=636
M2227 245 246 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=16870 $Y=5141 $D=636
M2228 246 187 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=16870 $Y=8691 $D=636
M2229 247 187 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=16870 $Y=41842 $D=636
M2230 248 247 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=16870 $Y=44992 $D=636
M2231 t_pxcb_n<4> 248 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=16870 $Y=46622 $D=636
M2232 vdd 142 639 vdd hvtpfet l=6e-08 w=3.2e-07 $X=17102 $Y=35913 $D=636
M2233 vdd 242 1229 vdd hvtpfet l=6e-08 w=4.8e-07 $X=17107 $Y=10476 $D=636
M2234 vdd 33 1230 vdd hvtpfet l=6e-08 w=8.23e-07 $X=17121 $Y=15520 $D=636
M2235 vdd 33 1231 vdd hvtpfet l=6e-08 w=8.23e-07 $X=17121 $Y=20589 $D=636
M2236 vdd 33 1232 vdd hvtpfet l=6e-08 w=8.23e-07 $X=17121 $Y=22440 $D=636
M2237 vdd 33 1233 vdd hvtpfet l=6e-08 w=8.23e-07 $X=17121 $Y=27509 $D=636
M2238 vdd 123 642 vdd hvtpfet l=6e-08 w=6e-07 $X=17126 $Y=29274 $D=636
M2239 vdd 245 b_pxcb_n<4> vdd hvtpfet l=6e-08 w=2.57e-06 $X=17130 $Y=1941 $D=636
M2240 vdd 246 245 vdd hvtpfet l=6e-08 w=1e-06 $X=17130 $Y=5141 $D=636
M2241 vdd 187 246 vdd hvtpfet l=6e-08 w=6e-07 $X=17130 $Y=8691 $D=636
M2242 vdd 187 247 vdd hvtpfet l=6e-08 w=6e-07 $X=17130 $Y=41842 $D=636
M2243 vdd 247 248 vdd hvtpfet l=6e-08 w=1e-06 $X=17130 $Y=44992 $D=636
M2244 vdd 248 t_pxcb_n<4> vdd hvtpfet l=6e-08 w=2.57e-06 $X=17130 $Y=46622 $D=636
M2245 244 229 vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=17362 $Y=35913 $D=636
M2246 1234 242 vdd vdd hvtpfet l=6e-08 w=4.8e-07 $X=17617 $Y=10476 $D=636
M2247 253 249 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=17631 $Y=15321 $D=636
M2248 1235 43 249 vdd hvtpfet l=6e-08 w=2.74e-07 $X=17631 $Y=16069 $D=636
M2249 1236 43 250 vdd hvtpfet l=6e-08 w=2.74e-07 $X=17631 $Y=20589 $D=636
M2250 254 250 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=17631 $Y=21405 $D=636
M2251 225 251 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=17631 $Y=22241 $D=636
M2252 1237 43 251 vdd hvtpfet l=6e-08 w=2.74e-07 $X=17631 $Y=22989 $D=636
M2253 1238 43 252 vdd hvtpfet l=6e-08 w=2.74e-07 $X=17631 $Y=27509 $D=636
M2254 237 252 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=17631 $Y=28325 $D=636
M2255 b_pxcb_n<5> 255 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=17640 $Y=1941 $D=636
M2256 255 256 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=17640 $Y=5141 $D=636
M2257 256 188 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=17640 $Y=8691 $D=636
M2258 257 188 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=17640 $Y=41842 $D=636
M2259 258 257 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=17640 $Y=44992 $D=636
M2260 t_pxcb_n<5> 258 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=17640 $Y=46622 $D=636
M2261 23 clkb vdd vdd hvtpfet l=6e-08 w=9e-07 $X=17646 $Y=29274 $D=636
M2262 647 tm<4> 1234 vdd hvtpfet l=6e-08 w=4.8e-07 $X=17877 $Y=10476 $D=636
M2263 vdd 249 253 vdd hvtpfet l=6e-08 w=2.06e-07 $X=17891 $Y=15321 $D=636
M2264 vdd 253 1235 vdd hvtpfet l=6e-08 w=2.74e-07 $X=17891 $Y=16069 $D=636
M2265 vdd 254 1236 vdd hvtpfet l=6e-08 w=2.74e-07 $X=17891 $Y=20589 $D=636
M2266 vdd 250 254 vdd hvtpfet l=6e-08 w=2.06e-07 $X=17891 $Y=21405 $D=636
M2267 vdd 251 225 vdd hvtpfet l=6e-08 w=2.06e-07 $X=17891 $Y=22241 $D=636
M2268 vdd 225 1237 vdd hvtpfet l=6e-08 w=2.74e-07 $X=17891 $Y=22989 $D=636
M2269 vdd 237 1238 vdd hvtpfet l=6e-08 w=2.74e-07 $X=17891 $Y=27509 $D=636
M2270 vdd 252 237 vdd hvtpfet l=6e-08 w=2.06e-07 $X=17891 $Y=28325 $D=636
M2271 vdd 255 b_pxcb_n<5> vdd hvtpfet l=6e-08 w=2.57e-06 $X=17900 $Y=1941 $D=636
M2272 vdd 256 255 vdd hvtpfet l=6e-08 w=1e-06 $X=17900 $Y=5141 $D=636
M2273 vdd 188 256 vdd hvtpfet l=6e-08 w=6e-07 $X=17900 $Y=8691 $D=636
M2274 vdd 188 257 vdd hvtpfet l=6e-08 w=6e-07 $X=17900 $Y=41842 $D=636
M2275 vdd 257 258 vdd hvtpfet l=6e-08 w=1e-06 $X=17900 $Y=44992 $D=636
M2276 vdd 258 t_pxcb_n<5> vdd hvtpfet l=6e-08 w=2.57e-06 $X=17900 $Y=46622 $D=636
M2277 vdd 260 273 vdd hvtpfet l=6e-08 w=4.11e-07 $X=18106 $Y=14280 $D=636
M2278 1239 wenb 232 vdd hvtpfet l=6e-08 w=8e-07 $X=18366 $Y=35907 $D=636
M2279 1240 tm<4> 648 vdd hvtpfet l=6e-08 w=4.8e-07 $X=18387 $Y=10476 $D=636
M2280 b_pxcb_n<6> 265 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=18410 $Y=1941 $D=636
M2281 265 266 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=18410 $Y=5141 $D=636
M2282 266 253 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=18410 $Y=8691 $D=636
M2283 267 253 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=18410 $Y=41842 $D=636
M2284 268 267 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=18410 $Y=44992 $D=636
M2285 t_pxcb_n<6> 268 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=18410 $Y=46622 $D=636
M2286 1241 ab<4> vdd vdd hvtpfet l=6e-08 w=4.8e-07 $X=18460 $Y=29394 $D=636
M2287 1242 wenb vdd vdd hvtpfet l=6e-08 w=4.8e-07 $X=18460 $Y=33942 $D=636
M2288 vdd tm<2> 173 vdd hvtpfet l=6e-08 w=4.11e-07 $X=18510 $Y=40177 $D=636
M2289 260 ab<1> vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=18616 $Y=14280 $D=636
M2290 vdd 264 1239 vdd hvtpfet l=6e-08 w=8e-07 $X=18626 $Y=35907 $D=636
M2291 1243 33 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=18641 $Y=15520 $D=636
M2292 1244 33 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=18641 $Y=20589 $D=636
M2293 1245 33 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=18641 $Y=22440 $D=636
M2294 1246 33 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=18641 $Y=27509 $D=636
M2295 vdd tm<3> 1240 vdd hvtpfet l=6e-08 w=4.8e-07 $X=18647 $Y=10476 $D=636
M2296 vdd 265 b_pxcb_n<6> vdd hvtpfet l=6e-08 w=2.57e-06 $X=18670 $Y=1941 $D=636
M2297 vdd 266 265 vdd hvtpfet l=6e-08 w=1e-06 $X=18670 $Y=5141 $D=636
M2298 vdd 253 266 vdd hvtpfet l=6e-08 w=6e-07 $X=18670 $Y=8691 $D=636
M2299 vdd 253 267 vdd hvtpfet l=6e-08 w=6e-07 $X=18670 $Y=41842 $D=636
M2300 vdd 267 268 vdd hvtpfet l=6e-08 w=1e-06 $X=18670 $Y=44992 $D=636
M2301 vdd 268 t_pxcb_n<6> vdd hvtpfet l=6e-08 w=2.57e-06 $X=18670 $Y=46622 $D=636
M2302 154 clkb 1241 vdd hvtpfet l=6e-08 w=4.8e-07 $X=18720 $Y=29394 $D=636
M2303 274 clkb 1242 vdd hvtpfet l=6e-08 w=4.8e-07 $X=18720 $Y=33942 $D=636
M2304 280 269 1243 vdd hvtpfet l=6e-08 w=4.11e-07 $X=18911 $Y=15932 $D=636
M2305 281 270 1244 vdd hvtpfet l=6e-08 w=4.11e-07 $X=18911 $Y=20589 $D=636
M2306 282 269 1245 vdd hvtpfet l=6e-08 w=4.11e-07 $X=18911 $Y=22852 $D=636
M2307 283 270 1246 vdd hvtpfet l=6e-08 w=4.11e-07 $X=18911 $Y=27509 $D=636
M2308 655 271 154 vdd hvtpfet l=6e-08 w=3.2e-07 $X=18980 $Y=29554 $D=636
M2309 656 272 274 vdd hvtpfet l=6e-08 w=3.2e-07 $X=18980 $Y=33942 $D=636
M2310 vdd 270 269 vdd hvtpfet l=6e-08 w=4.11e-07 $X=19126 $Y=14280 $D=636
M2311 1247 tm<3> vdd vdd hvtpfet l=6e-08 w=4.8e-07 $X=19157 $Y=10476 $D=636
M2312 1248 273 280 vdd hvtpfet l=6e-08 w=4.11e-07 $X=19171 $Y=15932 $D=636
M2313 1249 273 281 vdd hvtpfet l=6e-08 w=4.11e-07 $X=19171 $Y=20589 $D=636
M2314 1250 260 282 vdd hvtpfet l=6e-08 w=4.11e-07 $X=19171 $Y=22852 $D=636
M2315 1251 260 283 vdd hvtpfet l=6e-08 w=4.11e-07 $X=19171 $Y=27509 $D=636
M2316 b_pxcb_n<7> 275 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=19180 $Y=1941 $D=636
M2317 275 276 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=19180 $Y=5141 $D=636
M2318 276 254 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=19180 $Y=8691 $D=636
M2319 277 254 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=19180 $Y=41842 $D=636
M2320 278 277 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=19180 $Y=44992 $D=636
M2321 t_pxcb_n<7> 278 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=19180 $Y=46622 $D=636
M2322 vdd 23 655 vdd hvtpfet l=6e-08 w=3.2e-07 $X=19240 $Y=29554 $D=636
M2323 vdd 23 656 vdd hvtpfet l=6e-08 w=3.2e-07 $X=19240 $Y=33942 $D=636
M2324 659 243 1247 vdd hvtpfet l=6e-08 w=4.8e-07 $X=19417 $Y=10476 $D=636
M2325 vdd 275 b_pxcb_n<7> vdd hvtpfet l=6e-08 w=2.57e-06 $X=19440 $Y=1941 $D=636
M2326 vdd 276 275 vdd hvtpfet l=6e-08 w=1e-06 $X=19440 $Y=5141 $D=636
M2327 vdd 254 276 vdd hvtpfet l=6e-08 w=6e-07 $X=19440 $Y=8691 $D=636
M2328 vdd 254 277 vdd hvtpfet l=6e-08 w=6e-07 $X=19440 $Y=41842 $D=636
M2329 vdd 277 278 vdd hvtpfet l=6e-08 w=1e-06 $X=19440 $Y=44992 $D=636
M2330 vdd 278 t_pxcb_n<7> vdd hvtpfet l=6e-08 w=2.57e-06 $X=19440 $Y=46622 $D=636
M2331 vdd 33 1248 vdd hvtpfet l=6e-08 w=8.23e-07 $X=19441 $Y=15520 $D=636
M2332 vdd 33 1249 vdd hvtpfet l=6e-08 w=8.23e-07 $X=19441 $Y=20589 $D=636
M2333 vdd 33 1250 vdd hvtpfet l=6e-08 w=8.23e-07 $X=19441 $Y=22440 $D=636
M2334 vdd 33 1251 vdd hvtpfet l=6e-08 w=8.23e-07 $X=19441 $Y=27509 $D=636
M2335 271 154 vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=19500 $Y=29554 $D=636
M2336 272 274 vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=19500 $Y=33942 $D=636
M2337 270 ab<0> vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=19636 $Y=14280 $D=636
M2338 vdd 15 r_saeb_n vdd hvtpfet l=6e-08 w=1.43e-06 $X=19675 $Y=35277 $D=636
M2339 r_saeb_n 15 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=19935 $Y=35277 $D=636
M2340 212 280 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=19951 $Y=15321 $D=636
M2341 1252 43 280 vdd hvtpfet l=6e-08 w=2.74e-07 $X=19951 $Y=16069 $D=636
M2342 1253 43 281 vdd hvtpfet l=6e-08 w=2.74e-07 $X=19951 $Y=20589 $D=636
M2343 185 281 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=19951 $Y=21405 $D=636
M2344 155 282 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=19951 $Y=22241 $D=636
M2345 1254 43 282 vdd hvtpfet l=6e-08 w=2.74e-07 $X=19951 $Y=22989 $D=636
M2346 1255 43 283 vdd hvtpfet l=6e-08 w=2.74e-07 $X=19951 $Y=27509 $D=636
M2347 145 283 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=19951 $Y=28325 $D=636
M2348 vdd 11 rb_cb<0> vdd hvtpfet l=6e-08 w=1.43e-06 $X=20195 $Y=1506 $D=636
M2349 vdd 12 rb_cb<2> vdd hvtpfet l=6e-08 w=1.43e-06 $X=20195 $Y=3566 $D=636
M2350 vdd 13 rb_mb<0> vdd hvtpfet l=6e-08 w=1.43e-06 $X=20195 $Y=7966 $D=636
M2351 vdd 14 rb_mb<2> vdd hvtpfet l=6e-08 w=1.43e-06 $X=20195 $Y=10026 $D=636
M2352 vdd 15 r_saeb_n vdd hvtpfet l=6e-08 w=1.43e-06 $X=20195 $Y=35277 $D=636
M2353 vdd 16 rt_mb<2> vdd hvtpfet l=6e-08 w=1.43e-06 $X=20195 $Y=39677 $D=636
M2354 vdd 17 rt_mb<0> vdd hvtpfet l=6e-08 w=1.43e-06 $X=20195 $Y=41737 $D=636
M2355 vdd 18 rt_cb<2> vdd hvtpfet l=6e-08 w=1.43e-06 $X=20195 $Y=46137 $D=636
M2356 vdd 19 rt_cb<0> vdd hvtpfet l=6e-08 w=1.43e-06 $X=20195 $Y=48197 $D=636
M2357 vdd 280 212 vdd hvtpfet l=6e-08 w=2.06e-07 $X=20211 $Y=15321 $D=636
M2358 vdd 212 1252 vdd hvtpfet l=6e-08 w=2.74e-07 $X=20211 $Y=16069 $D=636
M2359 vdd 185 1253 vdd hvtpfet l=6e-08 w=2.74e-07 $X=20211 $Y=20589 $D=636
M2360 vdd 281 185 vdd hvtpfet l=6e-08 w=2.06e-07 $X=20211 $Y=21405 $D=636
M2361 vdd 282 155 vdd hvtpfet l=6e-08 w=2.06e-07 $X=20211 $Y=22241 $D=636
M2362 vdd 155 1254 vdd hvtpfet l=6e-08 w=2.74e-07 $X=20211 $Y=22989 $D=636
M2363 vdd 145 1255 vdd hvtpfet l=6e-08 w=2.74e-07 $X=20211 $Y=27509 $D=636
M2364 vdd 283 145 vdd hvtpfet l=6e-08 w=2.06e-07 $X=20211 $Y=28325 $D=636
M2365 rb_cb<0> 11 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=20455 $Y=1506 $D=636
M2366 rb_cb<2> 12 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=20455 $Y=3566 $D=636
M2367 rb_mb<0> 13 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=20455 $Y=7966 $D=636
M2368 rb_mb<2> 14 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=20455 $Y=10026 $D=636
M2369 r_saeb_n 15 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=20455 $Y=35277 $D=636
M2370 rt_mb<2> 16 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=20455 $Y=39677 $D=636
M2371 rt_mb<0> 17 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=20455 $Y=41737 $D=636
M2372 rt_cb<2> 18 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=20455 $Y=46137 $D=636
M2373 rt_cb<0> 19 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=20455 $Y=48197 $D=636
M2374 vdd 11 rb_cb<0> vdd hvtpfet l=6e-08 w=1.43e-06 $X=20715 $Y=1506 $D=636
M2375 vdd 12 rb_cb<2> vdd hvtpfet l=6e-08 w=1.43e-06 $X=20715 $Y=3566 $D=636
M2376 vdd 13 rb_mb<0> vdd hvtpfet l=6e-08 w=1.43e-06 $X=20715 $Y=7966 $D=636
M2377 vdd 14 rb_mb<2> vdd hvtpfet l=6e-08 w=1.43e-06 $X=20715 $Y=10026 $D=636
M2378 vdd 15 r_saeb_n vdd hvtpfet l=6e-08 w=1.43e-06 $X=20715 $Y=35277 $D=636
M2379 vdd 16 rt_mb<2> vdd hvtpfet l=6e-08 w=1.43e-06 $X=20715 $Y=39677 $D=636
M2380 vdd 17 rt_mb<0> vdd hvtpfet l=6e-08 w=1.43e-06 $X=20715 $Y=41737 $D=636
M2381 vdd 18 rt_cb<2> vdd hvtpfet l=6e-08 w=1.43e-06 $X=20715 $Y=46137 $D=636
M2382 vdd 19 rt_cb<0> vdd hvtpfet l=6e-08 w=1.43e-06 $X=20715 $Y=48197 $D=636
M2383 10 274 vdd vdd hvtpfet l=6e-08 w=1.2e-06 $X=20725 $Y=32684 $D=636
M2384 rb_cb<1> 34 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=20975 $Y=1506 $D=636
M2385 rb_cb<3> 35 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=20975 $Y=3566 $D=636
M2386 rb_mb<1> 36 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=20975 $Y=7966 $D=636
M2387 rb_mb<3> 37 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=20975 $Y=10026 $D=636
M2388 r_clk_dqb 8 vdd vdd hvtpfet l=6e-08 w=2.1e-06 $X=20975 $Y=23696 $D=636
M2389 r_clk_dqb_n 9 vdd vdd hvtpfet l=6e-08 w=2.1e-06 $X=20975 $Y=26512 $D=636
M2390 r_sa_preb_n 51 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=20975 $Y=35277 $D=636
M2391 rt_mb<3> 39 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=20975 $Y=39677 $D=636
M2392 rt_mb<1> 40 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=20975 $Y=41737 $D=636
M2393 rt_cb<3> 41 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=20975 $Y=46137 $D=636
M2394 rt_cb<1> 42 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=20975 $Y=48197 $D=636
M2395 vdd 34 rb_cb<1> vdd hvtpfet l=6e-08 w=1.43e-06 $X=21235 $Y=1506 $D=636
M2396 vdd 35 rb_cb<3> vdd hvtpfet l=6e-08 w=1.43e-06 $X=21235 $Y=3566 $D=636
M2397 vdd 36 rb_mb<1> vdd hvtpfet l=6e-08 w=1.43e-06 $X=21235 $Y=7966 $D=636
M2398 vdd 37 rb_mb<3> vdd hvtpfet l=6e-08 w=1.43e-06 $X=21235 $Y=10026 $D=636
M2399 rb_tm_preb_n 20 vdd vdd hvtpfet l=6e-08 w=2.145e-06 $X=21235 $Y=14887 $D=636
M2400 rt_tm_preb_n 21 vdd vdd hvtpfet l=6e-08 w=2.145e-06 $X=21235 $Y=17659 $D=636
M2401 vdd 8 r_clk_dqb vdd hvtpfet l=6e-08 w=2.1e-06 $X=21235 $Y=23696 $D=636
M2402 vdd 9 r_clk_dqb_n vdd hvtpfet l=6e-08 w=2.1e-06 $X=21235 $Y=26512 $D=636
M2403 r_lweb 10 vdd vdd hvtpfet l=6e-08 w=2.145e-06 $X=21235 $Y=32504 $D=636
M2404 vdd 51 r_sa_preb_n vdd hvtpfet l=6e-08 w=1.43e-06 $X=21235 $Y=35277 $D=636
M2405 vdd 39 rt_mb<3> vdd hvtpfet l=6e-08 w=1.43e-06 $X=21235 $Y=39677 $D=636
M2406 vdd 40 rt_mb<1> vdd hvtpfet l=6e-08 w=1.43e-06 $X=21235 $Y=41737 $D=636
M2407 vdd 41 rt_cb<3> vdd hvtpfet l=6e-08 w=1.43e-06 $X=21235 $Y=46137 $D=636
M2408 vdd 42 rt_cb<1> vdd hvtpfet l=6e-08 w=1.43e-06 $X=21235 $Y=48197 $D=636
M2409 rb_cb<1> 34 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=21495 $Y=1506 $D=636
M2410 rb_cb<3> 35 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=21495 $Y=3566 $D=636
M2411 rb_mb<1> 36 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=21495 $Y=7966 $D=636
M2412 rb_mb<3> 37 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=21495 $Y=10026 $D=636
M2413 vdd 20 rb_tm_preb_n vdd hvtpfet l=6e-08 w=2.145e-06 $X=21495 $Y=14887 $D=636
M2414 vdd 21 rt_tm_preb_n vdd hvtpfet l=6e-08 w=2.145e-06 $X=21495 $Y=17659 $D=636
M2415 r_clk_dqb 8 vdd vdd hvtpfet l=6e-08 w=2.1e-06 $X=21495 $Y=23696 $D=636
M2416 r_clk_dqb_n 9 vdd vdd hvtpfet l=6e-08 w=2.1e-06 $X=21495 $Y=26512 $D=636
M2417 vdd 10 r_lweb vdd hvtpfet l=6e-08 w=2.145e-06 $X=21495 $Y=32504 $D=636
M2418 r_sa_preb_n 51 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=21495 $Y=35277 $D=636
M2419 rt_mb<3> 39 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=21495 $Y=39677 $D=636
M2420 rt_mb<1> 40 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=21495 $Y=41737 $D=636
M2421 rt_cb<3> 41 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=21495 $Y=46137 $D=636
M2422 rt_cb<1> 42 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=21495 $Y=48197 $D=636
M2423 vdd 289 lb_ca<1> vdd hvtpfet l=6e-08 w=1.43e-06 $X=22005 $Y=1506 $D=636
M2424 vdd 290 lb_ca<3> vdd hvtpfet l=6e-08 w=1.43e-06 $X=22005 $Y=3566 $D=636
M2425 vdd 291 lb_ma<1> vdd hvtpfet l=6e-08 w=1.43e-06 $X=22005 $Y=7966 $D=636
M2426 vdd 292 lb_ma<3> vdd hvtpfet l=6e-08 w=1.43e-06 $X=22005 $Y=10026 $D=636
M2427 lb_tm_prea_n 285 vdd vdd hvtpfet l=6e-08 w=2.145e-06 $X=22005 $Y=14887 $D=636
M2428 lt_tm_prea_n 286 vdd vdd hvtpfet l=6e-08 w=2.145e-06 $X=22005 $Y=17659 $D=636
M2429 vdd 287 l_clk_dqa vdd hvtpfet l=6e-08 w=2.1e-06 $X=22005 $Y=23696 $D=636
M2430 vdd 288 l_clk_dqa_n vdd hvtpfet l=6e-08 w=2.1e-06 $X=22005 $Y=26512 $D=636
M2431 l_lwea 284 vdd vdd hvtpfet l=6e-08 w=2.145e-06 $X=22005 $Y=32504 $D=636
M2432 vdd 293 l_sa_prea_n vdd hvtpfet l=6e-08 w=1.43e-06 $X=22005 $Y=35277 $D=636
M2433 vdd 294 lt_ma<3> vdd hvtpfet l=6e-08 w=1.43e-06 $X=22005 $Y=39677 $D=636
M2434 vdd 295 lt_ma<1> vdd hvtpfet l=6e-08 w=1.43e-06 $X=22005 $Y=41737 $D=636
M2435 vdd 296 lt_ca<3> vdd hvtpfet l=6e-08 w=1.43e-06 $X=22005 $Y=46137 $D=636
M2436 vdd 297 lt_ca<1> vdd hvtpfet l=6e-08 w=1.43e-06 $X=22005 $Y=48197 $D=636
M2437 lb_ca<1> 289 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=22265 $Y=1506 $D=636
M2438 lb_ca<3> 290 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=22265 $Y=3566 $D=636
M2439 lb_ma<1> 291 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=22265 $Y=7966 $D=636
M2440 lb_ma<3> 292 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=22265 $Y=10026 $D=636
M2441 vdd 285 lb_tm_prea_n vdd hvtpfet l=6e-08 w=2.145e-06 $X=22265 $Y=14887 $D=636
M2442 vdd 286 lt_tm_prea_n vdd hvtpfet l=6e-08 w=2.145e-06 $X=22265 $Y=17659 $D=636
M2443 l_clk_dqa 287 vdd vdd hvtpfet l=6e-08 w=2.1e-06 $X=22265 $Y=23696 $D=636
M2444 l_clk_dqa_n 288 vdd vdd hvtpfet l=6e-08 w=2.1e-06 $X=22265 $Y=26512 $D=636
M2445 vdd 284 l_lwea vdd hvtpfet l=6e-08 w=2.145e-06 $X=22265 $Y=32504 $D=636
M2446 l_sa_prea_n 293 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=22265 $Y=35277 $D=636
M2447 lt_ma<3> 294 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=22265 $Y=39677 $D=636
M2448 lt_ma<1> 295 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=22265 $Y=41737 $D=636
M2449 lt_ca<3> 296 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=22265 $Y=46137 $D=636
M2450 lt_ca<1> 297 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=22265 $Y=48197 $D=636
M2451 vdd 289 lb_ca<1> vdd hvtpfet l=6e-08 w=1.43e-06 $X=22525 $Y=1506 $D=636
M2452 vdd 290 lb_ca<3> vdd hvtpfet l=6e-08 w=1.43e-06 $X=22525 $Y=3566 $D=636
M2453 vdd 291 lb_ma<1> vdd hvtpfet l=6e-08 w=1.43e-06 $X=22525 $Y=7966 $D=636
M2454 vdd 292 lb_ma<3> vdd hvtpfet l=6e-08 w=1.43e-06 $X=22525 $Y=10026 $D=636
M2455 vdd 287 l_clk_dqa vdd hvtpfet l=6e-08 w=2.1e-06 $X=22525 $Y=23696 $D=636
M2456 vdd 288 l_clk_dqa_n vdd hvtpfet l=6e-08 w=2.1e-06 $X=22525 $Y=26512 $D=636
M2457 vdd 293 l_sa_prea_n vdd hvtpfet l=6e-08 w=1.43e-06 $X=22525 $Y=35277 $D=636
M2458 vdd 294 lt_ma<3> vdd hvtpfet l=6e-08 w=1.43e-06 $X=22525 $Y=39677 $D=636
M2459 vdd 295 lt_ma<1> vdd hvtpfet l=6e-08 w=1.43e-06 $X=22525 $Y=41737 $D=636
M2460 vdd 296 lt_ca<3> vdd hvtpfet l=6e-08 w=1.43e-06 $X=22525 $Y=46137 $D=636
M2461 vdd 297 lt_ca<1> vdd hvtpfet l=6e-08 w=1.43e-06 $X=22525 $Y=48197 $D=636
M2462 vdd 298 284 vdd hvtpfet l=6e-08 w=1.2e-06 $X=22775 $Y=32684 $D=636
M2463 lb_ca<0> 299 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=22785 $Y=1506 $D=636
M2464 lb_ca<2> 300 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=22785 $Y=3566 $D=636
M2465 lb_ma<0> 301 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=22785 $Y=7966 $D=636
M2466 lb_ma<2> 302 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=22785 $Y=10026 $D=636
M2467 l_saea_n 303 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=22785 $Y=35277 $D=636
M2468 lt_ma<2> 304 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=22785 $Y=39677 $D=636
M2469 lt_ma<0> 305 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=22785 $Y=41737 $D=636
M2470 lt_ca<2> 306 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=22785 $Y=46137 $D=636
M2471 lt_ca<0> 307 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=22785 $Y=48197 $D=636
M2472 vdd 299 lb_ca<0> vdd hvtpfet l=6e-08 w=1.43e-06 $X=23045 $Y=1506 $D=636
M2473 vdd 300 lb_ca<2> vdd hvtpfet l=6e-08 w=1.43e-06 $X=23045 $Y=3566 $D=636
M2474 vdd 301 lb_ma<0> vdd hvtpfet l=6e-08 w=1.43e-06 $X=23045 $Y=7966 $D=636
M2475 vdd 302 lb_ma<2> vdd hvtpfet l=6e-08 w=1.43e-06 $X=23045 $Y=10026 $D=636
M2476 vdd 303 l_saea_n vdd hvtpfet l=6e-08 w=1.43e-06 $X=23045 $Y=35277 $D=636
M2477 vdd 304 lt_ma<2> vdd hvtpfet l=6e-08 w=1.43e-06 $X=23045 $Y=39677 $D=636
M2478 vdd 305 lt_ma<0> vdd hvtpfet l=6e-08 w=1.43e-06 $X=23045 $Y=41737 $D=636
M2479 vdd 306 lt_ca<2> vdd hvtpfet l=6e-08 w=1.43e-06 $X=23045 $Y=46137 $D=636
M2480 vdd 307 lt_ca<0> vdd hvtpfet l=6e-08 w=1.43e-06 $X=23045 $Y=48197 $D=636
M2481 308 312 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=23289 $Y=15321 $D=636
M2482 1256 308 vdd vdd hvtpfet l=6e-08 w=2.74e-07 $X=23289 $Y=16069 $D=636
M2483 1257 309 vdd vdd hvtpfet l=6e-08 w=2.74e-07 $X=23289 $Y=20589 $D=636
M2484 309 313 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=23289 $Y=21405 $D=636
M2485 310 314 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=23289 $Y=22241 $D=636
M2486 1258 310 vdd vdd hvtpfet l=6e-08 w=2.74e-07 $X=23289 $Y=22989 $D=636
M2487 1259 311 vdd vdd hvtpfet l=6e-08 w=2.74e-07 $X=23289 $Y=27509 $D=636
M2488 311 315 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=23289 $Y=28325 $D=636
M2489 lb_ca<0> 299 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=23305 $Y=1506 $D=636
M2490 lb_ca<2> 300 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=23305 $Y=3566 $D=636
M2491 lb_ma<0> 301 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=23305 $Y=7966 $D=636
M2492 lb_ma<2> 302 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=23305 $Y=10026 $D=636
M2493 l_saea_n 303 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=23305 $Y=35277 $D=636
M2494 lt_ma<2> 304 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=23305 $Y=39677 $D=636
M2495 lt_ma<0> 305 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=23305 $Y=41737 $D=636
M2496 lt_ca<2> 306 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=23305 $Y=46137 $D=636
M2497 lt_ca<0> 307 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=23305 $Y=48197 $D=636
M2498 vdd 312 308 vdd hvtpfet l=6e-08 w=2.06e-07 $X=23549 $Y=15321 $D=636
M2499 312 323 1256 vdd hvtpfet l=6e-08 w=2.74e-07 $X=23549 $Y=16069 $D=636
M2500 313 323 1257 vdd hvtpfet l=6e-08 w=2.74e-07 $X=23549 $Y=20589 $D=636
M2501 vdd 313 309 vdd hvtpfet l=6e-08 w=2.06e-07 $X=23549 $Y=21405 $D=636
M2502 vdd 314 310 vdd hvtpfet l=6e-08 w=2.06e-07 $X=23549 $Y=22241 $D=636
M2503 314 323 1258 vdd hvtpfet l=6e-08 w=2.74e-07 $X=23549 $Y=22989 $D=636
M2504 315 323 1259 vdd hvtpfet l=6e-08 w=2.74e-07 $X=23549 $Y=27509 $D=636
M2505 vdd 315 311 vdd hvtpfet l=6e-08 w=2.06e-07 $X=23549 $Y=28325 $D=636
M2506 vdd 303 l_saea_n vdd hvtpfet l=6e-08 w=1.43e-06 $X=23565 $Y=35277 $D=636
M2507 l_saea_n 303 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=23825 $Y=35277 $D=636
M2508 vdd aa<0> 327 vdd hvtpfet l=6e-08 w=4.11e-07 $X=23864 $Y=14280 $D=636
M2509 vdd 324 331 vdd hvtpfet l=6e-08 w=3.2e-07 $X=24000 $Y=29554 $D=636
M2510 vdd 298 332 vdd hvtpfet l=6e-08 w=3.2e-07 $X=24000 $Y=33942 $D=636
M2511 1261 317 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=24059 $Y=15520 $D=636
M2512 1262 317 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=24059 $Y=20589 $D=636
M2513 1263 317 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=24059 $Y=22440 $D=636
M2514 1264 317 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=24059 $Y=27509 $D=636
M2515 b_pxca_n<7> 318 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=24060 $Y=1941 $D=636
M2516 318 319 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=24060 $Y=5141 $D=636
M2517 319 320 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=24060 $Y=8691 $D=636
M2518 321 320 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=24060 $Y=41842 $D=636
M2519 322 321 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=24060 $Y=44992 $D=636
M2520 t_pxca_n<7> 322 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=24060 $Y=46622 $D=636
M2521 1260 325 709 vdd hvtpfet l=6e-08 w=4.8e-07 $X=24083 $Y=10476 $D=636
M2522 712 340 vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=24260 $Y=29554 $D=636
M2523 713 340 vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=24260 $Y=33942 $D=636
M2524 vdd 318 b_pxca_n<7> vdd hvtpfet l=6e-08 w=2.57e-06 $X=24320 $Y=1941 $D=636
M2525 vdd 319 318 vdd hvtpfet l=6e-08 w=1e-06 $X=24320 $Y=5141 $D=636
M2526 vdd 320 319 vdd hvtpfet l=6e-08 w=6e-07 $X=24320 $Y=8691 $D=636
M2527 vdd 320 321 vdd hvtpfet l=6e-08 w=6e-07 $X=24320 $Y=41842 $D=636
M2528 vdd 321 322 vdd hvtpfet l=6e-08 w=1e-06 $X=24320 $Y=44992 $D=636
M2529 vdd 322 t_pxca_n<7> vdd hvtpfet l=6e-08 w=2.57e-06 $X=24320 $Y=46622 $D=636
M2530 312 328 1261 vdd hvtpfet l=6e-08 w=4.11e-07 $X=24329 $Y=15932 $D=636
M2531 313 328 1262 vdd hvtpfet l=6e-08 w=4.11e-07 $X=24329 $Y=20589 $D=636
M2532 314 329 1263 vdd hvtpfet l=6e-08 w=4.11e-07 $X=24329 $Y=22852 $D=636
M2533 315 329 1264 vdd hvtpfet l=6e-08 w=4.11e-07 $X=24329 $Y=27509 $D=636
M2534 vdd tm<8> 1260 vdd hvtpfet l=6e-08 w=4.8e-07 $X=24343 $Y=10476 $D=636
M2535 334 327 vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=24374 $Y=14280 $D=636
M2536 vdd tm<5> 264 vdd hvtpfet l=6e-08 w=4.11e-07 $X=24518 $Y=40177 $D=636
M2537 324 331 712 vdd hvtpfet l=6e-08 w=3.2e-07 $X=24520 $Y=29554 $D=636
M2538 298 332 713 vdd hvtpfet l=6e-08 w=3.2e-07 $X=24520 $Y=33942 $D=636
M2539 1265 334 312 vdd hvtpfet l=6e-08 w=4.11e-07 $X=24589 $Y=15932 $D=636
M2540 1266 327 313 vdd hvtpfet l=6e-08 w=4.11e-07 $X=24589 $Y=20589 $D=636
M2541 1267 334 314 vdd hvtpfet l=6e-08 w=4.11e-07 $X=24589 $Y=22852 $D=636
M2542 1268 327 315 vdd hvtpfet l=6e-08 w=4.11e-07 $X=24589 $Y=27509 $D=636
M2543 1269 clka 324 vdd hvtpfet l=6e-08 w=4.8e-07 $X=24780 $Y=29394 $D=636
M2544 1270 clka 298 vdd hvtpfet l=6e-08 w=4.8e-07 $X=24780 $Y=33942 $D=636
M2545 b_pxca_n<6> 335 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=24830 $Y=1941 $D=636
M2546 335 336 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=24830 $Y=5141 $D=636
M2547 336 337 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=24830 $Y=8691 $D=636
M2548 338 337 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=24830 $Y=41842 $D=636
M2549 339 338 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=24830 $Y=44992 $D=636
M2550 t_pxca_n<6> 339 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=24830 $Y=46622 $D=636
M2551 1271 tm<8> vdd vdd hvtpfet l=6e-08 w=4.8e-07 $X=24853 $Y=10476 $D=636
M2552 vdd 317 1265 vdd hvtpfet l=6e-08 w=8.23e-07 $X=24859 $Y=15520 $D=636
M2553 vdd 317 1266 vdd hvtpfet l=6e-08 w=8.23e-07 $X=24859 $Y=20589 $D=636
M2554 vdd 317 1267 vdd hvtpfet l=6e-08 w=8.23e-07 $X=24859 $Y=22440 $D=636
M2555 vdd 317 1268 vdd hvtpfet l=6e-08 w=8.23e-07 $X=24859 $Y=27509 $D=636
M2556 1272 264 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=24874 $Y=35907 $D=636
M2557 vdd aa<1> 329 vdd hvtpfet l=6e-08 w=4.11e-07 $X=24884 $Y=14280 $D=636
M2558 vdd aa<4> 1269 vdd hvtpfet l=6e-08 w=4.8e-07 $X=25040 $Y=29394 $D=636
M2559 vdd wena 1270 vdd hvtpfet l=6e-08 w=4.8e-07 $X=25040 $Y=33942 $D=636
M2560 vdd 335 b_pxca_n<6> vdd hvtpfet l=6e-08 w=2.57e-06 $X=25090 $Y=1941 $D=636
M2561 vdd 336 335 vdd hvtpfet l=6e-08 w=1e-06 $X=25090 $Y=5141 $D=636
M2562 vdd 337 336 vdd hvtpfet l=6e-08 w=6e-07 $X=25090 $Y=8691 $D=636
M2563 vdd 337 338 vdd hvtpfet l=6e-08 w=6e-07 $X=25090 $Y=41842 $D=636
M2564 vdd 338 339 vdd hvtpfet l=6e-08 w=1e-06 $X=25090 $Y=44992 $D=636
M2565 vdd 339 t_pxca_n<6> vdd hvtpfet l=6e-08 w=2.57e-06 $X=25090 $Y=46622 $D=636
M2566 718 tm<9> 1271 vdd hvtpfet l=6e-08 w=4.8e-07 $X=25113 $Y=10476 $D=636
M2567 376 wena 1272 vdd hvtpfet l=6e-08 w=8e-07 $X=25134 $Y=35907 $D=636
M2568 328 329 vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=25394 $Y=14280 $D=636
M2569 b_pxca_n<5> 345 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=25600 $Y=1941 $D=636
M2570 345 346 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=25600 $Y=5141 $D=636
M2571 346 347 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=25600 $Y=8691 $D=636
M2572 348 347 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=25600 $Y=41842 $D=636
M2573 349 348 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=25600 $Y=44992 $D=636
M2574 t_pxca_n<5> 349 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=25600 $Y=46622 $D=636
M2575 337 352 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=25609 $Y=15321 $D=636
M2576 1273 337 vdd vdd hvtpfet l=6e-08 w=2.74e-07 $X=25609 $Y=16069 $D=636
M2577 1274 320 vdd vdd hvtpfet l=6e-08 w=2.74e-07 $X=25609 $Y=20589 $D=636
M2578 320 353 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=25609 $Y=21405 $D=636
M2579 350 354 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=25609 $Y=22241 $D=636
M2580 1275 350 vdd vdd hvtpfet l=6e-08 w=2.74e-07 $X=25609 $Y=22989 $D=636
M2581 1276 351 vdd vdd hvtpfet l=6e-08 w=2.74e-07 $X=25609 $Y=27509 $D=636
M2582 351 355 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=25609 $Y=28325 $D=636
M2583 1277 tm<9> 721 vdd hvtpfet l=6e-08 w=4.8e-07 $X=25623 $Y=10476 $D=636
M2584 vdd clka 340 vdd hvtpfet l=6e-08 w=9e-07 $X=25854 $Y=29274 $D=636
M2585 vdd 345 b_pxca_n<5> vdd hvtpfet l=6e-08 w=2.57e-06 $X=25860 $Y=1941 $D=636
M2586 vdd 346 345 vdd hvtpfet l=6e-08 w=1e-06 $X=25860 $Y=5141 $D=636
M2587 vdd 347 346 vdd hvtpfet l=6e-08 w=6e-07 $X=25860 $Y=8691 $D=636
M2588 vdd 347 348 vdd hvtpfet l=6e-08 w=6e-07 $X=25860 $Y=41842 $D=636
M2589 vdd 348 349 vdd hvtpfet l=6e-08 w=1e-06 $X=25860 $Y=44992 $D=636
M2590 vdd 349 t_pxca_n<5> vdd hvtpfet l=6e-08 w=2.57e-06 $X=25860 $Y=46622 $D=636
M2591 vdd 352 337 vdd hvtpfet l=6e-08 w=2.06e-07 $X=25869 $Y=15321 $D=636
M2592 352 323 1273 vdd hvtpfet l=6e-08 w=2.74e-07 $X=25869 $Y=16069 $D=636
M2593 353 323 1274 vdd hvtpfet l=6e-08 w=2.74e-07 $X=25869 $Y=20589 $D=636
M2594 vdd 353 320 vdd hvtpfet l=6e-08 w=2.06e-07 $X=25869 $Y=21405 $D=636
M2595 vdd 354 350 vdd hvtpfet l=6e-08 w=2.06e-07 $X=25869 $Y=22241 $D=636
M2596 354 323 1275 vdd hvtpfet l=6e-08 w=2.74e-07 $X=25869 $Y=22989 $D=636
M2597 355 323 1276 vdd hvtpfet l=6e-08 w=2.74e-07 $X=25869 $Y=27509 $D=636
M2598 vdd 355 351 vdd hvtpfet l=6e-08 w=2.06e-07 $X=25869 $Y=28325 $D=636
M2599 vdd 366 1277 vdd hvtpfet l=6e-08 w=4.8e-07 $X=25883 $Y=10476 $D=636
M2600 vdd 356 363 vdd hvtpfet l=6e-08 w=3.2e-07 $X=26138 $Y=35913 $D=636
M2601 b_pxca_n<4> 357 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=26370 $Y=1941 $D=636
M2602 357 358 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=26370 $Y=5141 $D=636
M2603 358 359 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=26370 $Y=8691 $D=636
M2604 360 359 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=26370 $Y=41842 $D=636
M2605 361 360 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=26370 $Y=44992 $D=636
M2606 t_pxca_n<4> 361 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=26370 $Y=46622 $D=636
M2607 729 123 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=26374 $Y=29274 $D=636
M2608 1279 317 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=26379 $Y=15520 $D=636
M2609 1280 317 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=26379 $Y=20589 $D=636
M2610 1281 317 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=26379 $Y=22440 $D=636
M2611 1282 317 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=26379 $Y=27509 $D=636
M2612 1278 366 vdd vdd hvtpfet l=6e-08 w=4.8e-07 $X=26393 $Y=10476 $D=636
M2613 725 368 vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=26398 $Y=35913 $D=636
M2614 vdd 357 b_pxca_n<4> vdd hvtpfet l=6e-08 w=2.57e-06 $X=26630 $Y=1941 $D=636
M2615 vdd 358 357 vdd hvtpfet l=6e-08 w=1e-06 $X=26630 $Y=5141 $D=636
M2616 vdd 359 358 vdd hvtpfet l=6e-08 w=6e-07 $X=26630 $Y=8691 $D=636
M2617 vdd 359 360 vdd hvtpfet l=6e-08 w=6e-07 $X=26630 $Y=41842 $D=636
M2618 vdd 360 361 vdd hvtpfet l=6e-08 w=1e-06 $X=26630 $Y=44992 $D=636
M2619 vdd 361 t_pxca_n<4> vdd hvtpfet l=6e-08 w=2.57e-06 $X=26630 $Y=46622 $D=636
M2620 vdd 123 729 vdd hvtpfet l=6e-08 w=6e-07 $X=26634 $Y=29274 $D=636
M2621 352 364 1279 vdd hvtpfet l=6e-08 w=4.11e-07 $X=26649 $Y=15932 $D=636
M2622 353 364 1280 vdd hvtpfet l=6e-08 w=4.11e-07 $X=26649 $Y=20589 $D=636
M2623 354 365 1281 vdd hvtpfet l=6e-08 w=4.11e-07 $X=26649 $Y=22852 $D=636
M2624 355 365 1282 vdd hvtpfet l=6e-08 w=4.11e-07 $X=26649 $Y=27509 $D=636
M2625 727 325 1278 vdd hvtpfet l=6e-08 w=4.8e-07 $X=26653 $Y=10476 $D=636
M2626 356 363 725 vdd hvtpfet l=6e-08 w=3.2e-07 $X=26658 $Y=35913 $D=636
M2627 vdd tm<7> 726 vdd hvtpfet l=6e-08 w=4.11e-07 $X=26820 $Y=40177 $D=636
M2628 1283 123 vdd vdd hvtpfet l=6e-08 w=4.8e-07 $X=26839 $Y=33942 $D=636
M2629 729 123 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=26894 $Y=29274 $D=636
M2630 1285 369 352 vdd hvtpfet l=6e-08 w=4.11e-07 $X=26909 $Y=15932 $D=636
M2631 1286 369 353 vdd hvtpfet l=6e-08 w=4.11e-07 $X=26909 $Y=20589 $D=636
M2632 1287 369 354 vdd hvtpfet l=6e-08 w=4.11e-07 $X=26909 $Y=22852 $D=636
M2633 1288 369 355 vdd hvtpfet l=6e-08 w=4.11e-07 $X=26909 $Y=27509 $D=636
M2634 1284 362 356 vdd hvtpfet l=6e-08 w=4.8e-07 $X=26918 $Y=35753 $D=636
M2635 vdd aa<10> 374 vdd hvtpfet l=6e-08 w=4.11e-07 $X=26924 $Y=14280 $D=636
M2636 379 131 1283 vdd hvtpfet l=6e-08 w=4.8e-07 $X=27099 $Y=33942 $D=636
M2637 b_pxca_n<3> 370 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=27140 $Y=1941 $D=636
M2638 370 371 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=27140 $Y=5141 $D=636
M2639 371 351 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=27140 $Y=8691 $D=636
M2640 372 351 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=27140 $Y=41842 $D=636
M2641 373 372 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=27140 $Y=44992 $D=636
M2642 t_pxca_n<3> 373 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=27140 $Y=46622 $D=636
M2643 vdd 123 729 vdd hvtpfet l=6e-08 w=6e-07 $X=27154 $Y=29274 $D=636
M2644 vdd tm<9> 325 vdd hvtpfet l=7e-08 w=4.8e-07 $X=27163 $Y=10476 $D=636
M2645 vdd 376 1284 vdd hvtpfet l=6e-08 w=4.8e-07 $X=27178 $Y=35753 $D=636
M2646 vdd 317 1285 vdd hvtpfet l=6e-08 w=8.23e-07 $X=27179 $Y=15520 $D=636
M2647 vdd 317 1286 vdd hvtpfet l=6e-08 w=8.23e-07 $X=27179 $Y=20589 $D=636
M2648 vdd 317 1287 vdd hvtpfet l=6e-08 w=8.23e-07 $X=27179 $Y=22440 $D=636
M2649 vdd 317 1288 vdd hvtpfet l=6e-08 w=8.23e-07 $X=27179 $Y=27509 $D=636
M2650 375 374 vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=27184 $Y=14280 $D=636
M2651 736 377 379 vdd hvtpfet l=6e-08 w=3.2e-07 $X=27359 $Y=33942 $D=636
M2652 vdd 370 b_pxca_n<3> vdd hvtpfet l=6e-08 w=2.57e-06 $X=27400 $Y=1941 $D=636
M2653 vdd 371 370 vdd hvtpfet l=6e-08 w=1e-06 $X=27400 $Y=5141 $D=636
M2654 vdd 351 371 vdd hvtpfet l=6e-08 w=6e-07 $X=27400 $Y=8691 $D=636
M2655 vdd 351 372 vdd hvtpfet l=6e-08 w=6e-07 $X=27400 $Y=41842 $D=636
M2656 vdd 372 373 vdd hvtpfet l=6e-08 w=1e-06 $X=27400 $Y=44992 $D=636
M2657 vdd 373 t_pxca_n<3> vdd hvtpfet l=6e-08 w=2.57e-06 $X=27400 $Y=46622 $D=636
M2658 366 tm<8> vdd vdd hvtpfet l=7e-08 w=4.8e-07 $X=27433 $Y=10476 $D=636
M2659 vdd 123 736 vdd hvtpfet l=6e-08 w=3.2e-07 $X=27619 $Y=33942 $D=636
M2660 vdd tm<1> 735 vdd hvtpfet l=6e-08 w=4.11e-07 $X=27620 $Y=40177 $D=636
M2661 317 323 vdd vdd hvtpfet l=6e-08 w=7e-07 $X=27664 $Y=29648 $D=636
M2662 1289 374 352 vdd hvtpfet l=6e-08 w=4.11e-07 $X=27689 $Y=15932 $D=636
M2663 1290 375 353 vdd hvtpfet l=6e-08 w=4.11e-07 $X=27689 $Y=20589 $D=636
M2664 1291 374 354 vdd hvtpfet l=6e-08 w=4.11e-07 $X=27689 $Y=22852 $D=636
M2665 1292 375 355 vdd hvtpfet l=6e-08 w=4.11e-07 $X=27689 $Y=27509 $D=636
M2666 vdd 380 369 vdd hvtpfet l=6e-08 w=4.11e-07 $X=27784 $Y=14280 $D=636
M2667 vdd 362 386 vdd hvtpfet l=6e-08 w=4e-07 $X=27858 $Y=35682 $D=636
M2668 377 379 vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=27879 $Y=33942 $D=636
M2669 b_pxca_n<2> 381 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=27910 $Y=1941 $D=636
M2670 381 382 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=27910 $Y=5141 $D=636
M2671 382 350 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=27910 $Y=8691 $D=636
M2672 383 350 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=27910 $Y=41842 $D=636
M2673 384 383 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=27910 $Y=44992 $D=636
M2674 t_pxca_n<2> 384 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=27910 $Y=46622 $D=636
M2675 vdd 323 317 vdd hvtpfet l=6e-08 w=7e-07 $X=27924 $Y=29648 $D=636
M2676 vdd 317 1289 vdd hvtpfet l=6e-08 w=8.23e-07 $X=27959 $Y=15520 $D=636
M2677 vdd 317 1290 vdd hvtpfet l=6e-08 w=8.23e-07 $X=27959 $Y=20589 $D=636
M2678 vdd 317 1291 vdd hvtpfet l=6e-08 w=8.23e-07 $X=27959 $Y=22440 $D=636
M2679 vdd 317 1292 vdd hvtpfet l=6e-08 w=8.23e-07 $X=27959 $Y=27509 $D=636
M2680 380 aa<11> vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=28044 $Y=14280 $D=636
M2681 386 356 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=28118 $Y=35682 $D=636
M2682 vdd 381 b_pxca_n<2> vdd hvtpfet l=6e-08 w=2.57e-06 $X=28170 $Y=1941 $D=636
M2683 vdd 382 381 vdd hvtpfet l=6e-08 w=1e-06 $X=28170 $Y=5141 $D=636
M2684 vdd 350 382 vdd hvtpfet l=6e-08 w=6e-07 $X=28170 $Y=8691 $D=636
M2685 vdd 350 383 vdd hvtpfet l=6e-08 w=6e-07 $X=28170 $Y=41842 $D=636
M2686 vdd 383 384 vdd hvtpfet l=6e-08 w=1e-06 $X=28170 $Y=44992 $D=636
M2687 vdd 384 t_pxca_n<2> vdd hvtpfet l=6e-08 w=2.57e-06 $X=28170 $Y=46622 $D=636
M2688 317 323 vdd vdd hvtpfet l=6e-08 w=7e-07 $X=28184 $Y=29648 $D=636
M2689 1293 317 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=28219 $Y=15520 $D=636
M2690 1294 317 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=28219 $Y=20589 $D=636
M2691 1295 317 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=28219 $Y=22440 $D=636
M2692 1296 317 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=28219 $Y=27509 $D=636
M2693 vdd 323 317 vdd hvtpfet l=6e-08 w=7e-07 $X=28444 $Y=29648 $D=636
M2694 407 374 1293 vdd hvtpfet l=6e-08 w=4.11e-07 $X=28489 $Y=15932 $D=636
M2695 408 375 1294 vdd hvtpfet l=6e-08 w=4.11e-07 $X=28489 $Y=20589 $D=636
M2696 409 374 1295 vdd hvtpfet l=6e-08 w=4.11e-07 $X=28489 $Y=22852 $D=636
M2697 410 375 1296 vdd hvtpfet l=6e-08 w=4.11e-07 $X=28489 $Y=27509 $D=636
M2698 vdd 392 541 vdd hvtpfet l=6e-08 w=4e-07 $X=28514 $Y=10167 $D=636
M2699 vdd 393 544 vdd hvtpfet l=6e-08 w=4e-07 $X=28514 $Y=40566 $D=636
M2700 494 386 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=28628 $Y=35682 $D=636
M2701 b_pxca_n<1> 387 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=28680 $Y=1941 $D=636
M2702 387 388 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=28680 $Y=5141 $D=636
M2703 388 389 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=28680 $Y=8691 $D=636
M2704 390 389 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=28680 $Y=41842 $D=636
M2705 391 390 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=28680 $Y=44992 $D=636
M2706 t_pxca_n<1> 391 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=28680 $Y=46622 $D=636
M2707 742 123 vdd vdd hvtpfet l=6e-08 w=1.2e-06 $X=28704 $Y=29148 $D=636
M2708 vdd 387 b_pxca_n<1> vdd hvtpfet l=6e-08 w=2.57e-06 $X=28940 $Y=1941 $D=636
M2709 vdd 388 387 vdd hvtpfet l=6e-08 w=1e-06 $X=28940 $Y=5141 $D=636
M2710 vdd 389 388 vdd hvtpfet l=6e-08 w=6e-07 $X=28940 $Y=8691 $D=636
M2711 vdd 389 390 vdd hvtpfet l=6e-08 w=6e-07 $X=28940 $Y=41842 $D=636
M2712 vdd 390 391 vdd hvtpfet l=6e-08 w=1e-06 $X=28940 $Y=44992 $D=636
M2713 vdd 391 t_pxca_n<1> vdd hvtpfet l=6e-08 w=2.57e-06 $X=28940 $Y=46622 $D=636
M2714 1297 317 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=28999 $Y=15520 $D=636
M2715 1298 317 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=28999 $Y=20589 $D=636
M2716 1299 317 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=28999 $Y=22440 $D=636
M2717 1300 317 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=28999 $Y=27509 $D=636
M2718 vdd 308 392 vdd hvtpfet l=6e-08 w=4.11e-07 $X=29024 $Y=10156 $D=636
M2719 vdd 308 393 vdd hvtpfet l=6e-08 w=4.11e-07 $X=29024 $Y=40566 $D=636
M2720 vdd aa<12> 365 vdd hvtpfet l=6e-08 w=4.11e-07 $X=29054 $Y=14280 $D=636
M2721 407 380 1297 vdd hvtpfet l=6e-08 w=4.11e-07 $X=29269 $Y=15932 $D=636
M2722 408 380 1298 vdd hvtpfet l=6e-08 w=4.11e-07 $X=29269 $Y=20589 $D=636
M2723 409 380 1299 vdd hvtpfet l=6e-08 w=4.11e-07 $X=29269 $Y=22852 $D=636
M2724 410 380 1300 vdd hvtpfet l=6e-08 w=4.11e-07 $X=29269 $Y=27509 $D=636
M2725 392 dwla<1> vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=29284 $Y=10156 $D=636
M2726 393 dwla<0> vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=29284 $Y=40566 $D=636
M2727 743 395 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=29298 $Y=33468 $D=636
M2728 b_pxca_n<0> 396 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=29450 $Y=1941 $D=636
M2729 396 397 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=29450 $Y=5141 $D=636
M2730 397 398 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=29450 $Y=8691 $D=636
M2731 399 398 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=29450 $Y=41842 $D=636
M2732 400 399 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=29450 $Y=44992 $D=636
M2733 t_pxca_n<0> 400 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=29450 $Y=46622 $D=636
M2734 748 403 456 vdd hvtpfet l=6e-08 w=1e-06 $X=29487 $Y=35707 $D=636
M2735 1301 364 407 vdd hvtpfet l=6e-08 w=4.11e-07 $X=29529 $Y=15932 $D=636
M2736 1302 364 408 vdd hvtpfet l=6e-08 w=4.11e-07 $X=29529 $Y=20589 $D=636
M2737 1303 365 409 vdd hvtpfet l=6e-08 w=4.11e-07 $X=29529 $Y=22852 $D=636
M2738 1304 365 410 vdd hvtpfet l=6e-08 w=4.11e-07 $X=29529 $Y=27509 $D=636
M2739 403 405 743 vdd hvtpfet l=6e-08 w=6e-07 $X=29558 $Y=33468 $D=636
M2740 364 365 vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=29564 $Y=14280 $D=636
M2741 vdd 404 395 vdd hvtpfet l=2.5e-07 w=5e-07 $X=29591 $Y=29813 $D=636
M2742 vdd 396 b_pxca_n<0> vdd hvtpfet l=6e-08 w=2.57e-06 $X=29710 $Y=1941 $D=636
M2743 vdd 397 396 vdd hvtpfet l=6e-08 w=1e-06 $X=29710 $Y=5141 $D=636
M2744 vdd 398 397 vdd hvtpfet l=6e-08 w=6e-07 $X=29710 $Y=8691 $D=636
M2745 vdd 398 399 vdd hvtpfet l=6e-08 w=6e-07 $X=29710 $Y=41842 $D=636
M2746 vdd 399 400 vdd hvtpfet l=6e-08 w=1e-06 $X=29710 $Y=44992 $D=636
M2747 vdd 400 t_pxca_n<0> vdd hvtpfet l=6e-08 w=2.57e-06 $X=29710 $Y=46622 $D=636
M2748 456 403 748 vdd hvtpfet l=6e-08 w=1e-06 $X=29747 $Y=35707 $D=636
M2749 vdd 317 1301 vdd hvtpfet l=6e-08 w=8.23e-07 $X=29799 $Y=15520 $D=636
M2750 vdd 317 1302 vdd hvtpfet l=6e-08 w=8.23e-07 $X=29799 $Y=20589 $D=636
M2751 vdd 317 1303 vdd hvtpfet l=6e-08 w=8.23e-07 $X=29799 $Y=22440 $D=636
M2752 vdd 317 1304 vdd hvtpfet l=6e-08 w=8.23e-07 $X=29799 $Y=27509 $D=636
M2753 748 403 456 vdd hvtpfet l=6e-08 w=1e-06 $X=30007 $Y=35707 $D=636
M2754 404 406 vdd vdd hvtpfet l=6e-08 w=5e-07 $X=30041 $Y=29813 $D=636
M2755 405 tm<7> vdd vdd hvtpfet l=6e-08 w=3e-07 $X=30068 $Y=33468 $D=636
M2756 dbl_pd_n<3> 131 vdd vdd hvtpfet l=6e-08 w=4.28e-07 $X=30204 $Y=14263 $D=636
M2757 b_pxba_n<7> 411 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=30220 $Y=1941 $D=636
M2758 411 412 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=30220 $Y=5141 $D=636
M2759 412 413 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=30220 $Y=8691 $D=636
M2760 414 413 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=30220 $Y=41842 $D=636
M2761 415 414 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=30220 $Y=44992 $D=636
M2762 t_pxba_n<7> 415 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=30220 $Y=46622 $D=636
M2763 753 416 748 vdd hvtpfet l=6e-08 w=1e-06 $X=30267 $Y=35707 $D=636
M2764 359 407 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=30309 $Y=15321 $D=636
M2765 1305 323 407 vdd hvtpfet l=6e-08 w=2.74e-07 $X=30309 $Y=16069 $D=636
M2766 1306 323 408 vdd hvtpfet l=6e-08 w=2.74e-07 $X=30309 $Y=20589 $D=636
M2767 347 408 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=30309 $Y=21405 $D=636
M2768 398 409 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=30309 $Y=22241 $D=636
M2769 1307 323 409 vdd hvtpfet l=6e-08 w=2.74e-07 $X=30309 $Y=22989 $D=636
M2770 1308 323 410 vdd hvtpfet l=6e-08 w=2.74e-07 $X=30309 $Y=27509 $D=636
M2771 389 410 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=30309 $Y=28325 $D=636
M2772 vdd 131 dbl_pd_n<3> vdd hvtpfet l=6e-08 w=4.28e-07 $X=30464 $Y=14263 $D=636
M2773 vdd 411 b_pxba_n<7> vdd hvtpfet l=6e-08 w=2.57e-06 $X=30480 $Y=1941 $D=636
M2774 vdd 412 411 vdd hvtpfet l=6e-08 w=1e-06 $X=30480 $Y=5141 $D=636
M2775 vdd 413 412 vdd hvtpfet l=6e-08 w=6e-07 $X=30480 $Y=8691 $D=636
M2776 vdd 413 414 vdd hvtpfet l=6e-08 w=6e-07 $X=30480 $Y=41842 $D=636
M2777 vdd 414 415 vdd hvtpfet l=6e-08 w=1e-06 $X=30480 $Y=44992 $D=636
M2778 vdd 415 t_pxba_n<7> vdd hvtpfet l=6e-08 w=2.57e-06 $X=30480 $Y=46622 $D=636
M2779 748 416 753 vdd hvtpfet l=6e-08 w=1e-06 $X=30527 $Y=35707 $D=636
M2780 vdd 407 359 vdd hvtpfet l=6e-08 w=2.06e-07 $X=30569 $Y=15321 $D=636
M2781 vdd 359 1305 vdd hvtpfet l=6e-08 w=2.74e-07 $X=30569 $Y=16069 $D=636
M2782 vdd 347 1306 vdd hvtpfet l=6e-08 w=2.74e-07 $X=30569 $Y=20589 $D=636
M2783 vdd 408 347 vdd hvtpfet l=6e-08 w=2.06e-07 $X=30569 $Y=21405 $D=636
M2784 vdd 409 398 vdd hvtpfet l=6e-08 w=2.06e-07 $X=30569 $Y=22241 $D=636
M2785 vdd 398 1307 vdd hvtpfet l=6e-08 w=2.74e-07 $X=30569 $Y=22989 $D=636
M2786 vdd 389 1308 vdd hvtpfet l=6e-08 w=2.74e-07 $X=30569 $Y=27509 $D=636
M2787 vdd 410 389 vdd hvtpfet l=6e-08 w=2.06e-07 $X=30569 $Y=28325 $D=636
M2788 vdd dwla<1> 426 vdd hvtpfet l=6e-08 w=4.11e-07 $X=30584 $Y=10156 $D=636
M2789 vdd dwla<0> 427 vdd hvtpfet l=6e-08 w=4.11e-07 $X=30584 $Y=40566 $D=636
M2790 749 406 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=30644 $Y=33468 $D=636
M2791 vdd 417 406 vdd hvtpfet l=2.5e-07 w=5e-07 $X=30711 $Y=29813 $D=636
M2792 dbl_pd_n<3> 131 vdd vdd hvtpfet l=6e-08 w=4.28e-07 $X=30724 $Y=14263 $D=636
M2793 753 416 748 vdd hvtpfet l=6e-08 w=1e-06 $X=30787 $Y=35707 $D=636
M2794 426 309 vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=30844 $Y=10156 $D=636
M2795 427 309 vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=30844 $Y=40566 $D=636
M2796 416 423 749 vdd hvtpfet l=6e-08 w=6e-07 $X=30904 $Y=33468 $D=636
M2797 b_pxba_n<6> 418 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=30990 $Y=1941 $D=636
M2798 418 419 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=30990 $Y=5141 $D=636
M2799 419 420 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=30990 $Y=8691 $D=636
M2800 421 420 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=30990 $Y=41842 $D=636
M2801 422 421 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=30990 $Y=44992 $D=636
M2802 t_pxba_n<6> 422 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=30990 $Y=46622 $D=636
M2803 vdd 362 753 vdd hvtpfet l=6e-08 w=1e-06 $X=31047 $Y=35707 $D=636
M2804 420 428 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=31079 $Y=15321 $D=636
M2805 1309 420 vdd vdd hvtpfet l=6e-08 w=2.74e-07 $X=31079 $Y=16069 $D=636
M2806 1310 413 vdd vdd hvtpfet l=6e-08 w=2.74e-07 $X=31079 $Y=20589 $D=636
M2807 413 429 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=31079 $Y=21405 $D=636
M2808 424 430 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=31079 $Y=22241 $D=636
M2809 1311 424 vdd vdd hvtpfet l=6e-08 w=2.74e-07 $X=31079 $Y=22989 $D=636
M2810 1312 425 vdd vdd hvtpfet l=6e-08 w=2.74e-07 $X=31079 $Y=27509 $D=636
M2811 425 431 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=31079 $Y=28325 $D=636
M2812 417 368 vdd vdd hvtpfet l=6e-08 w=5e-07 $X=31161 $Y=29813 $D=636
M2813 dbl_pd_n<1> tm<1> vdd vdd hvtpfet l=6e-08 w=4.28e-07 $X=31234 $Y=14263 $D=636
M2814 vdd 418 b_pxba_n<6> vdd hvtpfet l=6e-08 w=2.57e-06 $X=31250 $Y=1941 $D=636
M2815 vdd 419 418 vdd hvtpfet l=6e-08 w=1e-06 $X=31250 $Y=5141 $D=636
M2816 vdd 420 419 vdd hvtpfet l=6e-08 w=6e-07 $X=31250 $Y=8691 $D=636
M2817 vdd 420 421 vdd hvtpfet l=6e-08 w=6e-07 $X=31250 $Y=41842 $D=636
M2818 vdd 421 422 vdd hvtpfet l=6e-08 w=1e-06 $X=31250 $Y=44992 $D=636
M2819 vdd 422 t_pxba_n<6> vdd hvtpfet l=6e-08 w=2.57e-06 $X=31250 $Y=46622 $D=636
M2820 753 362 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=31307 $Y=35707 $D=636
M2821 vdd 428 420 vdd hvtpfet l=6e-08 w=2.06e-07 $X=31339 $Y=15321 $D=636
M2822 428 323 1309 vdd hvtpfet l=6e-08 w=2.74e-07 $X=31339 $Y=16069 $D=636
M2823 429 323 1310 vdd hvtpfet l=6e-08 w=2.74e-07 $X=31339 $Y=20589 $D=636
M2824 vdd 429 413 vdd hvtpfet l=6e-08 w=2.06e-07 $X=31339 $Y=21405 $D=636
M2825 vdd 430 424 vdd hvtpfet l=6e-08 w=2.06e-07 $X=31339 $Y=22241 $D=636
M2826 430 323 1311 vdd hvtpfet l=6e-08 w=2.74e-07 $X=31339 $Y=22989 $D=636
M2827 431 323 1312 vdd hvtpfet l=6e-08 w=2.74e-07 $X=31339 $Y=27509 $D=636
M2828 vdd 431 425 vdd hvtpfet l=6e-08 w=2.06e-07 $X=31339 $Y=28325 $D=636
M2829 556 426 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=31354 $Y=10167 $D=636
M2830 558 427 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=31354 $Y=40566 $D=636
M2831 vdd 173 423 vdd hvtpfet l=6e-08 w=3e-07 $X=31414 $Y=33468 $D=636
M2832 vdd tm<1> dbl_pd_n<1> vdd hvtpfet l=6e-08 w=4.28e-07 $X=31494 $Y=14263 $D=636
M2833 vdd 362 753 vdd hvtpfet l=6e-08 w=1e-06 $X=31567 $Y=35707 $D=636
M2834 dbl_pd_n<1> tm<1> vdd vdd hvtpfet l=6e-08 w=4.28e-07 $X=31754 $Y=14263 $D=636
M2835 b_pxba_n<5> 432 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=31760 $Y=1941 $D=636
M2836 432 433 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=31760 $Y=5141 $D=636
M2837 433 434 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=31760 $Y=8691 $D=636
M2838 435 434 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=31760 $Y=41842 $D=636
M2839 436 435 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=31760 $Y=44992 $D=636
M2840 t_pxba_n<5> 436 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=31760 $Y=46622 $D=636
M2841 vdd 368 362 vdd hvtpfet l=6e-08 w=4e-07 $X=31761 $Y=29948 $D=636
M2842 1313 317 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=31849 $Y=15520 $D=636
M2843 1314 317 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=31849 $Y=20589 $D=636
M2844 1315 317 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=31849 $Y=22440 $D=636
M2845 1316 317 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=31849 $Y=27509 $D=636
M2846 vdd 437 540 vdd hvtpfet l=6e-08 w=4e-07 $X=31864 $Y=10167 $D=636
M2847 vdd 438 545 vdd hvtpfet l=6e-08 w=4e-07 $X=31864 $Y=40566 $D=636
M2848 vdd 432 b_pxba_n<5> vdd hvtpfet l=6e-08 w=2.57e-06 $X=32020 $Y=1941 $D=636
M2849 vdd 433 432 vdd hvtpfet l=6e-08 w=1e-06 $X=32020 $Y=5141 $D=636
M2850 vdd 434 433 vdd hvtpfet l=6e-08 w=6e-07 $X=32020 $Y=8691 $D=636
M2851 vdd 434 435 vdd hvtpfet l=6e-08 w=6e-07 $X=32020 $Y=41842 $D=636
M2852 vdd 435 436 vdd hvtpfet l=6e-08 w=1e-06 $X=32020 $Y=44992 $D=636
M2853 vdd 436 t_pxba_n<5> vdd hvtpfet l=6e-08 w=2.57e-06 $X=32020 $Y=46622 $D=636
M2854 428 439 1313 vdd hvtpfet l=6e-08 w=4.11e-07 $X=32119 $Y=15932 $D=636
M2855 429 439 1314 vdd hvtpfet l=6e-08 w=4.11e-07 $X=32119 $Y=20589 $D=636
M2856 430 440 1315 vdd hvtpfet l=6e-08 w=4.11e-07 $X=32119 $Y=22852 $D=636
M2857 431 440 1316 vdd hvtpfet l=6e-08 w=4.11e-07 $X=32119 $Y=27509 $D=636
M2858 761 442 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=32271 $Y=29348 $D=636
M2859 762 442 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=32271 $Y=35707 $D=636
M2860 vdd 310 437 vdd hvtpfet l=6e-08 w=4.11e-07 $X=32374 $Y=10156 $D=636
M2861 vdd 310 438 vdd hvtpfet l=6e-08 w=4.11e-07 $X=32374 $Y=40566 $D=636
M2862 1317 443 428 vdd hvtpfet l=6e-08 w=4.11e-07 $X=32379 $Y=15932 $D=636
M2863 1318 443 429 vdd hvtpfet l=6e-08 w=4.11e-07 $X=32379 $Y=20589 $D=636
M2864 1319 443 430 vdd hvtpfet l=6e-08 w=4.11e-07 $X=32379 $Y=22852 $D=636
M2865 1320 443 431 vdd hvtpfet l=6e-08 w=4.11e-07 $X=32379 $Y=27509 $D=636
M2866 vdd aa<7> 449 vdd hvtpfet l=6e-08 w=4.11e-07 $X=32394 $Y=14280 $D=636
M2867 vdd 324 442 vdd hvtpfet l=6e-08 w=1e-06 $X=32394 $Y=33493 $D=636
M2868 b_pxba_n<4> 444 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=32530 $Y=1941 $D=636
M2869 444 445 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=32530 $Y=5141 $D=636
M2870 445 446 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=32530 $Y=8691 $D=636
M2871 447 446 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=32530 $Y=41842 $D=636
M2872 448 447 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=32530 $Y=44992 $D=636
M2873 t_pxba_n<4> 448 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=32530 $Y=46622 $D=636
M2874 vdd 442 761 vdd hvtpfet l=6e-08 w=1e-06 $X=32531 $Y=29348 $D=636
M2875 vdd 442 762 vdd hvtpfet l=6e-08 w=1e-06 $X=32531 $Y=35707 $D=636
M2876 437 dwla<1> vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=32634 $Y=10156 $D=636
M2877 438 dwla<0> vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=32634 $Y=40566 $D=636
M2878 vdd 317 1317 vdd hvtpfet l=6e-08 w=8.23e-07 $X=32649 $Y=15520 $D=636
M2879 vdd 317 1318 vdd hvtpfet l=6e-08 w=8.23e-07 $X=32649 $Y=20589 $D=636
M2880 vdd 317 1319 vdd hvtpfet l=6e-08 w=8.23e-07 $X=32649 $Y=22440 $D=636
M2881 vdd 317 1320 vdd hvtpfet l=6e-08 w=8.23e-07 $X=32649 $Y=27509 $D=636
M2882 450 449 vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=32654 $Y=14280 $D=636
M2883 vdd 444 b_pxba_n<4> vdd hvtpfet l=6e-08 w=2.57e-06 $X=32790 $Y=1941 $D=636
M2884 vdd 445 444 vdd hvtpfet l=6e-08 w=1e-06 $X=32790 $Y=5141 $D=636
M2885 vdd 446 445 vdd hvtpfet l=6e-08 w=6e-07 $X=32790 $Y=8691 $D=636
M2886 vdd 446 447 vdd hvtpfet l=6e-08 w=6e-07 $X=32790 $Y=41842 $D=636
M2887 vdd 447 448 vdd hvtpfet l=6e-08 w=1e-06 $X=32790 $Y=44992 $D=636
M2888 vdd 448 t_pxba_n<4> vdd hvtpfet l=6e-08 w=2.57e-06 $X=32790 $Y=46622 $D=636
M2889 dwla<1> 368 761 vdd hvtpfet l=6e-08 w=1e-06 $X=33041 $Y=29348 $D=636
M2890 497 456 762 vdd hvtpfet l=6e-08 w=1e-06 $X=33041 $Y=35707 $D=636
M2891 465 442 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=33094 $Y=33493 $D=636
M2892 vdd dwla<1> 458 vdd hvtpfet l=6e-08 w=4.11e-07 $X=33144 $Y=10156 $D=636
M2893 vdd dwla<0> 459 vdd hvtpfet l=6e-08 w=4.11e-07 $X=33144 $Y=40566 $D=636
M2894 1321 449 428 vdd hvtpfet l=6e-08 w=4.11e-07 $X=33159 $Y=15932 $D=636
M2895 1322 450 429 vdd hvtpfet l=6e-08 w=4.11e-07 $X=33159 $Y=20589 $D=636
M2896 1323 449 430 vdd hvtpfet l=6e-08 w=4.11e-07 $X=33159 $Y=22852 $D=636
M2897 1324 450 431 vdd hvtpfet l=6e-08 w=4.11e-07 $X=33159 $Y=27509 $D=636
M2898 vdd 455 443 vdd hvtpfet l=6e-08 w=4.11e-07 $X=33254 $Y=14280 $D=636
M2899 b_pxba_n<3> 451 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=33300 $Y=1941 $D=636
M2900 451 452 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=33300 $Y=5141 $D=636
M2901 452 425 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=33300 $Y=8691 $D=636
M2902 453 425 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=33300 $Y=41842 $D=636
M2903 454 453 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=33300 $Y=44992 $D=636
M2904 t_pxba_n<3> 454 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=33300 $Y=46622 $D=636
M2905 761 368 dwla<1> vdd hvtpfet l=6e-08 w=1e-06 $X=33301 $Y=29348 $D=636
M2906 762 456 497 vdd hvtpfet l=6e-08 w=1e-06 $X=33301 $Y=35707 $D=636
M2907 458 311 vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=33404 $Y=10156 $D=636
M2908 459 311 vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=33404 $Y=40566 $D=636
M2909 vdd 317 1321 vdd hvtpfet l=6e-08 w=8.23e-07 $X=33429 $Y=15520 $D=636
M2910 vdd 317 1322 vdd hvtpfet l=6e-08 w=8.23e-07 $X=33429 $Y=20589 $D=636
M2911 vdd 317 1323 vdd hvtpfet l=6e-08 w=8.23e-07 $X=33429 $Y=22440 $D=636
M2912 vdd 317 1324 vdd hvtpfet l=6e-08 w=8.23e-07 $X=33429 $Y=27509 $D=636
M2913 455 aa<8> vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=33514 $Y=14280 $D=636
M2914 vdd 451 b_pxba_n<3> vdd hvtpfet l=6e-08 w=2.57e-06 $X=33560 $Y=1941 $D=636
M2915 vdd 452 451 vdd hvtpfet l=6e-08 w=1e-06 $X=33560 $Y=5141 $D=636
M2916 vdd 425 452 vdd hvtpfet l=6e-08 w=6e-07 $X=33560 $Y=8691 $D=636
M2917 vdd 425 453 vdd hvtpfet l=6e-08 w=6e-07 $X=33560 $Y=41842 $D=636
M2918 vdd 453 454 vdd hvtpfet l=6e-08 w=1e-06 $X=33560 $Y=44992 $D=636
M2919 vdd 454 t_pxba_n<3> vdd hvtpfet l=6e-08 w=2.57e-06 $X=33560 $Y=46622 $D=636
M2920 1325 317 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=33689 $Y=15520 $D=636
M2921 1326 317 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=33689 $Y=20589 $D=636
M2922 1327 317 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=33689 $Y=22440 $D=636
M2923 1328 317 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=33689 $Y=27509 $D=636
M2924 dwla<0> 368 765 vdd hvtpfet l=6e-08 w=1e-06 $X=33811 $Y=29348 $D=636
M2925 498 456 766 vdd hvtpfet l=6e-08 w=1e-06 $X=33811 $Y=35707 $D=636
M2926 555 458 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=33914 $Y=10167 $D=636
M2927 559 459 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=33914 $Y=40566 $D=636
M2928 479 449 1325 vdd hvtpfet l=6e-08 w=4.11e-07 $X=33959 $Y=15932 $D=636
M2929 480 450 1326 vdd hvtpfet l=6e-08 w=4.11e-07 $X=33959 $Y=20589 $D=636
M2930 481 449 1327 vdd hvtpfet l=6e-08 w=4.11e-07 $X=33959 $Y=22852 $D=636
M2931 482 450 1328 vdd hvtpfet l=6e-08 w=4.11e-07 $X=33959 $Y=27509 $D=636
M2932 b_pxba_n<2> 460 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=34070 $Y=1941 $D=636
M2933 460 461 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=34070 $Y=5141 $D=636
M2934 461 424 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=34070 $Y=8691 $D=636
M2935 462 424 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=34070 $Y=41842 $D=636
M2936 463 462 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=34070 $Y=44992 $D=636
M2937 t_pxba_n<2> 463 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=34070 $Y=46622 $D=636
M2938 765 368 dwla<0> vdd hvtpfet l=6e-08 w=1e-06 $X=34071 $Y=29348 $D=636
M2939 766 456 498 vdd hvtpfet l=6e-08 w=1e-06 $X=34071 $Y=35707 $D=636
M2940 vdd 460 b_pxba_n<2> vdd hvtpfet l=6e-08 w=2.57e-06 $X=34330 $Y=1941 $D=636
M2941 vdd 461 460 vdd hvtpfet l=6e-08 w=1e-06 $X=34330 $Y=5141 $D=636
M2942 vdd 424 461 vdd hvtpfet l=6e-08 w=6e-07 $X=34330 $Y=8691 $D=636
M2943 vdd 424 462 vdd hvtpfet l=6e-08 w=6e-07 $X=34330 $Y=41842 $D=636
M2944 vdd 462 463 vdd hvtpfet l=6e-08 w=1e-06 $X=34330 $Y=44992 $D=636
M2945 vdd 463 t_pxba_n<2> vdd hvtpfet l=6e-08 w=2.57e-06 $X=34330 $Y=46622 $D=636
M2946 1329 317 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=34469 $Y=15520 $D=636
M2947 1330 317 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=34469 $Y=20589 $D=636
M2948 1331 317 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=34469 $Y=22440 $D=636
M2949 1332 317 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=34469 $Y=27509 $D=636
M2950 vdd aa<9> 440 vdd hvtpfet l=6e-08 w=4.11e-07 $X=34524 $Y=14280 $D=636
M2951 765 465 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=34581 $Y=29348 $D=636
M2952 766 465 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=34581 $Y=35707 $D=636
M2953 vdd vdd 535 vdd hvtpfet l=6e-08 w=6.4e-07 $X=34621 $Y=33468 $D=636
M2954 479 455 1329 vdd hvtpfet l=6e-08 w=4.11e-07 $X=34739 $Y=15932 $D=636
M2955 480 455 1330 vdd hvtpfet l=6e-08 w=4.11e-07 $X=34739 $Y=20589 $D=636
M2956 481 455 1331 vdd hvtpfet l=6e-08 w=4.11e-07 $X=34739 $Y=22852 $D=636
M2957 482 455 1332 vdd hvtpfet l=6e-08 w=4.11e-07 $X=34739 $Y=27509 $D=636
M2958 b_pxba_n<1> 466 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=34840 $Y=1941 $D=636
M2959 466 467 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=34840 $Y=5141 $D=636
M2960 467 468 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=34840 $Y=8691 $D=636
M2961 469 468 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=34840 $Y=41842 $D=636
M2962 470 469 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=34840 $Y=44992 $D=636
M2963 t_pxba_n<1> 470 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=34840 $Y=46622 $D=636
M2964 vdd 465 765 vdd hvtpfet l=6e-08 w=1e-06 $X=34841 $Y=29348 $D=636
M2965 vdd 465 766 vdd hvtpfet l=6e-08 w=1e-06 $X=34841 $Y=35707 $D=636
M2966 535 471 vdd vdd hvtpfet l=6e-08 w=6.4e-07 $X=34881 $Y=33468 $D=636
M2967 vdd 123 131 vdd hvtpfet l=6e-08 w=2e-07 $X=34906 $Y=10756 $D=636
M2968 1333 439 479 vdd hvtpfet l=6e-08 w=4.11e-07 $X=34999 $Y=15932 $D=636
M2969 1334 439 480 vdd hvtpfet l=6e-08 w=4.11e-07 $X=34999 $Y=20589 $D=636
M2970 1335 440 481 vdd hvtpfet l=6e-08 w=4.11e-07 $X=34999 $Y=22852 $D=636
M2971 1336 440 482 vdd hvtpfet l=6e-08 w=4.11e-07 $X=34999 $Y=27509 $D=636
M2972 439 440 vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=35034 $Y=14280 $D=636
M2973 vdd 466 b_pxba_n<1> vdd hvtpfet l=6e-08 w=2.57e-06 $X=35100 $Y=1941 $D=636
M2974 vdd 467 466 vdd hvtpfet l=6e-08 w=1e-06 $X=35100 $Y=5141 $D=636
M2975 vdd 468 467 vdd hvtpfet l=6e-08 w=6e-07 $X=35100 $Y=8691 $D=636
M2976 vdd 468 469 vdd hvtpfet l=6e-08 w=6e-07 $X=35100 $Y=41842 $D=636
M2977 vdd 469 470 vdd hvtpfet l=6e-08 w=1e-06 $X=35100 $Y=44992 $D=636
M2978 vdd 470 t_pxba_n<1> vdd hvtpfet l=6e-08 w=2.57e-06 $X=35100 $Y=46622 $D=636
M2979 vdd 317 1333 vdd hvtpfet l=6e-08 w=8.23e-07 $X=35269 $Y=15520 $D=636
M2980 vdd 317 1334 vdd hvtpfet l=6e-08 w=8.23e-07 $X=35269 $Y=20589 $D=636
M2981 vdd 317 1335 vdd hvtpfet l=6e-08 w=8.23e-07 $X=35269 $Y=22440 $D=636
M2982 vdd 317 1336 vdd hvtpfet l=6e-08 w=8.23e-07 $X=35269 $Y=27509 $D=636
M2983 vdd 473 484 vdd hvtpfet l=6e-08 w=3e-07 $X=35351 $Y=36377 $D=636
M2984 vdd 472 471 vdd hvtpfet l=2.5e-07 w=5e-07 $X=35416 $Y=33503 $D=636
M2985 b_pxba_n<0> 474 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=35610 $Y=1941 $D=636
M2986 474 475 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=35610 $Y=5141 $D=636
M2987 475 476 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=35610 $Y=8691 $D=636
M2988 477 476 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=35610 $Y=41842 $D=636
M2989 478 477 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=35610 $Y=44992 $D=636
M2990 t_pxba_n<0> 478 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=35610 $Y=46622 $D=636
M2991 446 479 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=35779 $Y=15321 $D=636
M2992 1337 323 479 vdd hvtpfet l=6e-08 w=2.74e-07 $X=35779 $Y=16069 $D=636
M2993 1338 323 480 vdd hvtpfet l=6e-08 w=2.74e-07 $X=35779 $Y=20589 $D=636
M2994 434 480 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=35779 $Y=21405 $D=636
M2995 476 481 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=35779 $Y=22241 $D=636
M2996 1339 323 481 vdd hvtpfet l=6e-08 w=2.74e-07 $X=35779 $Y=22989 $D=636
M2997 1340 323 482 vdd hvtpfet l=6e-08 w=2.74e-07 $X=35779 $Y=27509 $D=636
M2998 468 482 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=35779 $Y=28325 $D=636
M2999 473 484 vdd vdd hvtpfet l=1.2e-07 w=3e-07 $X=35861 $Y=36382 $D=636
M3000 472 483 vdd vdd hvtpfet l=6e-08 w=5e-07 $X=35866 $Y=33503 $D=636
M3001 vdd 474 b_pxba_n<0> vdd hvtpfet l=6e-08 w=2.57e-06 $X=35870 $Y=1941 $D=636
M3002 vdd 475 474 vdd hvtpfet l=6e-08 w=1e-06 $X=35870 $Y=5141 $D=636
M3003 vdd 476 475 vdd hvtpfet l=6e-08 w=6e-07 $X=35870 $Y=8691 $D=636
M3004 vdd 476 477 vdd hvtpfet l=6e-08 w=6e-07 $X=35870 $Y=41842 $D=636
M3005 vdd 477 478 vdd hvtpfet l=6e-08 w=1e-06 $X=35870 $Y=44992 $D=636
M3006 vdd 478 t_pxba_n<0> vdd hvtpfet l=6e-08 w=2.57e-06 $X=35870 $Y=46622 $D=636
M3007 368 495 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=35945 $Y=29548 $D=636
M3008 vdd 479 446 vdd hvtpfet l=6e-08 w=2.06e-07 $X=36039 $Y=15321 $D=636
M3009 vdd 446 1337 vdd hvtpfet l=6e-08 w=2.74e-07 $X=36039 $Y=16069 $D=636
M3010 vdd 434 1338 vdd hvtpfet l=6e-08 w=2.74e-07 $X=36039 $Y=20589 $D=636
M3011 vdd 480 434 vdd hvtpfet l=6e-08 w=2.06e-07 $X=36039 $Y=21405 $D=636
M3012 vdd 481 476 vdd hvtpfet l=6e-08 w=2.06e-07 $X=36039 $Y=22241 $D=636
M3013 vdd 476 1339 vdd hvtpfet l=6e-08 w=2.74e-07 $X=36039 $Y=22989 $D=636
M3014 vdd 468 1340 vdd hvtpfet l=6e-08 w=2.74e-07 $X=36039 $Y=27509 $D=636
M3015 vdd 482 468 vdd hvtpfet l=6e-08 w=2.06e-07 $X=36039 $Y=28325 $D=636
M3016 vdd 495 368 vdd hvtpfet l=6e-08 w=8e-07 $X=36205 $Y=29548 $D=636
M3017 vdd 491 509 vdd hvtpfet l=6e-08 w=4.11e-07 $X=36254 $Y=14280 $D=636
M3018 b_pxaa<3> 485 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=36380 $Y=1941 $D=636
M3019 485 486 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=36380 $Y=5141 $D=636
M3020 486 487 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=36380 $Y=8691 $D=636
M3021 vdd 492 487 vdd hvtpfet l=6e-08 w=4.11e-07 $X=36380 $Y=10156 $D=636
M3022 vdd 492 488 vdd hvtpfet l=6e-08 w=4.11e-07 $X=36380 $Y=40566 $D=636
M3023 489 488 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=36380 $Y=41842 $D=636
M3024 490 489 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=36380 $Y=44992 $D=636
M3025 t_pxaa<3> 490 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=36380 $Y=46622 $D=636
M3026 vdd 493 473 vdd hvtpfet l=6e-08 w=6.4e-07 $X=36431 $Y=35802 $D=636
M3027 vdd 496 483 vdd hvtpfet l=6e-08 w=6.4e-07 $X=36466 $Y=33468 $D=636
M3028 vdd 485 b_pxaa<3> vdd hvtpfet l=6e-08 w=2.57e-06 $X=36640 $Y=1941 $D=636
M3029 vdd 486 485 vdd hvtpfet l=6e-08 w=1e-06 $X=36640 $Y=5141 $D=636
M3030 vdd 487 486 vdd hvtpfet l=6e-08 w=6e-07 $X=36640 $Y=8691 $D=636
M3031 487 497 vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=36640 $Y=10156 $D=636
M3032 488 498 vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=36640 $Y=40566 $D=636
M3033 vdd 488 489 vdd hvtpfet l=6e-08 w=6e-07 $X=36640 $Y=41842 $D=636
M3034 vdd 489 490 vdd hvtpfet l=6e-08 w=1e-06 $X=36640 $Y=44992 $D=636
M3035 vdd 490 t_pxaa<3> vdd hvtpfet l=6e-08 w=2.57e-06 $X=36640 $Y=46622 $D=636
M3036 368 clka vdd vdd hvtpfet l=6e-08 w=8e-07 $X=36715 $Y=29548 $D=636
M3037 491 aa<6> vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=36764 $Y=14280 $D=636
M3038 1341 317 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=36789 $Y=15520 $D=636
M3039 1342 317 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=36789 $Y=20589 $D=636
M3040 1343 317 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=36789 $Y=22440 $D=636
M3041 1344 317 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=36789 $Y=27509 $D=636
M3042 vdd clka 368 vdd hvtpfet l=6e-08 w=8e-07 $X=36975 $Y=29548 $D=636
M3043 vdd 473 496 vdd hvtpfet l=6e-08 w=6.4e-07 $X=36976 $Y=33693 $D=636
M3044 519 501 1341 vdd hvtpfet l=6e-08 w=4.11e-07 $X=37059 $Y=15932 $D=636
M3045 520 502 1342 vdd hvtpfet l=6e-08 w=4.11e-07 $X=37059 $Y=20589 $D=636
M3046 521 501 1343 vdd hvtpfet l=6e-08 w=4.11e-07 $X=37059 $Y=22852 $D=636
M3047 522 502 1344 vdd hvtpfet l=6e-08 w=4.11e-07 $X=37059 $Y=27509 $D=636
M3048 b_pxaa<2> 503 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=37150 $Y=1941 $D=636
M3049 503 504 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=37150 $Y=5141 $D=636
M3050 504 505 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=37150 $Y=8691 $D=636
M3051 vdd 497 505 vdd hvtpfet l=6e-08 w=4.11e-07 $X=37150 $Y=10156 $D=636
M3052 vdd 498 506 vdd hvtpfet l=6e-08 w=4.11e-07 $X=37150 $Y=40566 $D=636
M3053 507 506 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=37150 $Y=41842 $D=636
M3054 508 507 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=37150 $Y=44992 $D=636
M3055 t_pxaa<2> 508 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=37150 $Y=46622 $D=636
M3056 776 ddqa_n vdd vdd hvtpfet l=6e-08 w=6.4e-07 $X=37161 $Y=35802 $D=636
M3057 vdd 502 501 vdd hvtpfet l=6e-08 w=4.11e-07 $X=37274 $Y=14280 $D=636
M3058 1345 509 519 vdd hvtpfet l=6e-08 w=4.11e-07 $X=37319 $Y=15932 $D=636
M3059 1346 509 520 vdd hvtpfet l=6e-08 w=4.11e-07 $X=37319 $Y=20589 $D=636
M3060 1347 491 521 vdd hvtpfet l=6e-08 w=4.11e-07 $X=37319 $Y=22852 $D=636
M3061 1348 491 522 vdd hvtpfet l=6e-08 w=4.11e-07 $X=37319 $Y=27509 $D=636
M3062 vdd 503 b_pxaa<2> vdd hvtpfet l=6e-08 w=2.57e-06 $X=37410 $Y=1941 $D=636
M3063 vdd 504 503 vdd hvtpfet l=6e-08 w=1e-06 $X=37410 $Y=5141 $D=636
M3064 vdd 505 504 vdd hvtpfet l=6e-08 w=6e-07 $X=37410 $Y=8691 $D=636
M3065 505 510 vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=37410 $Y=10156 $D=636
M3066 506 510 vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=37410 $Y=40566 $D=636
M3067 vdd 506 507 vdd hvtpfet l=6e-08 w=6e-07 $X=37410 $Y=41842 $D=636
M3068 vdd 507 508 vdd hvtpfet l=6e-08 w=1e-06 $X=37410 $Y=44992 $D=636
M3069 vdd 508 t_pxaa<2> vdd hvtpfet l=6e-08 w=2.57e-06 $X=37410 $Y=46622 $D=636
M3070 493 ddqa 776 vdd hvtpfet l=6e-08 w=6.4e-07 $X=37421 $Y=35802 $D=636
M3071 vdd clka 524 vdd hvtpfet l=6e-08 w=1.2e-06 $X=37485 $Y=29148 $D=636
M3072 vdd 317 1345 vdd hvtpfet l=6e-08 w=8.23e-07 $X=37589 $Y=15520 $D=636
M3073 vdd 317 1346 vdd hvtpfet l=6e-08 w=8.23e-07 $X=37589 $Y=20589 $D=636
M3074 vdd 317 1347 vdd hvtpfet l=6e-08 w=8.23e-07 $X=37589 $Y=22440 $D=636
M3075 vdd 317 1348 vdd hvtpfet l=6e-08 w=8.23e-07 $X=37589 $Y=27509 $D=636
M3076 vdd 496 557 vdd hvtpfet l=6e-08 w=6.4e-07 $X=37661 $Y=33693 $D=636
M3077 502 aa<5> vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=37784 $Y=14280 $D=636
M3078 b_pxaa<1> 512 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=37920 $Y=1941 $D=636
M3079 512 513 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=37920 $Y=5141 $D=636
M3080 513 514 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=37920 $Y=8691 $D=636
M3081 vdd 523 514 vdd hvtpfet l=6e-08 w=4.11e-07 $X=37920 $Y=10156 $D=636
M3082 vdd 523 515 vdd hvtpfet l=6e-08 w=4.11e-07 $X=37920 $Y=40566 $D=636
M3083 516 515 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=37920 $Y=41842 $D=636
M3084 517 516 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=37920 $Y=44992 $D=636
M3085 t_pxaa<1> 517 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=37920 $Y=46622 $D=636
M3086 557 386 vdd vdd hvtpfet l=6e-08 w=6.4e-07 $X=37921 $Y=33693 $D=636
M3087 492 519 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=38099 $Y=15321 $D=636
M3088 1349 323 519 vdd hvtpfet l=6e-08 w=2.74e-07 $X=38099 $Y=16069 $D=636
M3089 1350 323 520 vdd hvtpfet l=6e-08 w=2.74e-07 $X=38099 $Y=20589 $D=636
M3090 510 520 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=38099 $Y=21405 $D=636
M3091 523 521 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=38099 $Y=22241 $D=636
M3092 1351 323 521 vdd hvtpfet l=6e-08 w=2.74e-07 $X=38099 $Y=22989 $D=636
M3093 1352 323 522 vdd hvtpfet l=6e-08 w=2.74e-07 $X=38099 $Y=27509 $D=636
M3094 525 522 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=38099 $Y=28325 $D=636
M3095 vdd 493 526 vdd hvtpfet l=1.4e-07 w=6.4e-07 $X=38141 $Y=36067 $D=636
M3096 vdd 512 b_pxaa<1> vdd hvtpfet l=6e-08 w=2.57e-06 $X=38180 $Y=1941 $D=636
M3097 vdd 513 512 vdd hvtpfet l=6e-08 w=1e-06 $X=38180 $Y=5141 $D=636
M3098 vdd 514 513 vdd hvtpfet l=6e-08 w=6e-07 $X=38180 $Y=8691 $D=636
M3099 514 497 vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=38180 $Y=10156 $D=636
M3100 515 498 vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=38180 $Y=40566 $D=636
M3101 vdd 515 516 vdd hvtpfet l=6e-08 w=6e-07 $X=38180 $Y=41842 $D=636
M3102 vdd 516 517 vdd hvtpfet l=6e-08 w=1e-06 $X=38180 $Y=44992 $D=636
M3103 vdd 517 t_pxaa<1> vdd hvtpfet l=6e-08 w=2.57e-06 $X=38180 $Y=46622 $D=636
M3104 1353 524 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=38255 $Y=29525 $D=636
M3105 vdd 519 492 vdd hvtpfet l=6e-08 w=2.06e-07 $X=38359 $Y=15321 $D=636
M3106 vdd 492 1349 vdd hvtpfet l=6e-08 w=2.74e-07 $X=38359 $Y=16069 $D=636
M3107 vdd 510 1350 vdd hvtpfet l=6e-08 w=2.74e-07 $X=38359 $Y=20589 $D=636
M3108 vdd 520 510 vdd hvtpfet l=6e-08 w=2.06e-07 $X=38359 $Y=21405 $D=636
M3109 vdd 521 523 vdd hvtpfet l=6e-08 w=2.06e-07 $X=38359 $Y=22241 $D=636
M3110 vdd 523 1351 vdd hvtpfet l=6e-08 w=2.74e-07 $X=38359 $Y=22989 $D=636
M3111 vdd 525 1352 vdd hvtpfet l=6e-08 w=2.74e-07 $X=38359 $Y=27509 $D=636
M3112 vdd 522 525 vdd hvtpfet l=6e-08 w=2.06e-07 $X=38359 $Y=28325 $D=636
M3113 779 494 vdd vdd hvtpfet l=6e-08 w=6.4e-07 $X=38431 $Y=33468 $D=636
M3114 780 526 vdd vdd hvtpfet l=1.4e-07 w=6.4e-07 $X=38481 $Y=36067 $D=636
M3115 534 495 1353 vdd hvtpfet l=6e-08 w=8.23e-07 $X=38515 $Y=29525 $D=636
M3116 vdd 533 546 vdd hvtpfet l=6e-08 w=4.11e-07 $X=38574 $Y=14280 $D=636
M3117 b_pxaa<0> 527 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=38690 $Y=1941 $D=636
M3118 527 528 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=38690 $Y=5141 $D=636
M3119 528 529 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=38690 $Y=8691 $D=636
M3120 vdd 497 529 vdd hvtpfet l=6e-08 w=4.11e-07 $X=38690 $Y=10156 $D=636
M3121 vdd 498 530 vdd hvtpfet l=6e-08 w=4.11e-07 $X=38690 $Y=40566 $D=636
M3122 531 530 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=38690 $Y=41842 $D=636
M3123 532 531 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=38690 $Y=44992 $D=636
M3124 t_pxaa<0> 532 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=38690 $Y=46622 $D=636
M3125 vdd 527 b_pxaa<0> vdd hvtpfet l=6e-08 w=2.57e-06 $X=38950 $Y=1941 $D=636
M3126 vdd 528 527 vdd hvtpfet l=6e-08 w=1e-06 $X=38950 $Y=5141 $D=636
M3127 vdd 529 528 vdd hvtpfet l=6e-08 w=6e-07 $X=38950 $Y=8691 $D=636
M3128 529 525 vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=38950 $Y=10156 $D=636
M3129 530 525 vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=38950 $Y=40566 $D=636
M3130 vdd 530 531 vdd hvtpfet l=6e-08 w=6e-07 $X=38950 $Y=41842 $D=636
M3131 vdd 531 532 vdd hvtpfet l=6e-08 w=1e-06 $X=38950 $Y=44992 $D=636
M3132 vdd 532 t_pxaa<0> vdd hvtpfet l=6e-08 w=2.57e-06 $X=38950 $Y=46622 $D=636
M3133 1354 534 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=39025 $Y=29525 $D=636
M3134 533 aa<3> vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=39084 $Y=14280 $D=636
M3135 1355 317 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=39109 $Y=15520 $D=636
M3136 1356 317 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=39109 $Y=20589 $D=636
M3137 1357 317 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=39109 $Y=22440 $D=636
M3138 1358 317 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=39109 $Y=27509 $D=636
M3139 vdd clka 323 vdd hvtpfet l=6e-08 w=6e-07 $X=39174 $Y=33747 $D=636
M3140 293 535 vdd vdd hvtpfet l=6e-08 w=1.2e-06 $X=39185 $Y=35277 $D=636
M3141 495 539 1354 vdd hvtpfet l=6e-08 w=8.23e-07 $X=39285 $Y=29525 $D=636
M3142 549 537 1355 vdd hvtpfet l=6e-08 w=4.11e-07 $X=39379 $Y=15932 $D=636
M3143 550 538 1356 vdd hvtpfet l=6e-08 w=4.11e-07 $X=39379 $Y=20589 $D=636
M3144 551 537 1357 vdd hvtpfet l=6e-08 w=4.11e-07 $X=39379 $Y=22852 $D=636
M3145 552 538 1358 vdd hvtpfet l=6e-08 w=4.11e-07 $X=39379 $Y=27509 $D=636
M3146 323 clka vdd vdd hvtpfet l=6e-08 w=6e-07 $X=39434 $Y=33747 $D=636
M3147 vdd 538 537 vdd hvtpfet l=6e-08 w=4.11e-07 $X=39594 $Y=14280 $D=636
M3148 1359 546 549 vdd hvtpfet l=6e-08 w=4.11e-07 $X=39639 $Y=15932 $D=636
M3149 1360 546 550 vdd hvtpfet l=6e-08 w=4.11e-07 $X=39639 $Y=20589 $D=636
M3150 1361 533 551 vdd hvtpfet l=6e-08 w=4.11e-07 $X=39639 $Y=22852 $D=636
M3151 1362 533 552 vdd hvtpfet l=6e-08 w=4.11e-07 $X=39639 $Y=27509 $D=636
M3152 vdd clka 323 vdd hvtpfet l=6e-08 w=6e-07 $X=39694 $Y=33747 $D=636
M3153 r_sa_prea_n 293 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=39695 $Y=35277 $D=636
M3154 289 540 vdd vdd hvtpfet l=6e-08 w=1.2e-06 $X=39705 $Y=1736 $D=636
M3155 290 541 vdd vdd hvtpfet l=6e-08 w=1.2e-06 $X=39705 $Y=3566 $D=636
M3156 291 542 vdd vdd hvtpfet l=6e-08 w=1.2e-06 $X=39705 $Y=8196 $D=636
M3157 292 543 vdd vdd hvtpfet l=6e-08 w=1.2e-06 $X=39705 $Y=10026 $D=636
M3158 294 543 vdd vdd hvtpfet l=6e-08 w=1.2e-06 $X=39705 $Y=39907 $D=636
M3159 295 542 vdd vdd hvtpfet l=6e-08 w=1.2e-06 $X=39705 $Y=41737 $D=636
M3160 296 544 vdd vdd hvtpfet l=6e-08 w=1.2e-06 $X=39705 $Y=46367 $D=636
M3161 297 545 vdd vdd hvtpfet l=6e-08 w=1.2e-06 $X=39705 $Y=48197 $D=636
M3162 vdd stclka 539 vdd hvtpfet l=6e-08 w=4.11e-07 $X=39795 $Y=29937 $D=636
M3163 vdd 317 1359 vdd hvtpfet l=6e-08 w=8.23e-07 $X=39909 $Y=15520 $D=636
M3164 vdd 317 1360 vdd hvtpfet l=6e-08 w=8.23e-07 $X=39909 $Y=20589 $D=636
M3165 vdd 317 1361 vdd hvtpfet l=6e-08 w=8.23e-07 $X=39909 $Y=22440 $D=636
M3166 vdd 317 1362 vdd hvtpfet l=6e-08 w=8.23e-07 $X=39909 $Y=27509 $D=636
M3167 323 clka vdd vdd hvtpfet l=6e-08 w=6e-07 $X=39954 $Y=33747 $D=636
M3168 vdd 293 r_sa_prea_n vdd hvtpfet l=6e-08 w=1.43e-06 $X=39955 $Y=35277 $D=636
M3169 538 aa<2> vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=40104 $Y=14280 $D=636
M3170 rb_ca<1> 289 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=40215 $Y=1506 $D=636
M3171 rb_ca<3> 290 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=40215 $Y=3566 $D=636
M3172 rb_ma<1> 291 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=40215 $Y=7966 $D=636
M3173 rb_ma<3> 292 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=40215 $Y=10026 $D=636
M3174 r_sa_prea_n 293 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=40215 $Y=35277 $D=636
M3175 rt_ma<3> 294 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=40215 $Y=39677 $D=636
M3176 rt_ma<1> 295 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=40215 $Y=41737 $D=636
M3177 rt_ca<3> 296 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=40215 $Y=46137 $D=636
M3178 rt_ca<1> 297 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=40215 $Y=48197 $D=636
M3179 543 549 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=40419 $Y=15321 $D=636
M3180 1363 323 549 vdd hvtpfet l=6e-08 w=2.74e-07 $X=40419 $Y=16069 $D=636
M3181 1364 323 550 vdd hvtpfet l=6e-08 w=2.74e-07 $X=40419 $Y=20589 $D=636
M3182 553 550 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=40419 $Y=21405 $D=636
M3183 542 551 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=40419 $Y=22241 $D=636
M3184 1365 323 551 vdd hvtpfet l=6e-08 w=2.74e-07 $X=40419 $Y=22989 $D=636
M3185 1366 323 552 vdd hvtpfet l=6e-08 w=2.74e-07 $X=40419 $Y=27509 $D=636
M3186 554 552 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=40419 $Y=28325 $D=636
M3187 vdd 289 rb_ca<1> vdd hvtpfet l=6e-08 w=1.43e-06 $X=40475 $Y=1506 $D=636
M3188 vdd 290 rb_ca<3> vdd hvtpfet l=6e-08 w=1.43e-06 $X=40475 $Y=3566 $D=636
M3189 vdd 291 rb_ma<1> vdd hvtpfet l=6e-08 w=1.43e-06 $X=40475 $Y=7966 $D=636
M3190 vdd 292 rb_ma<3> vdd hvtpfet l=6e-08 w=1.43e-06 $X=40475 $Y=10026 $D=636
M3191 vdd 294 rt_ma<3> vdd hvtpfet l=6e-08 w=1.43e-06 $X=40475 $Y=39677 $D=636
M3192 vdd 295 rt_ma<1> vdd hvtpfet l=6e-08 w=1.43e-06 $X=40475 $Y=41737 $D=636
M3193 vdd 296 rt_ca<3> vdd hvtpfet l=6e-08 w=1.43e-06 $X=40475 $Y=46137 $D=636
M3194 vdd 297 rt_ca<1> vdd hvtpfet l=6e-08 w=1.43e-06 $X=40475 $Y=48197 $D=636
M3195 vdd 549 543 vdd hvtpfet l=6e-08 w=2.06e-07 $X=40679 $Y=15321 $D=636
M3196 vdd 543 1363 vdd hvtpfet l=6e-08 w=2.74e-07 $X=40679 $Y=16069 $D=636
M3197 vdd 553 1364 vdd hvtpfet l=6e-08 w=2.74e-07 $X=40679 $Y=20589 $D=636
M3198 vdd 550 553 vdd hvtpfet l=6e-08 w=2.06e-07 $X=40679 $Y=21405 $D=636
M3199 vdd 551 542 vdd hvtpfet l=6e-08 w=2.06e-07 $X=40679 $Y=22241 $D=636
M3200 vdd 542 1365 vdd hvtpfet l=6e-08 w=2.74e-07 $X=40679 $Y=22989 $D=636
M3201 vdd 554 1366 vdd hvtpfet l=6e-08 w=2.74e-07 $X=40679 $Y=27509 $D=636
M3202 vdd 552 554 vdd hvtpfet l=6e-08 w=2.06e-07 $X=40679 $Y=28325 $D=636
M3203 vdd 303 r_saea_n vdd hvtpfet l=6e-08 w=1.43e-06 $X=40725 $Y=35277 $D=636
M3204 rb_ca<1> 289 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=40735 $Y=1506 $D=636
M3205 rb_ca<3> 290 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=40735 $Y=3566 $D=636
M3206 rb_ma<1> 291 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=40735 $Y=7966 $D=636
M3207 rb_ma<3> 292 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=40735 $Y=10026 $D=636
M3208 rt_ma<3> 294 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=40735 $Y=39677 $D=636
M3209 rt_ma<1> 295 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=40735 $Y=41737 $D=636
M3210 rt_ca<3> 296 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=40735 $Y=46137 $D=636
M3211 rt_ca<1> 297 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=40735 $Y=48197 $D=636
M3212 r_saea_n 303 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=40985 $Y=35277 $D=636
M3213 vdd 299 rb_ca<0> vdd hvtpfet l=6e-08 w=1.43e-06 $X=41245 $Y=1506 $D=636
M3214 vdd 300 rb_ca<2> vdd hvtpfet l=6e-08 w=1.43e-06 $X=41245 $Y=3566 $D=636
M3215 vdd 301 rb_ma<0> vdd hvtpfet l=6e-08 w=1.43e-06 $X=41245 $Y=7966 $D=636
M3216 vdd 302 rb_ma<2> vdd hvtpfet l=6e-08 w=1.43e-06 $X=41245 $Y=10026 $D=636
M3217 vdd 303 r_saea_n vdd hvtpfet l=6e-08 w=1.43e-06 $X=41245 $Y=35277 $D=636
M3218 vdd 304 rt_ma<2> vdd hvtpfet l=6e-08 w=1.43e-06 $X=41245 $Y=39677 $D=636
M3219 vdd 305 rt_ma<0> vdd hvtpfet l=6e-08 w=1.43e-06 $X=41245 $Y=41737 $D=636
M3220 vdd 306 rt_ca<2> vdd hvtpfet l=6e-08 w=1.43e-06 $X=41245 $Y=46137 $D=636
M3221 vdd 307 rt_ca<0> vdd hvtpfet l=6e-08 w=1.43e-06 $X=41245 $Y=48197 $D=636
M3222 vdd clka 287 vdd hvtpfet l=6e-08 w=2.1e-06 $X=41495 $Y=23621 $D=636
M3223 vdd 340 288 vdd hvtpfet l=6e-08 w=2.1e-06 $X=41495 $Y=26587 $D=636
M3224 rb_ca<0> 299 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=41505 $Y=1506 $D=636
M3225 rb_ca<2> 300 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=41505 $Y=3566 $D=636
M3226 rb_ma<0> 301 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=41505 $Y=7966 $D=636
M3227 rb_ma<2> 302 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=41505 $Y=10026 $D=636
M3228 285 497 vdd vdd hvtpfet l=6e-08 w=1.2e-06 $X=41505 $Y=15067 $D=636
M3229 286 498 vdd vdd hvtpfet l=6e-08 w=1.2e-06 $X=41505 $Y=18424 $D=636
M3230 r_saea_n 303 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=41505 $Y=35277 $D=636
M3231 rt_ma<2> 304 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=41505 $Y=39677 $D=636
M3232 rt_ma<0> 305 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=41505 $Y=41737 $D=636
M3233 rt_ca<2> 306 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=41505 $Y=46137 $D=636
M3234 rt_ca<0> 307 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=41505 $Y=48197 $D=636
M3235 r_clk_dqa 287 vdd vdd hvtpfet l=6e-08 w=2.1e-06 $X=41755 $Y=23621 $D=636
M3236 r_clk_dqa_n 288 vdd vdd hvtpfet l=6e-08 w=2.1e-06 $X=41755 $Y=26587 $D=636
M3237 vdd 299 rb_ca<0> vdd hvtpfet l=6e-08 w=1.43e-06 $X=41765 $Y=1506 $D=636
M3238 vdd 300 rb_ca<2> vdd hvtpfet l=6e-08 w=1.43e-06 $X=41765 $Y=3566 $D=636
M3239 vdd 301 rb_ma<0> vdd hvtpfet l=6e-08 w=1.43e-06 $X=41765 $Y=7966 $D=636
M3240 vdd 302 rb_ma<2> vdd hvtpfet l=6e-08 w=1.43e-06 $X=41765 $Y=10026 $D=636
M3241 vdd 303 r_saea_n vdd hvtpfet l=6e-08 w=1.43e-06 $X=41765 $Y=35277 $D=636
M3242 vdd 304 rt_ma<2> vdd hvtpfet l=6e-08 w=1.43e-06 $X=41765 $Y=39677 $D=636
M3243 vdd 305 rt_ma<0> vdd hvtpfet l=6e-08 w=1.43e-06 $X=41765 $Y=41737 $D=636
M3244 vdd 306 rt_ca<2> vdd hvtpfet l=6e-08 w=1.43e-06 $X=41765 $Y=46137 $D=636
M3245 vdd 307 rt_ca<0> vdd hvtpfet l=6e-08 w=1.43e-06 $X=41765 $Y=48197 $D=636
M3246 rb_tm_prea_n 285 vdd vdd hvtpfet l=6e-08 w=2.145e-06 $X=42015 $Y=14887 $D=636
M3247 rt_tm_prea_n 286 vdd vdd hvtpfet l=6e-08 w=2.145e-06 $X=42015 $Y=17659 $D=636
M3248 vdd 287 r_clk_dqa vdd hvtpfet l=6e-08 w=2.1e-06 $X=42015 $Y=23621 $D=636
M3249 vdd 288 r_clk_dqa_n vdd hvtpfet l=6e-08 w=2.1e-06 $X=42015 $Y=26587 $D=636
M3250 r_lwea 284 vdd vdd hvtpfet l=6e-08 w=2.145e-06 $X=42015 $Y=32504 $D=636
M3251 vdd 555 299 vdd hvtpfet l=6e-08 w=1.2e-06 $X=42275 $Y=1736 $D=636
M3252 vdd 556 300 vdd hvtpfet l=6e-08 w=1.2e-06 $X=42275 $Y=3566 $D=636
M3253 vdd 554 301 vdd hvtpfet l=6e-08 w=1.2e-06 $X=42275 $Y=8196 $D=636
M3254 vdd 553 302 vdd hvtpfet l=6e-08 w=1.2e-06 $X=42275 $Y=10026 $D=636
M3255 vdd 285 rb_tm_prea_n vdd hvtpfet l=6e-08 w=2.145e-06 $X=42275 $Y=14887 $D=636
M3256 vdd 286 rt_tm_prea_n vdd hvtpfet l=6e-08 w=2.145e-06 $X=42275 $Y=17659 $D=636
M3257 r_clk_dqa 287 vdd vdd hvtpfet l=6e-08 w=2.1e-06 $X=42275 $Y=23621 $D=636
M3258 r_clk_dqa_n 288 vdd vdd hvtpfet l=6e-08 w=2.1e-06 $X=42275 $Y=26587 $D=636
M3259 vdd 284 r_lwea vdd hvtpfet l=6e-08 w=2.145e-06 $X=42275 $Y=32504 $D=636
M3260 vdd 557 303 vdd hvtpfet l=6e-08 w=1.2e-06 $X=42275 $Y=35277 $D=636
M3261 vdd 553 304 vdd hvtpfet l=6e-08 w=1.2e-06 $X=42275 $Y=39907 $D=636
M3262 vdd 554 305 vdd hvtpfet l=6e-08 w=1.2e-06 $X=42275 $Y=41737 $D=636
M3263 vdd 558 306 vdd hvtpfet l=6e-08 w=1.2e-06 $X=42275 $Y=46367 $D=636
M3264 vdd 559 307 vdd hvtpfet l=6e-08 w=1.2e-06 $X=42275 $Y=48197 $D=636
M3265 303 557 vdd vdd hvtpfet l=6e-08 w=1.2e-06 $X=42535 $Y=35277 $D=636
.ends

************************************************************************
* Library Name: XMC55_DPS
* Cell Name:    xmc55_dps_localc8io_bw
************************************************************************
.SUBCKT xmc55_dps_localc8io_bw b_bla<7> b_bla<6> b_bla<5> b_bla<4> b_bla<3> 
+ b_bla<2> b_bla<1> b_bla<0> b_bla_n<7> b_bla_n<6> b_bla_n<5> b_bla_n<4> 
+ b_bla_n<3> b_bla_n<2> b_bla_n<1> b_bla_n<0> b_blb<7> b_blb<6> b_blb<5> 
+ b_blb<4> b_blb<3> b_blb<2> b_blb<1> b_blb<0> b_blb_n<7> b_blb_n<6> 
+ b_blb_n<5> b_blb_n<4> b_blb_n<3> b_blb_n<2> b_blb_n<1> b_blb_n<0> b_ca<3> 
+ b_ca<2> b_ca<1> b_ca<0> b_cb<3> b_cb<2> b_cb<1> b_cb<0> b_ma<3> b_ma<2> 
+ b_ma<1> b_ma<0> b_mb<3> b_mb<2> b_mb<1> b_mb<0> b_tm_prea_n b_tm_preb_n 
+ bwena bwenb clk_dqa clk_dqa_n clk_dqb clk_dqb_n da db ddqa ddqa_n ddqb 
+ ddqb_n lwea lweb qa qb sa_prea_n sa_preb_n saea_n saeb_n t_bla<7> t_bla<6> 
+ t_bla<5> t_bla<4> t_bla<3> t_bla<2> t_bla<1> t_bla<0> t_bla_n<7> t_bla_n<6> 
+ t_bla_n<5> t_bla_n<4> t_bla_n<3> t_bla_n<2> t_bla_n<1> t_bla_n<0> t_blb<7> 
+ t_blb<6> t_blb<5> t_blb<4> t_blb<3> t_blb<2> t_blb<1> t_blb<0> t_blb_n<7> 
+ t_blb_n<6> t_blb_n<5> t_blb_n<4> t_blb_n<3> t_blb_n<2> t_blb_n<1> t_blb_n<0> 
+ t_ca<3> t_ca<2> t_ca<1> t_ca<0> t_cb<3> t_cb<2> t_cb<1> t_cb<0> t_ma<3> 
+ t_ma<2> t_ma<1> t_ma<0> t_mb<3> t_mb<2> t_mb<1> t_mb<0> t_tm_prea_n 
+ t_tm_preb_n vdd vss
** N=10332 EP=122 IP=0 FDC=1292
M0 195 8 b_blb<7> vss hvtnfet l=6e-08 w=6e-07 $X=210 $Y=2941 $D=616
M1 195 8 b_blb<7> vss hvtnfet l=6e-08 w=6e-07 $X=210 $Y=3201 $D=616
M2 204 16 b_bla_n<7> vss hvtnfet l=6e-08 w=6e-07 $X=210 $Y=3881 $D=616
M3 204 16 b_bla_n<7> vss hvtnfet l=6e-08 w=6e-07 $X=210 $Y=4141 $D=616
M4 t_bla_n<7> 17 204 vss hvtnfet l=6e-08 w=6e-07 $X=210 $Y=46932 $D=616
M5 204 17 t_bla_n<7> vss hvtnfet l=6e-08 w=6e-07 $X=210 $Y=47192 $D=616
M6 t_blb<7> 9 195 vss hvtnfet l=6e-08 w=6e-07 $X=210 $Y=47872 $D=616
M7 195 9 t_blb<7> vss hvtnfet l=6e-08 w=6e-07 $X=210 $Y=48132 $D=616
M8 8 5 vss vss hvtnfet l=6e-08 w=4e-07 $X=535 $Y=4836 $D=616
M9 549 b_cb<3> 5 vss hvtnfet l=6e-08 w=4e-07 $X=535 $Y=11331 $D=616
M10 550 5 2 vss hvtnfet l=6e-08 w=4e-07 $X=535 $Y=12191 $D=616
M11 551 6 3 vss hvtnfet l=6e-08 w=4e-07 $X=535 $Y=38542 $D=616
M12 552 t_cb<3> 6 vss hvtnfet l=6e-08 w=4e-07 $X=535 $Y=39402 $D=616
M13 9 6 vss vss hvtnfet l=6e-08 w=4e-07 $X=535 $Y=45897 $D=616
M14 215 vdd vss vss hvtnfet l=6e-08 w=2.5e-07 $X=540 $Y=17720 $D=616
M15 vss vss vss vss hvtnfet l=7e-08 w=3.2e-07 $X=610 $Y=33798 $D=616
M16 vss vss vss vss hvtnfet l=1.4e-07 w=7.5e-07 $X=650 $Y=34593 $D=616
M17 vss 11 8 vss hvtnfet l=6e-08 w=4e-07 $X=795 $Y=4836 $D=616
M18 vss b_mb<1> 549 vss hvtnfet l=6e-08 w=4e-07 $X=795 $Y=11331 $D=616
M19 vss 13 550 vss hvtnfet l=6e-08 w=4e-07 $X=795 $Y=12191 $D=616
M20 vss 14 551 vss hvtnfet l=6e-08 w=4e-07 $X=795 $Y=38542 $D=616
M21 vss t_mb<1> 552 vss hvtnfet l=6e-08 w=4e-07 $X=795 $Y=39402 $D=616
M22 vss 11 9 vss hvtnfet l=6e-08 w=4e-07 $X=795 $Y=45897 $D=616
M23 vss vdd 215 vss hvtnfet l=6e-08 w=2.5e-07 $X=800 $Y=17720 $D=616
M24 vss vss vss vss hvtnfet l=6e-08 w=3e-07 $X=867 $Y=31223 $D=616
M25 vss vss vss vss hvtnfet l=8e-08 w=3.75e-07 $X=890 $Y=33798 $D=616
M26 198 vdd vss vss hvtnfet l=6e-08 w=2e-07 $X=975 $Y=21427 $D=616
M27 199 vdd vss vss hvtnfet l=6e-08 w=2e-07 $X=975 $Y=23694 $D=616
M28 200 vdd vss vss hvtnfet l=6e-08 w=2e-07 $X=975 $Y=24394 $D=616
M29 201 vdd vss vss hvtnfet l=6e-08 w=2e-07 $X=975 $Y=24904 $D=616
M30 vss vss vss vss hvtnfet l=1.4e-07 w=7.5e-07 $X=990 $Y=34593 $D=616
M31 214 vdd vss vss hvtnfet l=6e-08 w=6e-07 $X=1007 $Y=26159 $D=616
M32 16 20 vss vss hvtnfet l=6e-08 w=4e-07 $X=1055 $Y=4836 $D=616
M33 553 b_ma<1> vss vss hvtnfet l=6e-08 w=4e-07 $X=1055 $Y=11331 $D=616
M34 554 22 vss vss hvtnfet l=6e-08 w=4e-07 $X=1055 $Y=12191 $D=616
M35 555 23 vss vss hvtnfet l=6e-08 w=4e-07 $X=1055 $Y=38542 $D=616
M36 556 t_ma<1> vss vss hvtnfet l=6e-08 w=4e-07 $X=1055 $Y=39402 $D=616
M37 17 20 vss vss hvtnfet l=6e-08 w=4e-07 $X=1055 $Y=45897 $D=616
M38 215 vdd vss vss hvtnfet l=6e-08 w=2.5e-07 $X=1060 $Y=17720 $D=616
M39 213 8 b_blb_n<7> vss hvtnfet l=6e-08 w=6e-07 $X=1100 $Y=2941 $D=616
M40 213 8 b_blb_n<7> vss hvtnfet l=6e-08 w=6e-07 $X=1100 $Y=3201 $D=616
M41 b_bla<7> 16 224 vss hvtnfet l=6e-08 w=6e-07 $X=1100 $Y=3881 $D=616
M42 b_bla<7> 16 224 vss hvtnfet l=6e-08 w=6e-07 $X=1100 $Y=4141 $D=616
M43 224 17 t_bla<7> vss hvtnfet l=6e-08 w=6e-07 $X=1100 $Y=46932 $D=616
M44 t_bla<7> 17 224 vss hvtnfet l=6e-08 w=6e-07 $X=1100 $Y=47192 $D=616
M45 t_blb_n<7> 9 213 vss hvtnfet l=6e-08 w=6e-07 $X=1100 $Y=47872 $D=616
M46 213 9 t_blb_n<7> vss hvtnfet l=6e-08 w=6e-07 $X=1100 $Y=48132 $D=616
M47 vss vss vss vss hvtnfet l=6e-08 w=3e-07 $X=1127 $Y=31223 $D=616
M48 vss vss vss vss hvtnfet l=8e-08 w=3.75e-07 $X=1170 $Y=33798 $D=616
M49 vss vdd 214 vss hvtnfet l=6e-08 w=6e-07 $X=1267 $Y=26159 $D=616
M50 vss 18 16 vss hvtnfet l=6e-08 w=4e-07 $X=1315 $Y=4836 $D=616
M51 18 b_ca<3> 553 vss hvtnfet l=6e-08 w=4e-07 $X=1315 $Y=11331 $D=616
M52 25 18 554 vss hvtnfet l=6e-08 w=4e-07 $X=1315 $Y=12191 $D=616
M53 26 19 555 vss hvtnfet l=6e-08 w=4e-07 $X=1315 $Y=38542 $D=616
M54 19 t_ca<3> 556 vss hvtnfet l=6e-08 w=4e-07 $X=1315 $Y=39402 $D=616
M55 vss 19 17 vss hvtnfet l=6e-08 w=4e-07 $X=1315 $Y=45897 $D=616
M56 vss vdd 215 vss hvtnfet l=6e-08 w=2.5e-07 $X=1320 $Y=17720 $D=616
M57 vss vss vss vss hvtnfet l=1.4e-07 w=7.5e-07 $X=1330 $Y=34593 $D=616
M58 vss vss vss vss hvtnfet l=8e-08 w=3.75e-07 $X=1450 $Y=33798 $D=616
M59 vss vss vss vss hvtnfet l=1.4e-07 w=7.5e-07 $X=1670 $Y=34593 $D=616
M60 vss vss vss vss hvtnfet l=8e-08 w=3.75e-07 $X=1730 $Y=33798 $D=616
M61 239 vdd 242 vss hvtnfet l=6e-08 w=8e-07 $X=1787 $Y=26159 $D=616
M62 233 vdd vss vss hvtnfet l=1.4e-07 w=2.1e-07 $X=1805 $Y=14550 $D=616
M63 234 vdd vss vss hvtnfet l=1.4e-07 w=2.1e-07 $X=1805 $Y=16760 $D=616
M64 249 vdd vss vss hvtnfet l=6e-08 w=3e-07 $X=1830 $Y=17670 $D=616
M65 vss vss vss vss hvtnfet l=6e-08 w=3.2e-07 $X=1920 $Y=19812 $D=616
M66 vss vss vss vss hvtnfet l=6e-08 w=3.2e-07 $X=1920 $Y=20072 $D=616
M67 vss vss vss vss hvtnfet l=6e-08 w=3.2e-07 $X=1920 $Y=21162 $D=616
M68 vss vss vss vss hvtnfet l=6e-08 w=3.2e-07 $X=1920 $Y=21422 $D=616
M69 vss vss vss vss hvtnfet l=6e-08 w=3.2e-07 $X=1920 $Y=21682 $D=616
M70 vss vss vss vss hvtnfet l=6e-08 w=3.2e-07 $X=1920 $Y=21942 $D=616
M71 vss vss vss vss hvtnfet l=6e-08 w=3.2e-07 $X=1920 $Y=22762 $D=616
M72 vss vss vss vss hvtnfet l=6e-08 w=3.2e-07 $X=1920 $Y=23879 $D=616
M73 vss vss vss vss hvtnfet l=6e-08 w=3.2e-07 $X=1920 $Y=24139 $D=616
M74 vss vss vss vss hvtnfet l=6e-08 w=3.2e-07 $X=1920 $Y=24399 $D=616
M75 vss vss vss vss hvtnfet l=6e-08 w=3.2e-07 $X=1920 $Y=24659 $D=616
M76 vss vss vss vss hvtnfet l=8e-08 w=3.75e-07 $X=2010 $Y=33798 $D=616
M77 vss vss vss vss hvtnfet l=1.4e-07 w=7.5e-07 $X=2010 $Y=34593 $D=616
M78 vss vss vss vss hvtnfet l=6e-08 w=3e-07 $X=2037 $Y=31223 $D=616
M79 242 vdd 239 vss hvtnfet l=6e-08 w=8e-07 $X=2047 $Y=26159 $D=616
M80 vss vdd 249 vss hvtnfet l=6e-08 w=3e-07 $X=2090 $Y=17670 $D=616
M81 213 39 b_blb_n<6> vss hvtnfet l=6e-08 w=6e-07 $X=2120 $Y=2941 $D=616
M82 213 39 b_blb_n<6> vss hvtnfet l=6e-08 w=6e-07 $X=2120 $Y=3201 $D=616
M83 b_bla<6> 35 224 vss hvtnfet l=6e-08 w=6e-07 $X=2120 $Y=3881 $D=616
M84 b_bla<6> 35 224 vss hvtnfet l=6e-08 w=6e-07 $X=2120 $Y=4141 $D=616
M85 224 36 t_bla<6> vss hvtnfet l=6e-08 w=6e-07 $X=2120 $Y=46932 $D=616
M86 t_bla<6> 36 224 vss hvtnfet l=6e-08 w=6e-07 $X=2120 $Y=47192 $D=616
M87 t_blb_n<6> 40 213 vss hvtnfet l=6e-08 w=6e-07 $X=2120 $Y=47872 $D=616
M88 213 40 t_blb_n<6> vss hvtnfet l=6e-08 w=6e-07 $X=2120 $Y=48132 $D=616
M89 vss vdd 233 vss hvtnfet l=1.4e-07 w=2.1e-07 $X=2145 $Y=14550 $D=616
M90 vss vdd 234 vss hvtnfet l=1.4e-07 w=2.1e-07 $X=2145 $Y=16760 $D=616
M91 vss vss vss vss hvtnfet l=8e-08 w=3.75e-07 $X=2290 $Y=33798 $D=616
M92 vss vss vss vss hvtnfet l=6e-08 w=3e-07 $X=2297 $Y=31223 $D=616
M93 vss vdd 242 vss hvtnfet l=6e-08 w=8e-07 $X=2307 $Y=26159 $D=616
M94 249 vdd vss vss hvtnfet l=6e-08 w=3e-07 $X=2350 $Y=17670 $D=616
M95 vss vss vss vss hvtnfet l=1.4e-07 w=7.5e-07 $X=2350 $Y=34593 $D=616
M96 35 30 vss vss hvtnfet l=6e-08 w=4e-07 $X=2445 $Y=4836 $D=616
M97 557 b_ca<2> 30 vss hvtnfet l=6e-08 w=4e-07 $X=2445 $Y=11331 $D=616
M98 558 30 33 vss hvtnfet l=6e-08 w=4e-07 $X=2445 $Y=12191 $D=616
M99 559 31 34 vss hvtnfet l=6e-08 w=4e-07 $X=2445 $Y=38542 $D=616
M100 560 t_ca<2> 31 vss hvtnfet l=6e-08 w=4e-07 $X=2445 $Y=39402 $D=616
M101 36 31 vss vss hvtnfet l=6e-08 w=4e-07 $X=2445 $Y=45897 $D=616
M102 vss vss vss vss hvtnfet l=6e-08 w=3e-07 $X=2557 $Y=31223 $D=616
M103 242 vdd vss vss hvtnfet l=6e-08 w=8e-07 $X=2567 $Y=26159 $D=616
M104 vss vss vss vss hvtnfet l=8e-08 w=3.75e-07 $X=2570 $Y=33798 $D=616
M105 vss vdd 249 vss hvtnfet l=6e-08 w=3e-07 $X=2610 $Y=17670 $D=616
M106 vss vss vss vss hvtnfet l=1.4e-07 w=7.5e-07 $X=2690 $Y=34593 $D=616
M107 vss 20 35 vss hvtnfet l=6e-08 w=4e-07 $X=2705 $Y=4836 $D=616
M108 vss b_ma<1> 557 vss hvtnfet l=6e-08 w=4e-07 $X=2705 $Y=11331 $D=616
M109 vss 22 558 vss hvtnfet l=6e-08 w=4e-07 $X=2705 $Y=12191 $D=616
M110 vss 23 559 vss hvtnfet l=6e-08 w=4e-07 $X=2705 $Y=38542 $D=616
M111 vss t_ma<1> 560 vss hvtnfet l=6e-08 w=4e-07 $X=2705 $Y=39402 $D=616
M112 vss 20 36 vss hvtnfet l=6e-08 w=4e-07 $X=2705 $Y=45897 $D=616
M113 247 vdd vss vss hvtnfet l=1.4e-07 w=2.1e-07 $X=2735 $Y=14550 $D=616
M114 248 vdd vss vss hvtnfet l=1.4e-07 w=2.1e-07 $X=2735 $Y=16760 $D=616
M115 vss vss vss vss hvtnfet l=6e-08 w=3e-07 $X=2817 $Y=31223 $D=616
M116 vss vss vss vss hvtnfet l=8e-08 w=3.75e-07 $X=2850 $Y=33798 $D=616
M117 249 vdd vss vss hvtnfet l=6e-08 w=3e-07 $X=2870 $Y=17670 $D=616
M118 39 11 vss vss hvtnfet l=6e-08 w=4e-07 $X=2965 $Y=4836 $D=616
M119 561 b_mb<1> vss vss hvtnfet l=6e-08 w=4e-07 $X=2965 $Y=11331 $D=616
M120 562 13 vss vss hvtnfet l=6e-08 w=4e-07 $X=2965 $Y=12191 $D=616
M121 563 14 vss vss hvtnfet l=6e-08 w=4e-07 $X=2965 $Y=38542 $D=616
M122 564 t_mb<1> vss vss hvtnfet l=6e-08 w=4e-07 $X=2965 $Y=39402 $D=616
M123 40 11 vss vss hvtnfet l=6e-08 w=4e-07 $X=2965 $Y=45897 $D=616
M124 195 39 b_blb<6> vss hvtnfet l=6e-08 w=6e-07 $X=3010 $Y=2941 $D=616
M125 195 39 b_blb<6> vss hvtnfet l=6e-08 w=6e-07 $X=3010 $Y=3201 $D=616
M126 204 35 b_bla_n<6> vss hvtnfet l=6e-08 w=6e-07 $X=3010 $Y=3881 $D=616
M127 204 35 b_bla_n<6> vss hvtnfet l=6e-08 w=6e-07 $X=3010 $Y=4141 $D=616
M128 t_bla_n<6> 36 204 vss hvtnfet l=6e-08 w=6e-07 $X=3010 $Y=46932 $D=616
M129 204 36 t_bla_n<6> vss hvtnfet l=6e-08 w=6e-07 $X=3010 $Y=47192 $D=616
M130 t_blb<6> 40 195 vss hvtnfet l=6e-08 w=6e-07 $X=3010 $Y=47872 $D=616
M131 195 40 t_blb<6> vss hvtnfet l=6e-08 w=6e-07 $X=3010 $Y=48132 $D=616
M132 vss vss vss vss hvtnfet l=1.4e-07 w=7.5e-07 $X=3030 $Y=34593 $D=616
M133 vss vdd 247 vss hvtnfet l=1.4e-07 w=2.1e-07 $X=3075 $Y=14550 $D=616
M134 vss vdd 248 vss hvtnfet l=1.4e-07 w=2.1e-07 $X=3075 $Y=16760 $D=616
M135 256 vdd vss vss hvtnfet l=6e-08 w=6e-07 $X=3077 $Y=26159 $D=616
M136 vss vdd 249 vss hvtnfet l=6e-08 w=3e-07 $X=3130 $Y=17670 $D=616
M137 vss vss vss vss hvtnfet l=7e-08 w=3.2e-07 $X=3140 $Y=33798 $D=616
M138 vss 37 39 vss hvtnfet l=6e-08 w=4e-07 $X=3225 $Y=4836 $D=616
M139 37 b_cb<2> 561 vss hvtnfet l=6e-08 w=4e-07 $X=3225 $Y=11331 $D=616
M140 41 37 562 vss hvtnfet l=6e-08 w=4e-07 $X=3225 $Y=12191 $D=616
M141 42 38 563 vss hvtnfet l=6e-08 w=4e-07 $X=3225 $Y=38542 $D=616
M142 38 t_cb<2> 564 vss hvtnfet l=6e-08 w=4e-07 $X=3225 $Y=39402 $D=616
M143 vss 38 40 vss hvtnfet l=6e-08 w=4e-07 $X=3225 $Y=45897 $D=616
M144 vss vdd 256 vss hvtnfet l=6e-08 w=6e-07 $X=3337 $Y=26159 $D=616
M145 195 54 b_blb<5> vss hvtnfet l=6e-08 w=6e-07 $X=4030 $Y=2941 $D=616
M146 195 54 b_blb<5> vss hvtnfet l=6e-08 w=6e-07 $X=4030 $Y=3201 $D=616
M147 204 62 b_bla_n<5> vss hvtnfet l=6e-08 w=6e-07 $X=4030 $Y=3881 $D=616
M148 204 62 b_bla_n<5> vss hvtnfet l=6e-08 w=6e-07 $X=4030 $Y=4141 $D=616
M149 t_bla_n<5> 63 204 vss hvtnfet l=6e-08 w=6e-07 $X=4030 $Y=46932 $D=616
M150 204 63 t_bla_n<5> vss hvtnfet l=6e-08 w=6e-07 $X=4030 $Y=47192 $D=616
M151 t_blb<5> 55 195 vss hvtnfet l=6e-08 w=6e-07 $X=4030 $Y=47872 $D=616
M152 195 55 t_blb<5> vss hvtnfet l=6e-08 w=6e-07 $X=4030 $Y=48132 $D=616
M153 204 61 vss vss hvtnfet l=6e-08 w=6e-07 $X=4243 $Y=26159 $D=616
M154 54 48 vss vss hvtnfet l=6e-08 w=4e-07 $X=4355 $Y=4836 $D=616
M155 565 b_cb<1> 48 vss hvtnfet l=6e-08 w=4e-07 $X=4355 $Y=11331 $D=616
M156 566 48 45 vss hvtnfet l=6e-08 w=4e-07 $X=4355 $Y=12191 $D=616
M157 567 49 46 vss hvtnfet l=6e-08 w=4e-07 $X=4355 $Y=38542 $D=616
M158 568 t_cb<1> 49 vss hvtnfet l=6e-08 w=4e-07 $X=4355 $Y=39402 $D=616
M159 55 49 vss vss hvtnfet l=6e-08 w=4e-07 $X=4355 $Y=45897 $D=616
M160 vss vdd 270 vss hvtnfet l=6e-08 w=3e-07 $X=4393 $Y=31223 $D=616
M161 vss bwena 64 vss hvtnfet l=1.4e-07 w=2.1e-07 $X=4425 $Y=14555 $D=616
M162 vss 56 76 vss hvtnfet l=1.4e-07 w=2.1e-07 $X=4425 $Y=16755 $D=616
M163 vss 57 ddqa_n vss hvtnfet l=7e-08 w=3.2e-07 $X=4430 $Y=33798 $D=616
M164 288 vdd vss vss hvtnfet l=6e-08 w=3e-07 $X=4450 $Y=17670 $D=616
M165 57 59 310 vss hvtnfet l=1.4e-07 w=7.5e-07 $X=4470 $Y=34593 $D=616
M166 vss 61 204 vss hvtnfet l=6e-08 w=6e-07 $X=4503 $Y=26159 $D=616
M167 vss 11 54 vss hvtnfet l=6e-08 w=4e-07 $X=4615 $Y=4836 $D=616
M168 vss b_mb<1> 565 vss hvtnfet l=6e-08 w=4e-07 $X=4615 $Y=11331 $D=616
M169 vss 13 566 vss hvtnfet l=6e-08 w=4e-07 $X=4615 $Y=12191 $D=616
M170 vss 14 567 vss hvtnfet l=6e-08 w=4e-07 $X=4615 $Y=38542 $D=616
M171 vss t_mb<1> 568 vss hvtnfet l=6e-08 w=4e-07 $X=4615 $Y=39402 $D=616
M172 vss 11 55 vss hvtnfet l=6e-08 w=4e-07 $X=4615 $Y=45897 $D=616
M173 vss vdd 288 vss hvtnfet l=6e-08 w=3e-07 $X=4710 $Y=17670 $D=616
M174 310 60 vss vss hvtnfet l=8e-08 w=3.75e-07 $X=4710 $Y=33798 $D=616
M175 72 64 vss vss hvtnfet l=1.4e-07 w=2.1e-07 $X=4765 $Y=14555 $D=616
M176 56 75 vss vss hvtnfet l=1.4e-07 w=2.1e-07 $X=4765 $Y=16755 $D=616
M177 310 59 57 vss hvtnfet l=1.4e-07 w=7.5e-07 $X=4810 $Y=34593 $D=616
M178 62 20 vss vss hvtnfet l=6e-08 w=4e-07 $X=4875 $Y=4836 $D=616
M179 569 b_ma<1> vss vss hvtnfet l=6e-08 w=4e-07 $X=4875 $Y=11331 $D=616
M180 570 22 vss vss hvtnfet l=6e-08 w=4e-07 $X=4875 $Y=12191 $D=616
M181 571 23 vss vss hvtnfet l=6e-08 w=4e-07 $X=4875 $Y=38542 $D=616
M182 572 t_ma<1> vss vss hvtnfet l=6e-08 w=4e-07 $X=4875 $Y=39402 $D=616
M183 63 20 vss vss hvtnfet l=6e-08 w=4e-07 $X=4875 $Y=45897 $D=616
M184 573 60 vss vss hvtnfet l=6e-08 w=3e-07 $X=4903 $Y=31223 $D=616
M185 213 54 b_blb_n<5> vss hvtnfet l=6e-08 w=6e-07 $X=4920 $Y=2941 $D=616
M186 213 54 b_blb_n<5> vss hvtnfet l=6e-08 w=6e-07 $X=4920 $Y=3201 $D=616
M187 b_bla<5> 62 224 vss hvtnfet l=6e-08 w=6e-07 $X=4920 $Y=3881 $D=616
M188 b_bla<5> 62 224 vss hvtnfet l=6e-08 w=6e-07 $X=4920 $Y=4141 $D=616
M189 224 63 t_bla<5> vss hvtnfet l=6e-08 w=6e-07 $X=4920 $Y=46932 $D=616
M190 t_bla<5> 63 224 vss hvtnfet l=6e-08 w=6e-07 $X=4920 $Y=47192 $D=616
M191 t_blb_n<5> 55 213 vss hvtnfet l=6e-08 w=6e-07 $X=4920 $Y=47872 $D=616
M192 213 55 t_blb_n<5> vss hvtnfet l=6e-08 w=6e-07 $X=4920 $Y=48132 $D=616
M193 288 vdd vss vss hvtnfet l=6e-08 w=3e-07 $X=4970 $Y=17670 $D=616
M194 vss 60 310 vss hvtnfet l=8e-08 w=3.75e-07 $X=4990 $Y=33798 $D=616
M195 vss 68 293 vss hvtnfet l=6e-08 w=8e-07 $X=5013 $Y=26159 $D=616
M196 82 57 573 vss hvtnfet l=6e-08 w=3e-07 $X=5093 $Y=31223 $D=616
M197 vss 65 62 vss hvtnfet l=6e-08 w=4e-07 $X=5135 $Y=4836 $D=616
M198 65 b_ca<1> 569 vss hvtnfet l=6e-08 w=4e-07 $X=5135 $Y=11331 $D=616
M199 69 65 570 vss hvtnfet l=6e-08 w=4e-07 $X=5135 $Y=12191 $D=616
M200 70 66 571 vss hvtnfet l=6e-08 w=4e-07 $X=5135 $Y=38542 $D=616
M201 66 t_ca<1> 572 vss hvtnfet l=6e-08 w=4e-07 $X=5135 $Y=39402 $D=616
M202 vss 66 63 vss hvtnfet l=6e-08 w=4e-07 $X=5135 $Y=45897 $D=616
M203 59 57 310 vss hvtnfet l=1.4e-07 w=7.5e-07 $X=5150 $Y=34593 $D=616
M204 vss vdd 288 vss hvtnfet l=6e-08 w=3e-07 $X=5230 $Y=17670 $D=616
M205 310 60 vss vss hvtnfet l=8e-08 w=3.75e-07 $X=5270 $Y=33798 $D=616
M206 293 68 vss vss hvtnfet l=6e-08 w=8e-07 $X=5273 $Y=26159 $D=616
M207 574 67 82 vss hvtnfet l=6e-08 w=3e-07 $X=5353 $Y=31223 $D=616
M208 vss 72 85 vss hvtnfet l=1.4e-07 w=2.1e-07 $X=5355 $Y=14555 $D=616
M209 vss 80 75 vss hvtnfet l=1.4e-07 w=2.1e-07 $X=5355 $Y=16755 $D=616
M210 qa 67 vss vss hvtnfet l=6e-08 w=4.5e-07 $X=5435 $Y=19812 $D=616
M211 vss 67 qa vss hvtnfet l=6e-08 w=4.5e-07 $X=5435 $Y=20072 $D=616
M212 575 76 vss vss hvtnfet l=6e-08 w=3.2e-07 $X=5435 $Y=21012 $D=616
M213 575 71 73 vss hvtnfet l=6e-08 w=3.2e-07 $X=5435 $Y=21202 $D=616
M214 576 53 73 vss hvtnfet l=6e-08 w=1.4e-07 $X=5435 $Y=21477 $D=616
M215 vss 51 576 vss hvtnfet l=6e-08 w=1.4e-07 $X=5435 $Y=21667 $D=616
M216 53 73 vss vss hvtnfet l=6e-08 w=2.1e-07 $X=5435 $Y=21942 $D=616
M217 vss 73 61 vss hvtnfet l=6e-08 w=3.2e-07 $X=5435 $Y=22762 $D=616
M218 577 77 vss vss hvtnfet l=6e-08 w=3.2e-07 $X=5435 $Y=23729 $D=616
M219 577 71 74 vss hvtnfet l=6e-08 w=3.2e-07 $X=5435 $Y=23919 $D=616
M220 578 52 74 vss hvtnfet l=6e-08 w=1.4e-07 $X=5435 $Y=24194 $D=616
M221 vss 51 578 vss hvtnfet l=6e-08 w=1.4e-07 $X=5435 $Y=24384 $D=616
M222 52 74 vss vss hvtnfet l=6e-08 w=2.1e-07 $X=5435 $Y=24659 $D=616
M223 288 vdd vss vss hvtnfet l=6e-08 w=3e-07 $X=5490 $Y=17670 $D=616
M224 310 57 59 vss hvtnfet l=1.4e-07 w=7.5e-07 $X=5490 $Y=34593 $D=616
M225 20 lwea 293 vss hvtnfet l=6e-08 w=8e-07 $X=5533 $Y=26159 $D=616
M226 vss saea_n 574 vss hvtnfet l=6e-08 w=3e-07 $X=5543 $Y=31223 $D=616
M227 vss 60 310 vss hvtnfet l=8e-08 w=3.75e-07 $X=5550 $Y=33798 $D=616
M228 77 85 vss vss hvtnfet l=1.4e-07 w=2.1e-07 $X=5695 $Y=14555 $D=616
M229 80 da vss vss hvtnfet l=1.4e-07 w=2.1e-07 $X=5695 $Y=16755 $D=616
M230 vss vdd 288 vss hvtnfet l=6e-08 w=3e-07 $X=5750 $Y=17670 $D=616
M231 293 lwea 20 vss hvtnfet l=6e-08 w=8e-07 $X=5793 $Y=26159 $D=616
M232 310 60 vss vss hvtnfet l=8e-08 w=3.75e-07 $X=5830 $Y=33798 $D=616
M233 57 59 310 vss hvtnfet l=1.4e-07 w=7.5e-07 $X=5830 $Y=34593 $D=616
M234 213 101 b_blb_n<4> vss hvtnfet l=6e-08 w=6e-07 $X=5940 $Y=2941 $D=616
M235 213 101 b_blb_n<4> vss hvtnfet l=6e-08 w=6e-07 $X=5940 $Y=3201 $D=616
M236 b_bla<4> 94 224 vss hvtnfet l=6e-08 w=6e-07 $X=5940 $Y=3881 $D=616
M237 b_bla<4> 94 224 vss hvtnfet l=6e-08 w=6e-07 $X=5940 $Y=4141 $D=616
M238 224 95 t_bla<4> vss hvtnfet l=6e-08 w=6e-07 $X=5940 $Y=46932 $D=616
M239 t_bla<4> 95 224 vss hvtnfet l=6e-08 w=6e-07 $X=5940 $Y=47192 $D=616
M240 t_blb_n<4> 102 213 vss hvtnfet l=6e-08 w=6e-07 $X=5940 $Y=47872 $D=616
M241 213 102 t_blb_n<4> vss hvtnfet l=6e-08 w=6e-07 $X=5940 $Y=48132 $D=616
M242 vss 60 310 vss hvtnfet l=8e-08 w=3.75e-07 $X=6110 $Y=33798 $D=616
M243 310 59 57 vss hvtnfet l=1.4e-07 w=7.5e-07 $X=6170 $Y=34593 $D=616
M244 22 b_tm_prea_n vss vss hvtnfet l=6e-08 w=2.5e-07 $X=6260 $Y=17720 $D=616
M245 94 88 vss vss hvtnfet l=6e-08 w=4e-07 $X=6265 $Y=4836 $D=616
M246 579 b_ca<0> 88 vss hvtnfet l=6e-08 w=4e-07 $X=6265 $Y=11331 $D=616
M247 580 88 91 vss hvtnfet l=6e-08 w=4e-07 $X=6265 $Y=12191 $D=616
M248 581 89 92 vss hvtnfet l=6e-08 w=4e-07 $X=6265 $Y=38542 $D=616
M249 582 t_ca<0> 89 vss hvtnfet l=6e-08 w=4e-07 $X=6265 $Y=39402 $D=616
M250 95 89 vss vss hvtnfet l=6e-08 w=4e-07 $X=6265 $Y=45897 $D=616
M251 224 73 vss vss hvtnfet l=6e-08 w=6e-07 $X=6313 $Y=26159 $D=616
M252 310 60 vss vss hvtnfet l=8e-08 w=3.75e-07 $X=6390 $Y=33798 $D=616
M253 vss 82 67 vss hvtnfet l=6e-08 w=3e-07 $X=6453 $Y=31223 $D=616
M254 71 clk_dqa vss vss hvtnfet l=6e-08 w=2e-07 $X=6465 $Y=21427 $D=616
M255 51 clk_dqa_n vss vss hvtnfet l=6e-08 w=2e-07 $X=6465 $Y=23694 $D=616
M256 98 74 vss vss hvtnfet l=6e-08 w=2e-07 $X=6465 $Y=24394 $D=616
M257 68 98 vss vss hvtnfet l=6e-08 w=2e-07 $X=6465 $Y=24904 $D=616
M258 59 57 310 vss hvtnfet l=1.4e-07 w=7.5e-07 $X=6510 $Y=34593 $D=616
M259 vss b_tm_prea_n 22 vss hvtnfet l=6e-08 w=2.5e-07 $X=6520 $Y=17720 $D=616
M260 vss 20 94 vss hvtnfet l=6e-08 w=4e-07 $X=6525 $Y=4836 $D=616
M261 vss b_ma<1> 579 vss hvtnfet l=6e-08 w=4e-07 $X=6525 $Y=11331 $D=616
M262 vss 22 580 vss hvtnfet l=6e-08 w=4e-07 $X=6525 $Y=12191 $D=616
M263 vss 23 581 vss hvtnfet l=6e-08 w=4e-07 $X=6525 $Y=38542 $D=616
M264 vss t_ma<1> 582 vss hvtnfet l=6e-08 w=4e-07 $X=6525 $Y=39402 $D=616
M265 vss 20 95 vss hvtnfet l=6e-08 w=4e-07 $X=6525 $Y=45897 $D=616
M266 vss 73 224 vss hvtnfet l=6e-08 w=6e-07 $X=6573 $Y=26159 $D=616
M267 vss 60 310 vss hvtnfet l=8e-08 w=3.75e-07 $X=6670 $Y=33798 $D=616
M268 60 saea_n vss vss hvtnfet l=6e-08 w=3e-07 $X=6713 $Y=31223 $D=616
M269 23 t_tm_prea_n vss vss hvtnfet l=6e-08 w=2.5e-07 $X=6780 $Y=17720 $D=616
M270 101 11 vss vss hvtnfet l=6e-08 w=4e-07 $X=6785 $Y=4836 $D=616
M271 583 b_mb<1> vss vss hvtnfet l=6e-08 w=4e-07 $X=6785 $Y=11331 $D=616
M272 584 13 vss vss hvtnfet l=6e-08 w=4e-07 $X=6785 $Y=12191 $D=616
M273 585 14 vss vss hvtnfet l=6e-08 w=4e-07 $X=6785 $Y=38542 $D=616
M274 586 t_mb<1> vss vss hvtnfet l=6e-08 w=4e-07 $X=6785 $Y=39402 $D=616
M275 102 11 vss vss hvtnfet l=6e-08 w=4e-07 $X=6785 $Y=45897 $D=616
M276 195 101 b_blb<4> vss hvtnfet l=6e-08 w=6e-07 $X=6830 $Y=2941 $D=616
M277 195 101 b_blb<4> vss hvtnfet l=6e-08 w=6e-07 $X=6830 $Y=3201 $D=616
M278 204 94 b_bla_n<4> vss hvtnfet l=6e-08 w=6e-07 $X=6830 $Y=3881 $D=616
M279 204 94 b_bla_n<4> vss hvtnfet l=6e-08 w=6e-07 $X=6830 $Y=4141 $D=616
M280 t_bla_n<4> 95 204 vss hvtnfet l=6e-08 w=6e-07 $X=6830 $Y=46932 $D=616
M281 204 95 t_bla_n<4> vss hvtnfet l=6e-08 w=6e-07 $X=6830 $Y=47192 $D=616
M282 t_blb<4> 102 195 vss hvtnfet l=6e-08 w=6e-07 $X=6830 $Y=47872 $D=616
M283 195 102 t_blb<4> vss hvtnfet l=6e-08 w=6e-07 $X=6830 $Y=48132 $D=616
M284 310 57 59 vss hvtnfet l=1.4e-07 w=7.5e-07 $X=6850 $Y=34593 $D=616
M285 ddqa 59 vss vss hvtnfet l=7e-08 w=3.2e-07 $X=6960 $Y=33798 $D=616
M286 vss t_tm_prea_n 23 vss hvtnfet l=6e-08 w=2.5e-07 $X=7040 $Y=17720 $D=616
M287 vss 99 101 vss hvtnfet l=6e-08 w=4e-07 $X=7045 $Y=4836 $D=616
M288 99 b_cb<0> 583 vss hvtnfet l=6e-08 w=4e-07 $X=7045 $Y=11331 $D=616
M289 103 99 584 vss hvtnfet l=6e-08 w=4e-07 $X=7045 $Y=12191 $D=616
M290 104 100 585 vss hvtnfet l=6e-08 w=4e-07 $X=7045 $Y=38542 $D=616
M291 100 t_cb<0> 586 vss hvtnfet l=6e-08 w=4e-07 $X=7045 $Y=39402 $D=616
M292 vss 100 102 vss hvtnfet l=6e-08 w=4e-07 $X=7045 $Y=45897 $D=616
M293 316 59 vss vss hvtnfet l=6e-08 w=3e-07 $X=7223 $Y=31223 $D=616
M294 195 114 b_blb<3> vss hvtnfet l=6e-08 w=6e-07 $X=7850 $Y=2941 $D=616
M295 195 114 b_blb<3> vss hvtnfet l=6e-08 w=6e-07 $X=7850 $Y=3201 $D=616
M296 204 124 b_bla_n<3> vss hvtnfet l=6e-08 w=6e-07 $X=7850 $Y=3881 $D=616
M297 204 124 b_bla_n<3> vss hvtnfet l=6e-08 w=6e-07 $X=7850 $Y=4141 $D=616
M298 t_bla_n<3> 125 204 vss hvtnfet l=6e-08 w=6e-07 $X=7850 $Y=46932 $D=616
M299 204 125 t_bla_n<3> vss hvtnfet l=6e-08 w=6e-07 $X=7850 $Y=47192 $D=616
M300 t_blb<3> 115 195 vss hvtnfet l=6e-08 w=6e-07 $X=7850 $Y=47872 $D=616
M301 195 115 t_blb<3> vss hvtnfet l=6e-08 w=6e-07 $X=7850 $Y=48132 $D=616
M302 vss 108 323 vss hvtnfet l=6e-08 w=3e-07 $X=7997 $Y=31223 $D=616
M303 114 111 vss vss hvtnfet l=6e-08 w=4e-07 $X=8175 $Y=4836 $D=616
M304 587 b_cb<3> 111 vss hvtnfet l=6e-08 w=4e-07 $X=8175 $Y=11331 $D=616
M305 588 111 109 vss hvtnfet l=6e-08 w=4e-07 $X=8175 $Y=12191 $D=616
M306 589 112 110 vss hvtnfet l=6e-08 w=4e-07 $X=8175 $Y=38542 $D=616
M307 590 t_cb<3> 112 vss hvtnfet l=6e-08 w=4e-07 $X=8175 $Y=39402 $D=616
M308 115 112 vss vss hvtnfet l=6e-08 w=4e-07 $X=8175 $Y=45897 $D=616
M309 14 t_tm_preb_n vss vss hvtnfet l=6e-08 w=2.5e-07 $X=8180 $Y=17720 $D=616
M310 vss 108 ddqb vss hvtnfet l=7e-08 w=3.2e-07 $X=8250 $Y=33798 $D=616
M311 108 116 366 vss hvtnfet l=1.4e-07 w=7.5e-07 $X=8290 $Y=34593 $D=616
M312 vss 11 114 vss hvtnfet l=6e-08 w=4e-07 $X=8435 $Y=4836 $D=616
M313 vss b_mb<0> 587 vss hvtnfet l=6e-08 w=4e-07 $X=8435 $Y=11331 $D=616
M314 vss 13 588 vss hvtnfet l=6e-08 w=4e-07 $X=8435 $Y=12191 $D=616
M315 vss 14 589 vss hvtnfet l=6e-08 w=4e-07 $X=8435 $Y=38542 $D=616
M316 vss t_mb<0> 590 vss hvtnfet l=6e-08 w=4e-07 $X=8435 $Y=39402 $D=616
M317 vss 11 115 vss hvtnfet l=6e-08 w=4e-07 $X=8435 $Y=45897 $D=616
M318 vss t_tm_preb_n 14 vss hvtnfet l=6e-08 w=2.5e-07 $X=8440 $Y=17720 $D=616
M319 vss saeb_n 117 vss hvtnfet l=6e-08 w=3e-07 $X=8507 $Y=31223 $D=616
M320 366 117 vss vss hvtnfet l=8e-08 w=3.75e-07 $X=8530 $Y=33798 $D=616
M321 140 clk_dqb vss vss hvtnfet l=6e-08 w=2e-07 $X=8615 $Y=21427 $D=616
M322 138 clk_dqb_n vss vss hvtnfet l=6e-08 w=2e-07 $X=8615 $Y=23694 $D=616
M323 122 121 vss vss hvtnfet l=6e-08 w=2e-07 $X=8615 $Y=24394 $D=616
M324 148 122 vss vss hvtnfet l=6e-08 w=2e-07 $X=8615 $Y=24904 $D=616
M325 366 116 108 vss hvtnfet l=1.4e-07 w=7.5e-07 $X=8630 $Y=34593 $D=616
M326 195 126 vss vss hvtnfet l=6e-08 w=6e-07 $X=8647 $Y=26159 $D=616
M327 124 20 vss vss hvtnfet l=6e-08 w=4e-07 $X=8695 $Y=4836 $D=616
M328 591 b_ma<0> vss vss hvtnfet l=6e-08 w=4e-07 $X=8695 $Y=11331 $D=616
M329 592 22 vss vss hvtnfet l=6e-08 w=4e-07 $X=8695 $Y=12191 $D=616
M330 593 23 vss vss hvtnfet l=6e-08 w=4e-07 $X=8695 $Y=38542 $D=616
M331 594 t_ma<0> vss vss hvtnfet l=6e-08 w=4e-07 $X=8695 $Y=39402 $D=616
M332 125 20 vss vss hvtnfet l=6e-08 w=4e-07 $X=8695 $Y=45897 $D=616
M333 13 b_tm_preb_n vss vss hvtnfet l=6e-08 w=2.5e-07 $X=8700 $Y=17720 $D=616
M334 213 114 b_blb_n<3> vss hvtnfet l=6e-08 w=6e-07 $X=8740 $Y=2941 $D=616
M335 213 114 b_blb_n<3> vss hvtnfet l=6e-08 w=6e-07 $X=8740 $Y=3201 $D=616
M336 b_bla<3> 124 224 vss hvtnfet l=6e-08 w=6e-07 $X=8740 $Y=3881 $D=616
M337 b_bla<3> 124 224 vss hvtnfet l=6e-08 w=6e-07 $X=8740 $Y=4141 $D=616
M338 224 125 t_bla<3> vss hvtnfet l=6e-08 w=6e-07 $X=8740 $Y=46932 $D=616
M339 t_bla<3> 125 224 vss hvtnfet l=6e-08 w=6e-07 $X=8740 $Y=47192 $D=616
M340 t_blb_n<3> 115 213 vss hvtnfet l=6e-08 w=6e-07 $X=8740 $Y=47872 $D=616
M341 213 115 t_blb_n<3> vss hvtnfet l=6e-08 w=6e-07 $X=8740 $Y=48132 $D=616
M342 137 142 vss vss hvtnfet l=6e-08 w=3e-07 $X=8767 $Y=31223 $D=616
M343 vss 117 366 vss hvtnfet l=8e-08 w=3.75e-07 $X=8810 $Y=33798 $D=616
M344 vss 126 195 vss hvtnfet l=6e-08 w=6e-07 $X=8907 $Y=26159 $D=616
M345 vss 127 124 vss hvtnfet l=6e-08 w=4e-07 $X=8955 $Y=4836 $D=616
M346 127 b_ca<3> 591 vss hvtnfet l=6e-08 w=4e-07 $X=8955 $Y=11331 $D=616
M347 132 127 592 vss hvtnfet l=6e-08 w=4e-07 $X=8955 $Y=12191 $D=616
M348 133 128 593 vss hvtnfet l=6e-08 w=4e-07 $X=8955 $Y=38542 $D=616
M349 128 t_ca<3> 594 vss hvtnfet l=6e-08 w=4e-07 $X=8955 $Y=39402 $D=616
M350 vss 128 125 vss hvtnfet l=6e-08 w=4e-07 $X=8955 $Y=45897 $D=616
M351 vss b_tm_preb_n 13 vss hvtnfet l=6e-08 w=2.5e-07 $X=8960 $Y=17720 $D=616
M352 116 108 366 vss hvtnfet l=1.4e-07 w=7.5e-07 $X=8970 $Y=34593 $D=616
M353 366 117 vss vss hvtnfet l=8e-08 w=3.75e-07 $X=9090 $Y=33798 $D=616
M354 366 108 116 vss hvtnfet l=1.4e-07 w=7.5e-07 $X=9310 $Y=34593 $D=616
M355 vss 117 366 vss hvtnfet l=8e-08 w=3.75e-07 $X=9370 $Y=33798 $D=616
M356 qb 137 vss vss hvtnfet l=6e-08 w=4.5e-07 $X=9395 $Y=19812 $D=616
M357 vss 137 qb vss hvtnfet l=6e-08 w=4.5e-07 $X=9395 $Y=20072 $D=616
M358 11 lweb 354 vss hvtnfet l=6e-08 w=8e-07 $X=9427 $Y=26159 $D=616
M359 vss 139 150 vss hvtnfet l=1.4e-07 w=2.1e-07 $X=9445 $Y=14555 $D=616
M360 vss db 143 vss hvtnfet l=1.4e-07 w=2.1e-07 $X=9445 $Y=16755 $D=616
M361 359 vdd vss vss hvtnfet l=6e-08 w=3e-07 $X=9470 $Y=17670 $D=616
M362 595 149 vss vss hvtnfet l=6e-08 w=3.2e-07 $X=9525 $Y=21012 $D=616
M363 595 140 126 vss hvtnfet l=6e-08 w=3.2e-07 $X=9525 $Y=21202 $D=616
M364 vss 126 156 vss hvtnfet l=6e-08 w=3.2e-07 $X=9525 $Y=22762 $D=616
M365 596 150 vss vss hvtnfet l=6e-08 w=3.2e-07 $X=9525 $Y=23729 $D=616
M366 596 140 121 vss hvtnfet l=6e-08 w=3.2e-07 $X=9525 $Y=23919 $D=616
M367 165 126 vss vss hvtnfet l=6e-08 w=2.1e-07 $X=9635 $Y=21942 $D=616
M368 166 121 vss vss hvtnfet l=6e-08 w=2.1e-07 $X=9635 $Y=24659 $D=616
M369 366 117 vss vss hvtnfet l=8e-08 w=3.75e-07 $X=9650 $Y=33798 $D=616
M370 108 116 366 vss hvtnfet l=1.4e-07 w=7.5e-07 $X=9650 $Y=34593 $D=616
M371 599 saeb_n vss vss hvtnfet l=6e-08 w=3e-07 $X=9677 $Y=31223 $D=616
M372 354 lweb 11 vss hvtnfet l=6e-08 w=8e-07 $X=9687 $Y=26159 $D=616
M373 597 165 126 vss hvtnfet l=6e-08 w=1.4e-07 $X=9705 $Y=21477 $D=616
M374 vss 138 597 vss hvtnfet l=6e-08 w=1.4e-07 $X=9705 $Y=21667 $D=616
M375 598 166 121 vss hvtnfet l=6e-08 w=1.4e-07 $X=9705 $Y=24194 $D=616
M376 vss 138 598 vss hvtnfet l=6e-08 w=1.4e-07 $X=9705 $Y=24384 $D=616
M377 vss vdd 359 vss hvtnfet l=6e-08 w=3e-07 $X=9730 $Y=17670 $D=616
M378 213 159 b_blb_n<2> vss hvtnfet l=6e-08 w=6e-07 $X=9760 $Y=2941 $D=616
M379 213 159 b_blb_n<2> vss hvtnfet l=6e-08 w=6e-07 $X=9760 $Y=3201 $D=616
M380 b_bla<2> 153 224 vss hvtnfet l=6e-08 w=6e-07 $X=9760 $Y=3881 $D=616
M381 b_bla<2> 153 224 vss hvtnfet l=6e-08 w=6e-07 $X=9760 $Y=4141 $D=616
M382 224 154 t_bla<2> vss hvtnfet l=6e-08 w=6e-07 $X=9760 $Y=46932 $D=616
M383 t_bla<2> 154 224 vss hvtnfet l=6e-08 w=6e-07 $X=9760 $Y=47192 $D=616
M384 t_blb_n<2> 160 213 vss hvtnfet l=6e-08 w=6e-07 $X=9760 $Y=47872 $D=616
M385 213 160 t_blb_n<2> vss hvtnfet l=6e-08 w=6e-07 $X=9760 $Y=48132 $D=616
M386 139 152 vss vss hvtnfet l=1.4e-07 w=2.1e-07 $X=9785 $Y=14555 $D=616
M387 151 143 vss vss hvtnfet l=1.4e-07 w=2.1e-07 $X=9785 $Y=16755 $D=616
M388 142 137 599 vss hvtnfet l=6e-08 w=3e-07 $X=9867 $Y=31223 $D=616
M389 vss 117 366 vss hvtnfet l=8e-08 w=3.75e-07 $X=9930 $Y=33798 $D=616
M390 vss 148 354 vss hvtnfet l=6e-08 w=8e-07 $X=9947 $Y=26159 $D=616
M391 359 vdd vss vss hvtnfet l=6e-08 w=3e-07 $X=9990 $Y=17670 $D=616
M392 366 116 108 vss hvtnfet l=1.4e-07 w=7.5e-07 $X=9990 $Y=34593 $D=616
M393 153 144 vss vss hvtnfet l=6e-08 w=4e-07 $X=10085 $Y=4836 $D=616
M394 600 b_ca<2> 144 vss hvtnfet l=6e-08 w=4e-07 $X=10085 $Y=11331 $D=616
M395 601 144 146 vss hvtnfet l=6e-08 w=4e-07 $X=10085 $Y=12191 $D=616
M396 602 145 147 vss hvtnfet l=6e-08 w=4e-07 $X=10085 $Y=38542 $D=616
M397 603 t_ca<2> 145 vss hvtnfet l=6e-08 w=4e-07 $X=10085 $Y=39402 $D=616
M398 154 145 vss vss hvtnfet l=6e-08 w=4e-07 $X=10085 $Y=45897 $D=616
M399 604 116 142 vss hvtnfet l=6e-08 w=3e-07 $X=10127 $Y=31223 $D=616
M400 354 148 vss vss hvtnfet l=6e-08 w=8e-07 $X=10207 $Y=26159 $D=616
M401 366 117 vss vss hvtnfet l=8e-08 w=3.75e-07 $X=10210 $Y=33798 $D=616
M402 vss vdd 359 vss hvtnfet l=6e-08 w=3e-07 $X=10250 $Y=17670 $D=616
M403 vss 117 604 vss hvtnfet l=6e-08 w=3e-07 $X=10317 $Y=31223 $D=616
M404 116 108 366 vss hvtnfet l=1.4e-07 w=7.5e-07 $X=10330 $Y=34593 $D=616
M405 vss 20 153 vss hvtnfet l=6e-08 w=4e-07 $X=10345 $Y=4836 $D=616
M406 vss b_ma<0> 600 vss hvtnfet l=6e-08 w=4e-07 $X=10345 $Y=11331 $D=616
M407 vss 22 601 vss hvtnfet l=6e-08 w=4e-07 $X=10345 $Y=12191 $D=616
M408 vss 23 602 vss hvtnfet l=6e-08 w=4e-07 $X=10345 $Y=38542 $D=616
M409 vss t_ma<0> 603 vss hvtnfet l=6e-08 w=4e-07 $X=10345 $Y=39402 $D=616
M410 vss 20 154 vss hvtnfet l=6e-08 w=4e-07 $X=10345 $Y=45897 $D=616
M411 vss 155 152 vss hvtnfet l=1.4e-07 w=2.1e-07 $X=10375 $Y=14555 $D=616
M412 vss 151 164 vss hvtnfet l=1.4e-07 w=2.1e-07 $X=10375 $Y=16755 $D=616
M413 vss 117 366 vss hvtnfet l=8e-08 w=3.75e-07 $X=10490 $Y=33798 $D=616
M414 359 vdd vss vss hvtnfet l=6e-08 w=3e-07 $X=10510 $Y=17670 $D=616
M415 159 11 vss vss hvtnfet l=6e-08 w=4e-07 $X=10605 $Y=4836 $D=616
M416 605 b_mb<0> vss vss hvtnfet l=6e-08 w=4e-07 $X=10605 $Y=11331 $D=616
M417 606 13 vss vss hvtnfet l=6e-08 w=4e-07 $X=10605 $Y=12191 $D=616
M418 607 14 vss vss hvtnfet l=6e-08 w=4e-07 $X=10605 $Y=38542 $D=616
M419 608 t_mb<0> vss vss hvtnfet l=6e-08 w=4e-07 $X=10605 $Y=39402 $D=616
M420 160 11 vss vss hvtnfet l=6e-08 w=4e-07 $X=10605 $Y=45897 $D=616
M421 195 159 b_blb<2> vss hvtnfet l=6e-08 w=6e-07 $X=10650 $Y=2941 $D=616
M422 195 159 b_blb<2> vss hvtnfet l=6e-08 w=6e-07 $X=10650 $Y=3201 $D=616
M423 204 153 b_bla_n<2> vss hvtnfet l=6e-08 w=6e-07 $X=10650 $Y=3881 $D=616
M424 204 153 b_bla_n<2> vss hvtnfet l=6e-08 w=6e-07 $X=10650 $Y=4141 $D=616
M425 t_bla_n<2> 154 204 vss hvtnfet l=6e-08 w=6e-07 $X=10650 $Y=46932 $D=616
M426 204 154 t_bla_n<2> vss hvtnfet l=6e-08 w=6e-07 $X=10650 $Y=47192 $D=616
M427 t_blb<2> 160 195 vss hvtnfet l=6e-08 w=6e-07 $X=10650 $Y=47872 $D=616
M428 195 160 t_blb<2> vss hvtnfet l=6e-08 w=6e-07 $X=10650 $Y=48132 $D=616
M429 366 108 116 vss hvtnfet l=1.4e-07 w=7.5e-07 $X=10670 $Y=34593 $D=616
M430 155 bwenb vss vss hvtnfet l=1.4e-07 w=2.1e-07 $X=10715 $Y=14555 $D=616
M431 149 164 vss vss hvtnfet l=1.4e-07 w=2.1e-07 $X=10715 $Y=16755 $D=616
M432 213 156 vss vss hvtnfet l=6e-08 w=6e-07 $X=10717 $Y=26159 $D=616
M433 vss vdd 359 vss hvtnfet l=6e-08 w=3e-07 $X=10770 $Y=17670 $D=616
M434 ddqb_n 116 vss vss hvtnfet l=7e-08 w=3.2e-07 $X=10780 $Y=33798 $D=616
M435 370 vdd vss vss hvtnfet l=6e-08 w=3e-07 $X=10827 $Y=31223 $D=616
M436 vss 157 159 vss hvtnfet l=6e-08 w=4e-07 $X=10865 $Y=4836 $D=616
M437 157 b_cb<2> 605 vss hvtnfet l=6e-08 w=4e-07 $X=10865 $Y=11331 $D=616
M438 162 157 606 vss hvtnfet l=6e-08 w=4e-07 $X=10865 $Y=12191 $D=616
M439 163 158 607 vss hvtnfet l=6e-08 w=4e-07 $X=10865 $Y=38542 $D=616
M440 158 t_cb<2> 608 vss hvtnfet l=6e-08 w=4e-07 $X=10865 $Y=39402 $D=616
M441 vss 158 160 vss hvtnfet l=6e-08 w=4e-07 $X=10865 $Y=45897 $D=616
M442 vss 156 213 vss hvtnfet l=6e-08 w=6e-07 $X=10977 $Y=26159 $D=616
M443 195 171 b_blb<1> vss hvtnfet l=6e-08 w=6e-07 $X=11670 $Y=2941 $D=616
M444 195 171 b_blb<1> vss hvtnfet l=6e-08 w=6e-07 $X=11670 $Y=3201 $D=616
M445 204 173 b_bla_n<1> vss hvtnfet l=6e-08 w=6e-07 $X=11670 $Y=3881 $D=616
M446 204 173 b_bla_n<1> vss hvtnfet l=6e-08 w=6e-07 $X=11670 $Y=4141 $D=616
M447 t_bla_n<1> 174 204 vss hvtnfet l=6e-08 w=6e-07 $X=11670 $Y=46932 $D=616
M448 204 174 t_bla_n<1> vss hvtnfet l=6e-08 w=6e-07 $X=11670 $Y=47192 $D=616
M449 t_blb<1> 172 195 vss hvtnfet l=6e-08 w=6e-07 $X=11670 $Y=47872 $D=616
M450 195 172 t_blb<1> vss hvtnfet l=6e-08 w=6e-07 $X=11670 $Y=48132 $D=616
M451 381 vdd vss vss hvtnfet l=6e-08 w=6e-07 $X=11883 $Y=26159 $D=616
M452 171 169 vss vss hvtnfet l=6e-08 w=4e-07 $X=11995 $Y=4836 $D=616
M453 609 b_cb<1> 169 vss hvtnfet l=6e-08 w=4e-07 $X=11995 $Y=11331 $D=616
M454 610 169 167 vss hvtnfet l=6e-08 w=4e-07 $X=11995 $Y=12191 $D=616
M455 611 170 168 vss hvtnfet l=6e-08 w=4e-07 $X=11995 $Y=38542 $D=616
M456 612 t_cb<1> 170 vss hvtnfet l=6e-08 w=4e-07 $X=11995 $Y=39402 $D=616
M457 172 170 vss vss hvtnfet l=6e-08 w=4e-07 $X=11995 $Y=45897 $D=616
M458 384 vdd vss vss hvtnfet l=1.4e-07 w=2.1e-07 $X=12065 $Y=14550 $D=616
M459 385 vdd vss vss hvtnfet l=1.4e-07 w=2.1e-07 $X=12065 $Y=16760 $D=616
M460 vss vss vss vss hvtnfet l=7e-08 w=3.2e-07 $X=12070 $Y=33798 $D=616
M461 402 vdd vss vss hvtnfet l=6e-08 w=3e-07 $X=12090 $Y=17670 $D=616
M462 vss vss vss vss hvtnfet l=1.4e-07 w=7.5e-07 $X=12110 $Y=34593 $D=616
M463 vss vdd 381 vss hvtnfet l=6e-08 w=6e-07 $X=12143 $Y=26159 $D=616
M464 vss 11 171 vss hvtnfet l=6e-08 w=4e-07 $X=12255 $Y=4836 $D=616
M465 vss b_mb<0> 609 vss hvtnfet l=6e-08 w=4e-07 $X=12255 $Y=11331 $D=616
M466 vss 13 610 vss hvtnfet l=6e-08 w=4e-07 $X=12255 $Y=12191 $D=616
M467 vss 14 611 vss hvtnfet l=6e-08 w=4e-07 $X=12255 $Y=38542 $D=616
M468 vss t_mb<0> 612 vss hvtnfet l=6e-08 w=4e-07 $X=12255 $Y=39402 $D=616
M469 vss 11 172 vss hvtnfet l=6e-08 w=4e-07 $X=12255 $Y=45897 $D=616
M470 vss vdd 402 vss hvtnfet l=6e-08 w=3e-07 $X=12350 $Y=17670 $D=616
M471 vss vss vss vss hvtnfet l=8e-08 w=3.75e-07 $X=12350 $Y=33798 $D=616
M472 vss vss vss vss hvtnfet l=6e-08 w=3e-07 $X=12403 $Y=31223 $D=616
M473 vss vdd 384 vss hvtnfet l=1.4e-07 w=2.1e-07 $X=12405 $Y=14550 $D=616
M474 vss vdd 385 vss hvtnfet l=1.4e-07 w=2.1e-07 $X=12405 $Y=16760 $D=616
M475 vss vss vss vss hvtnfet l=1.4e-07 w=7.5e-07 $X=12450 $Y=34593 $D=616
M476 173 20 vss vss hvtnfet l=6e-08 w=4e-07 $X=12515 $Y=4836 $D=616
M477 613 b_ma<0> vss vss hvtnfet l=6e-08 w=4e-07 $X=12515 $Y=11331 $D=616
M478 614 22 vss vss hvtnfet l=6e-08 w=4e-07 $X=12515 $Y=12191 $D=616
M479 615 23 vss vss hvtnfet l=6e-08 w=4e-07 $X=12515 $Y=38542 $D=616
M480 616 t_ma<0> vss vss hvtnfet l=6e-08 w=4e-07 $X=12515 $Y=39402 $D=616
M481 174 20 vss vss hvtnfet l=6e-08 w=4e-07 $X=12515 $Y=45897 $D=616
M482 213 171 b_blb_n<1> vss hvtnfet l=6e-08 w=6e-07 $X=12560 $Y=2941 $D=616
M483 213 171 b_blb_n<1> vss hvtnfet l=6e-08 w=6e-07 $X=12560 $Y=3201 $D=616
M484 b_bla<1> 173 224 vss hvtnfet l=6e-08 w=6e-07 $X=12560 $Y=3881 $D=616
M485 b_bla<1> 173 224 vss hvtnfet l=6e-08 w=6e-07 $X=12560 $Y=4141 $D=616
M486 224 174 t_bla<1> vss hvtnfet l=6e-08 w=6e-07 $X=12560 $Y=46932 $D=616
M487 t_bla<1> 174 224 vss hvtnfet l=6e-08 w=6e-07 $X=12560 $Y=47192 $D=616
M488 t_blb_n<1> 172 213 vss hvtnfet l=6e-08 w=6e-07 $X=12560 $Y=47872 $D=616
M489 213 172 t_blb_n<1> vss hvtnfet l=6e-08 w=6e-07 $X=12560 $Y=48132 $D=616
M490 402 vdd vss vss hvtnfet l=6e-08 w=3e-07 $X=12610 $Y=17670 $D=616
M491 vss vss vss vss hvtnfet l=8e-08 w=3.75e-07 $X=12630 $Y=33798 $D=616
M492 vss vdd 408 vss hvtnfet l=6e-08 w=8e-07 $X=12653 $Y=26159 $D=616
M493 vss vss vss vss hvtnfet l=6e-08 w=3e-07 $X=12663 $Y=31223 $D=616
M494 vss 175 173 vss hvtnfet l=6e-08 w=4e-07 $X=12775 $Y=4836 $D=616
M495 175 b_ca<1> 613 vss hvtnfet l=6e-08 w=4e-07 $X=12775 $Y=11331 $D=616
M496 177 175 614 vss hvtnfet l=6e-08 w=4e-07 $X=12775 $Y=12191 $D=616
M497 178 176 615 vss hvtnfet l=6e-08 w=4e-07 $X=12775 $Y=38542 $D=616
M498 176 t_ca<1> 616 vss hvtnfet l=6e-08 w=4e-07 $X=12775 $Y=39402 $D=616
M499 vss 176 174 vss hvtnfet l=6e-08 w=4e-07 $X=12775 $Y=45897 $D=616
M500 vss vss vss vss hvtnfet l=1.4e-07 w=7.5e-07 $X=12790 $Y=34593 $D=616
M501 vss vdd 402 vss hvtnfet l=6e-08 w=3e-07 $X=12870 $Y=17670 $D=616
M502 vss vss vss vss hvtnfet l=8e-08 w=3.75e-07 $X=12910 $Y=33798 $D=616
M503 408 vdd vss vss hvtnfet l=6e-08 w=8e-07 $X=12913 $Y=26159 $D=616
M504 vss vss vss vss hvtnfet l=6e-08 w=3e-07 $X=12923 $Y=31223 $D=616
M505 400 vdd vss vss hvtnfet l=1.4e-07 w=2.1e-07 $X=12995 $Y=14550 $D=616
M506 401 vdd vss vss hvtnfet l=1.4e-07 w=2.1e-07 $X=12995 $Y=16760 $D=616
M507 vss vss vss vss hvtnfet l=6e-08 w=3.2e-07 $X=13040 $Y=19812 $D=616
M508 vss vss vss vss hvtnfet l=6e-08 w=3.2e-07 $X=13040 $Y=20072 $D=616
M509 vss vss vss vss hvtnfet l=6e-08 w=3.2e-07 $X=13040 $Y=21162 $D=616
M510 vss vss vss vss hvtnfet l=6e-08 w=3.2e-07 $X=13040 $Y=21422 $D=616
M511 vss vss vss vss hvtnfet l=6e-08 w=3.2e-07 $X=13040 $Y=21682 $D=616
M512 vss vss vss vss hvtnfet l=6e-08 w=3.2e-07 $X=13040 $Y=21942 $D=616
M513 vss vss vss vss hvtnfet l=6e-08 w=3.2e-07 $X=13040 $Y=22762 $D=616
M514 vss vss vss vss hvtnfet l=6e-08 w=3.2e-07 $X=13040 $Y=23879 $D=616
M515 vss vss vss vss hvtnfet l=6e-08 w=3.2e-07 $X=13040 $Y=24139 $D=616
M516 vss vss vss vss hvtnfet l=6e-08 w=3.2e-07 $X=13040 $Y=24399 $D=616
M517 vss vss vss vss hvtnfet l=6e-08 w=3.2e-07 $X=13040 $Y=24659 $D=616
M518 402 vdd vss vss hvtnfet l=6e-08 w=3e-07 $X=13130 $Y=17670 $D=616
M519 vss vss vss vss hvtnfet l=1.4e-07 w=7.5e-07 $X=13130 $Y=34593 $D=616
M520 403 vdd 408 vss hvtnfet l=6e-08 w=8e-07 $X=13173 $Y=26159 $D=616
M521 vss vss vss vss hvtnfet l=6e-08 w=3e-07 $X=13183 $Y=31223 $D=616
M522 vss vss vss vss hvtnfet l=8e-08 w=3.75e-07 $X=13190 $Y=33798 $D=616
M523 vss vdd 400 vss hvtnfet l=1.4e-07 w=2.1e-07 $X=13335 $Y=14550 $D=616
M524 vss vdd 401 vss hvtnfet l=1.4e-07 w=2.1e-07 $X=13335 $Y=16760 $D=616
M525 vss vdd 402 vss hvtnfet l=6e-08 w=3e-07 $X=13390 $Y=17670 $D=616
M526 408 vdd 403 vss hvtnfet l=6e-08 w=8e-07 $X=13433 $Y=26159 $D=616
M527 vss vss vss vss hvtnfet l=8e-08 w=3.75e-07 $X=13470 $Y=33798 $D=616
M528 vss vss vss vss hvtnfet l=1.4e-07 w=7.5e-07 $X=13470 $Y=34593 $D=616
M529 213 187 b_blb_n<0> vss hvtnfet l=6e-08 w=6e-07 $X=13580 $Y=2941 $D=616
M530 213 187 b_blb_n<0> vss hvtnfet l=6e-08 w=6e-07 $X=13580 $Y=3201 $D=616
M531 b_bla<0> 183 224 vss hvtnfet l=6e-08 w=6e-07 $X=13580 $Y=3881 $D=616
M532 b_bla<0> 183 224 vss hvtnfet l=6e-08 w=6e-07 $X=13580 $Y=4141 $D=616
M533 224 184 t_bla<0> vss hvtnfet l=6e-08 w=6e-07 $X=13580 $Y=46932 $D=616
M534 t_bla<0> 184 224 vss hvtnfet l=6e-08 w=6e-07 $X=13580 $Y=47192 $D=616
M535 t_blb_n<0> 188 213 vss hvtnfet l=6e-08 w=6e-07 $X=13580 $Y=47872 $D=616
M536 213 188 t_blb_n<0> vss hvtnfet l=6e-08 w=6e-07 $X=13580 $Y=48132 $D=616
M537 vss vss vss vss hvtnfet l=8e-08 w=3.75e-07 $X=13750 $Y=33798 $D=616
M538 vss vss vss vss hvtnfet l=1.4e-07 w=7.5e-07 $X=13810 $Y=34593 $D=616
M539 426 vdd vss vss hvtnfet l=6e-08 w=2.5e-07 $X=13900 $Y=17720 $D=616
M540 183 179 vss vss hvtnfet l=6e-08 w=4e-07 $X=13905 $Y=4836 $D=616
M541 617 b_ca<0> 179 vss hvtnfet l=6e-08 w=4e-07 $X=13905 $Y=11331 $D=616
M542 618 179 181 vss hvtnfet l=6e-08 w=4e-07 $X=13905 $Y=12191 $D=616
M543 619 180 182 vss hvtnfet l=6e-08 w=4e-07 $X=13905 $Y=38542 $D=616
M544 620 t_ca<0> 180 vss hvtnfet l=6e-08 w=4e-07 $X=13905 $Y=39402 $D=616
M545 184 180 vss vss hvtnfet l=6e-08 w=4e-07 $X=13905 $Y=45897 $D=616
M546 415 vdd vss vss hvtnfet l=6e-08 w=6e-07 $X=13953 $Y=26159 $D=616
M547 vss vss vss vss hvtnfet l=8e-08 w=3.75e-07 $X=14030 $Y=33798 $D=616
M548 vss vss vss vss hvtnfet l=6e-08 w=3e-07 $X=14093 $Y=31223 $D=616
M549 416 vdd vss vss hvtnfet l=6e-08 w=2e-07 $X=14105 $Y=21427 $D=616
M550 417 vdd vss vss hvtnfet l=6e-08 w=2e-07 $X=14105 $Y=23694 $D=616
M551 418 vdd vss vss hvtnfet l=6e-08 w=2e-07 $X=14105 $Y=24394 $D=616
M552 419 vdd vss vss hvtnfet l=6e-08 w=2e-07 $X=14105 $Y=24904 $D=616
M553 vss vss vss vss hvtnfet l=1.4e-07 w=7.5e-07 $X=14150 $Y=34593 $D=616
M554 vss vdd 426 vss hvtnfet l=6e-08 w=2.5e-07 $X=14160 $Y=17720 $D=616
M555 vss 20 183 vss hvtnfet l=6e-08 w=4e-07 $X=14165 $Y=4836 $D=616
M556 vss b_ma<0> 617 vss hvtnfet l=6e-08 w=4e-07 $X=14165 $Y=11331 $D=616
M557 vss 22 618 vss hvtnfet l=6e-08 w=4e-07 $X=14165 $Y=12191 $D=616
M558 vss 23 619 vss hvtnfet l=6e-08 w=4e-07 $X=14165 $Y=38542 $D=616
M559 vss t_ma<0> 620 vss hvtnfet l=6e-08 w=4e-07 $X=14165 $Y=39402 $D=616
M560 vss 20 184 vss hvtnfet l=6e-08 w=4e-07 $X=14165 $Y=45897 $D=616
M561 vss vdd 415 vss hvtnfet l=6e-08 w=6e-07 $X=14213 $Y=26159 $D=616
M562 vss vss vss vss hvtnfet l=8e-08 w=3.75e-07 $X=14310 $Y=33798 $D=616
M563 vss vss vss vss hvtnfet l=6e-08 w=3e-07 $X=14353 $Y=31223 $D=616
M564 426 vdd vss vss hvtnfet l=6e-08 w=2.5e-07 $X=14420 $Y=17720 $D=616
M565 187 11 vss vss hvtnfet l=6e-08 w=4e-07 $X=14425 $Y=4836 $D=616
M566 621 b_mb<0> vss vss hvtnfet l=6e-08 w=4e-07 $X=14425 $Y=11331 $D=616
M567 622 13 vss vss hvtnfet l=6e-08 w=4e-07 $X=14425 $Y=12191 $D=616
M568 623 14 vss vss hvtnfet l=6e-08 w=4e-07 $X=14425 $Y=38542 $D=616
M569 624 t_mb<0> vss vss hvtnfet l=6e-08 w=4e-07 $X=14425 $Y=39402 $D=616
M570 188 11 vss vss hvtnfet l=6e-08 w=4e-07 $X=14425 $Y=45897 $D=616
M571 195 187 b_blb<0> vss hvtnfet l=6e-08 w=6e-07 $X=14470 $Y=2941 $D=616
M572 195 187 b_blb<0> vss hvtnfet l=6e-08 w=6e-07 $X=14470 $Y=3201 $D=616
M573 204 183 b_bla_n<0> vss hvtnfet l=6e-08 w=6e-07 $X=14470 $Y=3881 $D=616
M574 204 183 b_bla_n<0> vss hvtnfet l=6e-08 w=6e-07 $X=14470 $Y=4141 $D=616
M575 t_bla_n<0> 184 204 vss hvtnfet l=6e-08 w=6e-07 $X=14470 $Y=46932 $D=616
M576 204 184 t_bla_n<0> vss hvtnfet l=6e-08 w=6e-07 $X=14470 $Y=47192 $D=616
M577 t_blb<0> 188 195 vss hvtnfet l=6e-08 w=6e-07 $X=14470 $Y=47872 $D=616
M578 195 188 t_blb<0> vss hvtnfet l=6e-08 w=6e-07 $X=14470 $Y=48132 $D=616
M579 vss vss vss vss hvtnfet l=1.4e-07 w=7.5e-07 $X=14490 $Y=34593 $D=616
M580 vss vss vss vss hvtnfet l=7e-08 w=3.2e-07 $X=14600 $Y=33798 $D=616
M581 vss vdd 426 vss hvtnfet l=6e-08 w=2.5e-07 $X=14680 $Y=17720 $D=616
M582 vss 185 187 vss hvtnfet l=6e-08 w=4e-07 $X=14685 $Y=4836 $D=616
M583 185 b_cb<0> 621 vss hvtnfet l=6e-08 w=4e-07 $X=14685 $Y=11331 $D=616
M584 189 185 622 vss hvtnfet l=6e-08 w=4e-07 $X=14685 $Y=12191 $D=616
M585 190 186 623 vss hvtnfet l=6e-08 w=4e-07 $X=14685 $Y=38542 $D=616
M586 186 t_cb<0> 624 vss hvtnfet l=6e-08 w=4e-07 $X=14685 $Y=39402 $D=616
M587 vss 186 188 vss hvtnfet l=6e-08 w=4e-07 $X=14685 $Y=45897 $D=616
M588 b_blb_n<7> 2 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=187 $Y=-170 $D=636
M589 t_blb_n<7> 3 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=187 $Y=50503 $D=636
M590 vdd vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=205 $Y=35893 $D=636
M591 192 5 b_blb<7> vdd hvtpfet l=6e-08 w=3e-07 $X=210 $Y=1094 $D=636
M592 b_blb<7> 5 192 vdd hvtpfet l=6e-08 w=3e-07 $X=210 $Y=1354 $D=636
M593 b_blb_n<7> 5 193 vdd hvtpfet l=6e-08 w=3e-07 $X=210 $Y=1864 $D=636
M594 193 5 b_blb_n<7> vdd hvtpfet l=6e-08 w=3e-07 $X=210 $Y=2124 $D=636
M595 t_blb_n<7> 6 193 vdd hvtpfet l=6e-08 w=3e-07 $X=210 $Y=48949 $D=636
M596 193 6 t_blb_n<7> vdd hvtpfet l=6e-08 w=3e-07 $X=210 $Y=49209 $D=636
M597 192 6 t_blb<7> vdd hvtpfet l=6e-08 w=3e-07 $X=210 $Y=49719 $D=636
M598 t_blb<7> 6 192 vdd hvtpfet l=6e-08 w=3e-07 $X=210 $Y=49979 $D=636
M599 198 vdd vdd vdd hvtpfet l=6e-08 w=4e-07 $X=255 $Y=21427 $D=636
M600 199 vdd vdd vdd hvtpfet l=6e-08 w=4e-07 $X=255 $Y=23694 $D=636
M601 200 vdd vdd vdd hvtpfet l=6e-08 w=4e-07 $X=255 $Y=24394 $D=636
M602 201 vdd vdd vdd hvtpfet l=6e-08 w=4e-07 $X=255 $Y=24904 $D=636
M603 b_blb<7> 2 b_blb_n<7> vdd hvtpfet l=6e-08 w=8e-07 $X=447 $Y=-170 $D=636
M604 t_blb<7> 3 t_blb_n<7> vdd hvtpfet l=6e-08 w=8e-07 $X=447 $Y=50503 $D=636
M605 629 5 8 vdd hvtpfet l=6e-08 w=8e-07 $X=535 $Y=5556 $D=636
M606 5 b_cb<3> vdd vdd hvtpfet l=6e-08 w=4e-07 $X=535 $Y=10611 $D=636
M607 2 5 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=535 $Y=12911 $D=636
M608 3 6 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=535 $Y=37822 $D=636
M609 6 t_cb<3> vdd vdd hvtpfet l=6e-08 w=4e-07 $X=535 $Y=40122 $D=636
M610 630 6 9 vdd hvtpfet l=6e-08 w=8e-07 $X=535 $Y=44777 $D=636
M611 215 vdd vdd vdd hvtpfet l=6e-08 w=5e-07 $X=540 $Y=18290 $D=636
M612 vdd vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=650 $Y=35893 $D=636
M613 vdd vdd vdd vdd hvtpfet l=1e-07 w=2e-07 $X=685 $Y=36723 $D=636
M614 vdd 2 b_blb<7> vdd hvtpfet l=6e-08 w=8e-07 $X=707 $Y=-170 $D=636
M615 vdd 3 t_blb<7> vdd hvtpfet l=6e-08 w=8e-07 $X=707 $Y=50503 $D=636
M616 vdd 11 629 vdd hvtpfet l=6e-08 w=8e-07 $X=795 $Y=5556 $D=636
M617 vdd b_mb<1> 5 vdd hvtpfet l=6e-08 w=4e-07 $X=795 $Y=10611 $D=636
M618 vdd 13 2 vdd hvtpfet l=6e-08 w=4e-07 $X=795 $Y=12911 $D=636
M619 vdd 14 3 vdd hvtpfet l=6e-08 w=4e-07 $X=795 $Y=37822 $D=636
M620 vdd t_mb<1> 6 vdd hvtpfet l=6e-08 w=4e-07 $X=795 $Y=40122 $D=636
M621 vdd 11 630 vdd hvtpfet l=6e-08 w=8e-07 $X=795 $Y=44777 $D=636
M622 vdd vdd 215 vdd hvtpfet l=6e-08 w=5e-07 $X=800 $Y=18290 $D=636
M623 vdd vdd vdd vdd hvtpfet l=6e-08 w=6e-07 $X=867 $Y=29008 $D=636
M624 vdd vdd vdd vdd hvtpfet l=1e-07 w=2e-07 $X=985 $Y=36723 $D=636
M625 vdd vdd vdd vdd hvtpfet l=7e-08 w=3.2e-07 $X=990 $Y=32628 $D=636
M626 vdd vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=990 $Y=35893 $D=636
M627 631 20 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=1055 $Y=5556 $D=636
M628 18 b_ma<1> vdd vdd hvtpfet l=6e-08 w=4e-07 $X=1055 $Y=10611 $D=636
M629 25 22 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=1055 $Y=12911 $D=636
M630 26 23 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=1055 $Y=37822 $D=636
M631 19 t_ma<1> vdd vdd hvtpfet l=6e-08 w=4e-07 $X=1055 $Y=40122 $D=636
M632 632 20 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=1055 $Y=44777 $D=636
M633 215 vdd vdd vdd hvtpfet l=6e-08 w=5e-07 $X=1060 $Y=18290 $D=636
M634 vdd vdd vdd vdd hvtpfet l=6e-08 w=6e-07 $X=1127 $Y=29008 $D=636
M635 b_bla_n<7> 25 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=1143 $Y=-170 $D=636
M636 t_bla_n<7> 26 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=1143 $Y=50503 $D=636
M637 vdd vdd 214 vdd hvtpfet l=6e-08 w=6e-07 $X=1267 $Y=27488 $D=636
M638 vdd vdd vdd vdd hvtpfet l=7e-08 w=3.2e-07 $X=1280 $Y=32628 $D=636
M639 vdd vdd vdd vdd hvtpfet l=1e-07 w=2e-07 $X=1285 $Y=36723 $D=636
M640 16 18 631 vdd hvtpfet l=6e-08 w=8e-07 $X=1315 $Y=5556 $D=636
M641 vdd b_ca<3> 18 vdd hvtpfet l=6e-08 w=4e-07 $X=1315 $Y=10611 $D=636
M642 vdd 18 25 vdd hvtpfet l=6e-08 w=4e-07 $X=1315 $Y=12911 $D=636
M643 vdd 19 26 vdd hvtpfet l=6e-08 w=4e-07 $X=1315 $Y=37822 $D=636
M644 vdd t_ca<3> 19 vdd hvtpfet l=6e-08 w=4e-07 $X=1315 $Y=40122 $D=636
M645 17 19 632 vdd hvtpfet l=6e-08 w=8e-07 $X=1315 $Y=44777 $D=636
M646 vdd vdd 215 vdd hvtpfet l=6e-08 w=5e-07 $X=1320 $Y=18290 $D=636
M647 vdd vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=1330 $Y=35893 $D=636
M648 221 18 b_bla<7> vdd hvtpfet l=6e-08 w=3e-07 $X=1400 $Y=1094 $D=636
M649 b_bla<7> 18 221 vdd hvtpfet l=6e-08 w=3e-07 $X=1400 $Y=1354 $D=636
M650 b_bla_n<7> 18 222 vdd hvtpfet l=6e-08 w=3e-07 $X=1400 $Y=1864 $D=636
M651 222 18 b_bla_n<7> vdd hvtpfet l=6e-08 w=3e-07 $X=1400 $Y=2124 $D=636
M652 t_bla_n<7> 19 222 vdd hvtpfet l=6e-08 w=3e-07 $X=1400 $Y=48949 $D=636
M653 222 19 t_bla_n<7> vdd hvtpfet l=6e-08 w=3e-07 $X=1400 $Y=49209 $D=636
M654 221 19 t_bla<7> vdd hvtpfet l=6e-08 w=3e-07 $X=1400 $Y=49719 $D=636
M655 t_bla<7> 19 221 vdd hvtpfet l=6e-08 w=3e-07 $X=1400 $Y=49979 $D=636
M656 b_bla<7> 25 b_bla_n<7> vdd hvtpfet l=6e-08 w=8e-07 $X=1403 $Y=-170 $D=636
M657 t_bla<7> 26 t_bla_n<7> vdd hvtpfet l=6e-08 w=8e-07 $X=1403 $Y=50503 $D=636
M658 vdd vdd vdd vdd hvtpfet l=1e-07 w=6e-07 $X=1560 $Y=32628 $D=636
M659 vdd vdd vdd vdd hvtpfet l=1e-07 w=2e-07 $X=1585 $Y=36723 $D=636
M660 vdd 25 b_bla<7> vdd hvtpfet l=6e-08 w=8e-07 $X=1663 $Y=-170 $D=636
M661 vdd 26 t_bla<7> vdd hvtpfet l=6e-08 w=8e-07 $X=1663 $Y=50503 $D=636
M662 vdd vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=1670 $Y=35893 $D=636
M663 239 vdd vdd vdd hvtpfet l=6e-08 w=8e-07 $X=1787 $Y=27288 $D=636
M664 233 vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=1805 $Y=15090 $D=636
M665 234 vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=1805 $Y=16110 $D=636
M666 249 vdd vdd vdd hvtpfet l=6e-08 w=6e-07 $X=1830 $Y=18290 $D=636
M667 vdd vdd vdd vdd hvtpfet l=1e-07 w=6e-07 $X=1860 $Y=32628 $D=636
M668 vdd vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=2010 $Y=35893 $D=636
M669 vdd vdd vdd vdd hvtpfet l=6e-08 w=6e-07 $X=2037 $Y=29008 $D=636
M670 vdd vdd 239 vdd hvtpfet l=6e-08 w=8e-07 $X=2047 $Y=27288 $D=636
M671 vdd vdd 249 vdd hvtpfet l=6e-08 w=6e-07 $X=2090 $Y=18290 $D=636
M672 b_bla<6> 33 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=2097 $Y=-170 $D=636
M673 t_bla<6> 34 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=2097 $Y=50503 $D=636
M674 221 30 b_bla<6> vdd hvtpfet l=6e-08 w=3e-07 $X=2120 $Y=1094 $D=636
M675 b_bla<6> 30 221 vdd hvtpfet l=6e-08 w=3e-07 $X=2120 $Y=1354 $D=636
M676 b_bla_n<6> 30 222 vdd hvtpfet l=6e-08 w=3e-07 $X=2120 $Y=1864 $D=636
M677 222 30 b_bla_n<6> vdd hvtpfet l=6e-08 w=3e-07 $X=2120 $Y=2124 $D=636
M678 t_bla_n<6> 31 222 vdd hvtpfet l=6e-08 w=3e-07 $X=2120 $Y=48949 $D=636
M679 222 31 t_bla_n<6> vdd hvtpfet l=6e-08 w=3e-07 $X=2120 $Y=49209 $D=636
M680 221 31 t_bla<6> vdd hvtpfet l=6e-08 w=3e-07 $X=2120 $Y=49719 $D=636
M681 t_bla<6> 31 221 vdd hvtpfet l=6e-08 w=3e-07 $X=2120 $Y=49979 $D=636
M682 vdd vdd vdd vdd hvtpfet l=1e-07 w=2e-07 $X=2135 $Y=36723 $D=636
M683 vdd vdd 233 vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=2145 $Y=15090 $D=636
M684 vdd vdd 234 vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=2145 $Y=16110 $D=636
M685 vdd vdd vdd vdd hvtpfet l=1e-07 w=6e-07 $X=2160 $Y=32628 $D=636
M686 vdd vdd vdd vdd hvtpfet l=6e-08 w=6e-07 $X=2297 $Y=29008 $D=636
M687 239 vdd vdd vdd hvtpfet l=6e-08 w=8e-07 $X=2307 $Y=27288 $D=636
M688 249 vdd vdd vdd hvtpfet l=6e-08 w=6e-07 $X=2350 $Y=18290 $D=636
M689 vdd vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=2350 $Y=35893 $D=636
M690 b_bla_n<6> 33 b_bla<6> vdd hvtpfet l=6e-08 w=8e-07 $X=2357 $Y=-170 $D=636
M691 t_bla_n<6> 34 t_bla<6> vdd hvtpfet l=6e-08 w=8e-07 $X=2357 $Y=50503 $D=636
M692 vdd vdd vdd vdd hvtpfet l=1e-07 w=2e-07 $X=2435 $Y=36723 $D=636
M693 637 30 35 vdd hvtpfet l=6e-08 w=8e-07 $X=2445 $Y=5556 $D=636
M694 30 b_ca<2> vdd vdd hvtpfet l=6e-08 w=4e-07 $X=2445 $Y=10611 $D=636
M695 33 30 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=2445 $Y=12911 $D=636
M696 34 31 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=2445 $Y=37822 $D=636
M697 31 t_ca<2> vdd vdd hvtpfet l=6e-08 w=4e-07 $X=2445 $Y=40122 $D=636
M698 638 31 36 vdd hvtpfet l=6e-08 w=8e-07 $X=2445 $Y=44777 $D=636
M699 vdd vdd vdd vdd hvtpfet l=7e-08 w=3.2e-07 $X=2470 $Y=32628 $D=636
M700 vdd vdd vdd vdd hvtpfet l=6e-08 w=6e-07 $X=2557 $Y=29008 $D=636
M701 vdd vdd 239 vdd hvtpfet l=6e-08 w=8e-07 $X=2567 $Y=27288 $D=636
M702 vdd vdd 249 vdd hvtpfet l=6e-08 w=6e-07 $X=2610 $Y=18290 $D=636
M703 vdd 33 b_bla_n<6> vdd hvtpfet l=6e-08 w=8e-07 $X=2617 $Y=-170 $D=636
M704 vdd 34 t_bla_n<6> vdd hvtpfet l=6e-08 w=8e-07 $X=2617 $Y=50503 $D=636
M705 vdd vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=2690 $Y=35893 $D=636
M706 vdd 20 637 vdd hvtpfet l=6e-08 w=8e-07 $X=2705 $Y=5556 $D=636
M707 vdd b_ma<1> 30 vdd hvtpfet l=6e-08 w=4e-07 $X=2705 $Y=10611 $D=636
M708 vdd 22 33 vdd hvtpfet l=6e-08 w=4e-07 $X=2705 $Y=12911 $D=636
M709 vdd 23 34 vdd hvtpfet l=6e-08 w=4e-07 $X=2705 $Y=37822 $D=636
M710 vdd t_ma<1> 31 vdd hvtpfet l=6e-08 w=4e-07 $X=2705 $Y=40122 $D=636
M711 vdd 20 638 vdd hvtpfet l=6e-08 w=8e-07 $X=2705 $Y=44777 $D=636
M712 247 vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=2735 $Y=15090 $D=636
M713 248 vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=2735 $Y=16110 $D=636
M714 vdd vdd vdd vdd hvtpfet l=1e-07 w=2e-07 $X=2735 $Y=36723 $D=636
M715 vdd vdd vdd vdd hvtpfet l=7e-08 w=3.2e-07 $X=2760 $Y=32628 $D=636
M716 vdd vdd vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=2806 $Y=19812 $D=636
M717 vdd vdd vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=2806 $Y=20072 $D=636
M718 vdd vdd vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=2806 $Y=21162 $D=636
M719 vdd vdd vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=2806 $Y=21422 $D=636
M720 vdd vdd vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=2806 $Y=21682 $D=636
M721 vdd vdd vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=2806 $Y=21942 $D=636
M722 vdd vdd vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=2806 $Y=22762 $D=636
M723 vdd vdd vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=2806 $Y=23879 $D=636
M724 vdd vdd vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=2806 $Y=24139 $D=636
M725 vdd vdd vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=2806 $Y=24399 $D=636
M726 vdd vdd vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=2806 $Y=24659 $D=636
M727 vdd vdd vdd vdd hvtpfet l=6e-08 w=6e-07 $X=2817 $Y=29008 $D=636
M728 249 vdd vdd vdd hvtpfet l=6e-08 w=6e-07 $X=2870 $Y=18290 $D=636
M729 639 11 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=2965 $Y=5556 $D=636
M730 37 b_mb<1> vdd vdd hvtpfet l=6e-08 w=4e-07 $X=2965 $Y=10611 $D=636
M731 41 13 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=2965 $Y=12911 $D=636
M732 42 14 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=2965 $Y=37822 $D=636
M733 38 t_mb<1> vdd vdd hvtpfet l=6e-08 w=4e-07 $X=2965 $Y=40122 $D=636
M734 640 11 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=2965 $Y=44777 $D=636
M735 vdd vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=3030 $Y=35893 $D=636
M736 vdd vdd vdd vdd hvtpfet l=1e-07 w=2e-07 $X=3035 $Y=36723 $D=636
M737 b_blb<6> 41 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=3053 $Y=-170 $D=636
M738 t_blb<6> 42 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=3053 $Y=50503 $D=636
M739 vdd vdd 247 vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=3075 $Y=15090 $D=636
M740 vdd vdd 248 vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=3075 $Y=16110 $D=636
M741 256 vdd vdd vdd hvtpfet l=6e-08 w=6e-07 $X=3077 $Y=27488 $D=636
M742 vdd vdd 249 vdd hvtpfet l=6e-08 w=6e-07 $X=3130 $Y=18290 $D=636
M743 39 37 639 vdd hvtpfet l=6e-08 w=8e-07 $X=3225 $Y=5556 $D=636
M744 vdd b_cb<2> 37 vdd hvtpfet l=6e-08 w=4e-07 $X=3225 $Y=10611 $D=636
M745 vdd 37 41 vdd hvtpfet l=6e-08 w=4e-07 $X=3225 $Y=12911 $D=636
M746 vdd 38 42 vdd hvtpfet l=6e-08 w=4e-07 $X=3225 $Y=37822 $D=636
M747 vdd t_cb<2> 38 vdd hvtpfet l=6e-08 w=4e-07 $X=3225 $Y=40122 $D=636
M748 40 38 640 vdd hvtpfet l=6e-08 w=8e-07 $X=3225 $Y=44777 $D=636
M749 192 37 b_blb<6> vdd hvtpfet l=6e-08 w=3e-07 $X=3310 $Y=1094 $D=636
M750 b_blb<6> 37 192 vdd hvtpfet l=6e-08 w=3e-07 $X=3310 $Y=1354 $D=636
M751 b_blb_n<6> 37 193 vdd hvtpfet l=6e-08 w=3e-07 $X=3310 $Y=1864 $D=636
M752 193 37 b_blb_n<6> vdd hvtpfet l=6e-08 w=3e-07 $X=3310 $Y=2124 $D=636
M753 t_blb_n<6> 38 193 vdd hvtpfet l=6e-08 w=3e-07 $X=3310 $Y=48949 $D=636
M754 193 38 t_blb_n<6> vdd hvtpfet l=6e-08 w=3e-07 $X=3310 $Y=49209 $D=636
M755 192 38 t_blb<6> vdd hvtpfet l=6e-08 w=3e-07 $X=3310 $Y=49719 $D=636
M756 t_blb<6> 38 192 vdd hvtpfet l=6e-08 w=3e-07 $X=3310 $Y=49979 $D=636
M757 b_blb_n<6> 41 b_blb<6> vdd hvtpfet l=6e-08 w=8e-07 $X=3313 $Y=-170 $D=636
M758 t_blb_n<6> 42 t_blb<6> vdd hvtpfet l=6e-08 w=8e-07 $X=3313 $Y=50503 $D=636
M759 vdd vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=3475 $Y=35893 $D=636
M760 vdd 41 b_blb_n<6> vdd hvtpfet l=6e-08 w=8e-07 $X=3573 $Y=-170 $D=636
M761 vdd 42 t_blb_n<6> vdd hvtpfet l=6e-08 w=8e-07 $X=3573 $Y=50503 $D=636
M762 b_blb_n<5> 45 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=4007 $Y=-170 $D=636
M763 t_blb_n<5> 46 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=4007 $Y=50503 $D=636
M764 vdd vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=4025 $Y=35893 $D=636
M765 192 48 b_blb<5> vdd hvtpfet l=6e-08 w=3e-07 $X=4030 $Y=1094 $D=636
M766 b_blb<5> 48 192 vdd hvtpfet l=6e-08 w=3e-07 $X=4030 $Y=1354 $D=636
M767 b_blb_n<5> 48 193 vdd hvtpfet l=6e-08 w=3e-07 $X=4030 $Y=1864 $D=636
M768 193 48 b_blb_n<5> vdd hvtpfet l=6e-08 w=3e-07 $X=4030 $Y=2124 $D=636
M769 t_blb_n<5> 49 193 vdd hvtpfet l=6e-08 w=3e-07 $X=4030 $Y=48949 $D=636
M770 193 49 t_blb_n<5> vdd hvtpfet l=6e-08 w=3e-07 $X=4030 $Y=49209 $D=636
M771 192 49 t_blb<5> vdd hvtpfet l=6e-08 w=3e-07 $X=4030 $Y=49719 $D=636
M772 t_blb<5> 49 192 vdd hvtpfet l=6e-08 w=3e-07 $X=4030 $Y=49979 $D=636
M773 qa 67 vdd vdd hvtpfet l=6e-08 w=9e-07 $X=4118 $Y=19812 $D=636
M774 qa 67 vdd vdd hvtpfet l=6e-08 w=9e-07 $X=4118 $Y=20072 $D=636
M775 b_blb<5> 45 b_blb_n<5> vdd hvtpfet l=6e-08 w=8e-07 $X=4267 $Y=-170 $D=636
M776 t_blb<5> 46 t_blb_n<5> vdd hvtpfet l=6e-08 w=8e-07 $X=4267 $Y=50503 $D=636
M777 645 48 54 vdd hvtpfet l=6e-08 w=8e-07 $X=4355 $Y=5556 $D=636
M778 48 b_cb<1> vdd vdd hvtpfet l=6e-08 w=4e-07 $X=4355 $Y=10611 $D=636
M779 45 48 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=4355 $Y=12911 $D=636
M780 46 49 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=4355 $Y=37822 $D=636
M781 49 t_cb<1> vdd vdd hvtpfet l=6e-08 w=4e-07 $X=4355 $Y=40122 $D=636
M782 646 49 55 vdd hvtpfet l=6e-08 w=8e-07 $X=4355 $Y=44777 $D=636
M783 vdd vdd 270 vdd hvtpfet l=6e-08 w=6e-07 $X=4393 $Y=29008 $D=636
M784 vdd bwena 64 vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=4425 $Y=15085 $D=636
M785 vdd 56 76 vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=4425 $Y=16115 $D=636
M786 288 vdd vdd vdd hvtpfet l=6e-08 w=6e-07 $X=4450 $Y=18290 $D=636
M787 57 59 vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=4470 $Y=35893 $D=636
M788 647 76 vdd vdd hvtpfet l=6e-08 w=4.8e-07 $X=4473 $Y=21012 $D=636
M789 647 51 73 vdd hvtpfet l=6e-08 w=4.8e-07 $X=4473 $Y=21202 $D=636
M790 61 73 vdd vdd hvtpfet l=6e-08 w=4.8e-07 $X=4473 $Y=22762 $D=636
M791 648 77 vdd vdd hvtpfet l=6e-08 w=4.8e-07 $X=4473 $Y=23729 $D=636
M792 648 51 74 vdd hvtpfet l=6e-08 w=4.8e-07 $X=4473 $Y=23919 $D=636
M793 vdd 61 204 vdd hvtpfet l=6e-08 w=6e-07 $X=4503 $Y=27488 $D=636
M794 57 60 221 vdd hvtpfet l=1e-07 w=2e-07 $X=4505 $Y=36723 $D=636
M795 vdd 45 b_blb<5> vdd hvtpfet l=6e-08 w=8e-07 $X=4527 $Y=-170 $D=636
M796 vdd 46 t_blb<5> vdd hvtpfet l=6e-08 w=8e-07 $X=4527 $Y=50503 $D=636
M797 vdd 11 645 vdd hvtpfet l=6e-08 w=8e-07 $X=4615 $Y=5556 $D=636
M798 vdd b_mb<1> 48 vdd hvtpfet l=6e-08 w=4e-07 $X=4615 $Y=10611 $D=636
M799 vdd 13 45 vdd hvtpfet l=6e-08 w=4e-07 $X=4615 $Y=12911 $D=636
M800 vdd 14 46 vdd hvtpfet l=6e-08 w=4e-07 $X=4615 $Y=37822 $D=636
M801 vdd t_mb<1> 49 vdd hvtpfet l=6e-08 w=4e-07 $X=4615 $Y=40122 $D=636
M802 vdd 11 646 vdd hvtpfet l=6e-08 w=8e-07 $X=4615 $Y=44777 $D=636
M803 vdd 73 53 vdd hvtpfet l=6e-08 w=3.2e-07 $X=4633 $Y=21942 $D=636
M804 vdd 74 52 vdd hvtpfet l=6e-08 w=3.2e-07 $X=4633 $Y=24659 $D=636
M805 vdd vdd 288 vdd hvtpfet l=6e-08 w=6e-07 $X=4710 $Y=18290 $D=636
M806 649 53 73 vdd hvtpfet l=6e-08 w=2.1e-07 $X=4743 $Y=21477 $D=636
M807 649 71 vdd vdd hvtpfet l=6e-08 w=2.1e-07 $X=4743 $Y=21667 $D=636
M808 650 52 74 vdd hvtpfet l=6e-08 w=2.1e-07 $X=4743 $Y=24194 $D=636
M809 650 71 vdd vdd hvtpfet l=6e-08 w=2.1e-07 $X=4743 $Y=24384 $D=636
M810 72 64 vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=4765 $Y=15085 $D=636
M811 56 75 vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=4765 $Y=16115 $D=636
M812 221 60 57 vdd hvtpfet l=1e-07 w=2e-07 $X=4805 $Y=36723 $D=636
M813 ddqa_n 57 vdd vdd hvtpfet l=7e-08 w=3.2e-07 $X=4810 $Y=32628 $D=636
M814 vdd 59 57 vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=4810 $Y=35893 $D=636
M815 651 20 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=4875 $Y=5556 $D=636
M816 65 b_ma<1> vdd vdd hvtpfet l=6e-08 w=4e-07 $X=4875 $Y=10611 $D=636
M817 69 22 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=4875 $Y=12911 $D=636
M818 70 23 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=4875 $Y=37822 $D=636
M819 66 t_ma<1> vdd vdd hvtpfet l=6e-08 w=4e-07 $X=4875 $Y=40122 $D=636
M820 652 20 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=4875 $Y=44777 $D=636
M821 653 60 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=4903 $Y=29008 $D=636
M822 b_bla_n<5> 69 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=4963 $Y=-170 $D=636
M823 t_bla_n<5> 70 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=4963 $Y=50503 $D=636
M824 288 vdd vdd vdd hvtpfet l=6e-08 w=6e-07 $X=4970 $Y=18290 $D=636
M825 20 68 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=5013 $Y=27288 $D=636
M826 82 67 653 vdd hvtpfet l=6e-08 w=6e-07 $X=5093 $Y=29008 $D=636
M827 vdd 57 ddqa_n vdd hvtpfet l=7e-08 w=3.2e-07 $X=5100 $Y=32628 $D=636
M828 57 60 221 vdd hvtpfet l=1e-07 w=2e-07 $X=5105 $Y=36723 $D=636
M829 62 65 651 vdd hvtpfet l=6e-08 w=8e-07 $X=5135 $Y=5556 $D=636
M830 vdd b_ca<1> 65 vdd hvtpfet l=6e-08 w=4e-07 $X=5135 $Y=10611 $D=636
M831 vdd 65 69 vdd hvtpfet l=6e-08 w=4e-07 $X=5135 $Y=12911 $D=636
M832 vdd 66 70 vdd hvtpfet l=6e-08 w=4e-07 $X=5135 $Y=37822 $D=636
M833 vdd t_ca<1> 66 vdd hvtpfet l=6e-08 w=4e-07 $X=5135 $Y=40122 $D=636
M834 63 66 652 vdd hvtpfet l=6e-08 w=8e-07 $X=5135 $Y=44777 $D=636
M835 59 57 vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=5150 $Y=35893 $D=636
M836 221 65 b_bla<5> vdd hvtpfet l=6e-08 w=3e-07 $X=5220 $Y=1094 $D=636
M837 b_bla<5> 65 221 vdd hvtpfet l=6e-08 w=3e-07 $X=5220 $Y=1354 $D=636
M838 b_bla_n<5> 65 222 vdd hvtpfet l=6e-08 w=3e-07 $X=5220 $Y=1864 $D=636
M839 222 65 b_bla_n<5> vdd hvtpfet l=6e-08 w=3e-07 $X=5220 $Y=2124 $D=636
M840 t_bla_n<5> 66 222 vdd hvtpfet l=6e-08 w=3e-07 $X=5220 $Y=48949 $D=636
M841 222 66 t_bla_n<5> vdd hvtpfet l=6e-08 w=3e-07 $X=5220 $Y=49209 $D=636
M842 221 66 t_bla<5> vdd hvtpfet l=6e-08 w=3e-07 $X=5220 $Y=49719 $D=636
M843 t_bla<5> 66 221 vdd hvtpfet l=6e-08 w=3e-07 $X=5220 $Y=49979 $D=636
M844 b_bla<5> 69 b_bla_n<5> vdd hvtpfet l=6e-08 w=8e-07 $X=5223 $Y=-170 $D=636
M845 t_bla<5> 70 t_bla_n<5> vdd hvtpfet l=6e-08 w=8e-07 $X=5223 $Y=50503 $D=636
M846 vdd vdd 288 vdd hvtpfet l=6e-08 w=6e-07 $X=5230 $Y=18290 $D=636
M847 vdd 68 20 vdd hvtpfet l=6e-08 w=8e-07 $X=5273 $Y=27288 $D=636
M848 654 57 82 vdd hvtpfet l=6e-08 w=6e-07 $X=5353 $Y=29008 $D=636
M849 vdd 72 85 vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=5355 $Y=15085 $D=636
M850 vdd 80 75 vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=5355 $Y=16115 $D=636
M851 57 sa_prea_n vdd vdd hvtpfet l=1e-07 w=6e-07 $X=5380 $Y=32628 $D=636
M852 221 60 57 vdd hvtpfet l=1e-07 w=2e-07 $X=5405 $Y=36723 $D=636
M853 vdd 69 b_bla<5> vdd hvtpfet l=6e-08 w=8e-07 $X=5483 $Y=-170 $D=636
M854 vdd 70 t_bla<5> vdd hvtpfet l=6e-08 w=8e-07 $X=5483 $Y=50503 $D=636
M855 288 vdd vdd vdd hvtpfet l=6e-08 w=6e-07 $X=5490 $Y=18290 $D=636
M856 vdd 57 59 vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=5490 $Y=35893 $D=636
M857 20 lwea vdd vdd hvtpfet l=6e-08 w=8e-07 $X=5533 $Y=27288 $D=636
M858 vdd saea_n 654 vdd hvtpfet l=6e-08 w=6e-07 $X=5543 $Y=29008 $D=636
M859 59 sa_prea_n 57 vdd hvtpfet l=1e-07 w=6e-07 $X=5680 $Y=32628 $D=636
M860 77 85 vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=5695 $Y=15085 $D=636
M861 80 da vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=5695 $Y=16115 $D=636
M862 vdd vdd 288 vdd hvtpfet l=6e-08 w=6e-07 $X=5750 $Y=18290 $D=636
M863 vdd lwea 20 vdd hvtpfet l=6e-08 w=8e-07 $X=5793 $Y=27288 $D=636
M864 57 59 vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=5830 $Y=35893 $D=636
M865 b_bla<4> 91 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=5917 $Y=-170 $D=636
M866 t_bla<4> 92 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=5917 $Y=50503 $D=636
M867 221 88 b_bla<4> vdd hvtpfet l=6e-08 w=3e-07 $X=5940 $Y=1094 $D=636
M868 b_bla<4> 88 221 vdd hvtpfet l=6e-08 w=3e-07 $X=5940 $Y=1354 $D=636
M869 b_bla_n<4> 88 222 vdd hvtpfet l=6e-08 w=3e-07 $X=5940 $Y=1864 $D=636
M870 222 88 b_bla_n<4> vdd hvtpfet l=6e-08 w=3e-07 $X=5940 $Y=2124 $D=636
M871 t_bla_n<4> 89 222 vdd hvtpfet l=6e-08 w=3e-07 $X=5940 $Y=48949 $D=636
M872 222 89 t_bla_n<4> vdd hvtpfet l=6e-08 w=3e-07 $X=5940 $Y=49209 $D=636
M873 221 89 t_bla<4> vdd hvtpfet l=6e-08 w=3e-07 $X=5940 $Y=49719 $D=636
M874 t_bla<4> 89 221 vdd hvtpfet l=6e-08 w=3e-07 $X=5940 $Y=49979 $D=636
M875 59 60 222 vdd hvtpfet l=1e-07 w=2e-07 $X=5955 $Y=36723 $D=636
M876 vdd sa_prea_n 59 vdd hvtpfet l=1e-07 w=6e-07 $X=5980 $Y=32628 $D=636
M877 vdd 59 57 vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=6170 $Y=35893 $D=636
M878 b_bla_n<4> 91 b_bla<4> vdd hvtpfet l=6e-08 w=8e-07 $X=6177 $Y=-170 $D=636
M879 t_bla_n<4> 92 t_bla<4> vdd hvtpfet l=6e-08 w=8e-07 $X=6177 $Y=50503 $D=636
M880 222 60 59 vdd hvtpfet l=1e-07 w=2e-07 $X=6255 $Y=36723 $D=636
M881 22 b_tm_prea_n vdd vdd hvtpfet l=6e-08 w=5e-07 $X=6260 $Y=18290 $D=636
M882 659 88 94 vdd hvtpfet l=6e-08 w=8e-07 $X=6265 $Y=5556 $D=636
M883 88 b_ca<0> vdd vdd hvtpfet l=6e-08 w=4e-07 $X=6265 $Y=10611 $D=636
M884 91 88 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=6265 $Y=12911 $D=636
M885 92 89 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=6265 $Y=37822 $D=636
M886 89 t_ca<0> vdd vdd hvtpfet l=6e-08 w=4e-07 $X=6265 $Y=40122 $D=636
M887 660 89 95 vdd hvtpfet l=6e-08 w=8e-07 $X=6265 $Y=44777 $D=636
M888 ddqa 59 vdd vdd hvtpfet l=7e-08 w=3.2e-07 $X=6290 $Y=32628 $D=636
M889 224 73 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=6313 $Y=27488 $D=636
M890 vdd 91 b_bla_n<4> vdd hvtpfet l=6e-08 w=8e-07 $X=6437 $Y=-170 $D=636
M891 vdd 92 t_bla_n<4> vdd hvtpfet l=6e-08 w=8e-07 $X=6437 $Y=50503 $D=636
M892 vdd 82 67 vdd hvtpfet l=6e-08 w=6e-07 $X=6453 $Y=29008 $D=636
M893 59 57 vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=6510 $Y=35893 $D=636
M894 vdd b_tm_prea_n 22 vdd hvtpfet l=6e-08 w=5e-07 $X=6520 $Y=18290 $D=636
M895 vdd 20 659 vdd hvtpfet l=6e-08 w=8e-07 $X=6525 $Y=5556 $D=636
M896 vdd b_ma<1> 88 vdd hvtpfet l=6e-08 w=4e-07 $X=6525 $Y=10611 $D=636
M897 vdd 22 91 vdd hvtpfet l=6e-08 w=4e-07 $X=6525 $Y=12911 $D=636
M898 vdd 23 92 vdd hvtpfet l=6e-08 w=4e-07 $X=6525 $Y=37822 $D=636
M899 vdd t_ma<1> 89 vdd hvtpfet l=6e-08 w=4e-07 $X=6525 $Y=40122 $D=636
M900 vdd 20 660 vdd hvtpfet l=6e-08 w=8e-07 $X=6525 $Y=44777 $D=636
M901 59 60 222 vdd hvtpfet l=1e-07 w=2e-07 $X=6555 $Y=36723 $D=636
M902 vdd 59 ddqa vdd hvtpfet l=7e-08 w=3.2e-07 $X=6580 $Y=32628 $D=636
M903 60 saea_n vdd vdd hvtpfet l=6e-08 w=6e-07 $X=6713 $Y=29008 $D=636
M904 23 t_tm_prea_n vdd vdd hvtpfet l=6e-08 w=5e-07 $X=6780 $Y=18290 $D=636
M905 661 11 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=6785 $Y=5556 $D=636
M906 99 b_mb<1> vdd vdd hvtpfet l=6e-08 w=4e-07 $X=6785 $Y=10611 $D=636
M907 103 13 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=6785 $Y=12911 $D=636
M908 104 14 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=6785 $Y=37822 $D=636
M909 100 t_mb<1> vdd vdd hvtpfet l=6e-08 w=4e-07 $X=6785 $Y=40122 $D=636
M910 662 11 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=6785 $Y=44777 $D=636
M911 vdd 57 59 vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=6850 $Y=35893 $D=636
M912 222 60 59 vdd hvtpfet l=1e-07 w=2e-07 $X=6855 $Y=36723 $D=636
M913 b_blb<4> 103 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=6873 $Y=-170 $D=636
M914 t_blb<4> 104 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=6873 $Y=50503 $D=636
M915 71 clk_dqa vdd vdd hvtpfet l=6e-08 w=4e-07 $X=6985 $Y=21427 $D=636
M916 51 clk_dqa_n vdd vdd hvtpfet l=6e-08 w=4e-07 $X=6985 $Y=23694 $D=636
M917 98 74 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=6985 $Y=24394 $D=636
M918 68 98 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=6985 $Y=24904 $D=636
M919 vdd t_tm_prea_n 23 vdd hvtpfet l=6e-08 w=5e-07 $X=7040 $Y=18290 $D=636
M920 101 99 661 vdd hvtpfet l=6e-08 w=8e-07 $X=7045 $Y=5556 $D=636
M921 vdd b_cb<0> 99 vdd hvtpfet l=6e-08 w=4e-07 $X=7045 $Y=10611 $D=636
M922 vdd 99 103 vdd hvtpfet l=6e-08 w=4e-07 $X=7045 $Y=12911 $D=636
M923 vdd 100 104 vdd hvtpfet l=6e-08 w=4e-07 $X=7045 $Y=37822 $D=636
M924 vdd t_cb<0> 100 vdd hvtpfet l=6e-08 w=4e-07 $X=7045 $Y=40122 $D=636
M925 102 100 662 vdd hvtpfet l=6e-08 w=8e-07 $X=7045 $Y=44777 $D=636
M926 192 99 b_blb<4> vdd hvtpfet l=6e-08 w=3e-07 $X=7130 $Y=1094 $D=636
M927 b_blb<4> 99 192 vdd hvtpfet l=6e-08 w=3e-07 $X=7130 $Y=1354 $D=636
M928 b_blb_n<4> 99 193 vdd hvtpfet l=6e-08 w=3e-07 $X=7130 $Y=1864 $D=636
M929 193 99 b_blb_n<4> vdd hvtpfet l=6e-08 w=3e-07 $X=7130 $Y=2124 $D=636
M930 t_blb_n<4> 100 193 vdd hvtpfet l=6e-08 w=3e-07 $X=7130 $Y=48949 $D=636
M931 193 100 t_blb_n<4> vdd hvtpfet l=6e-08 w=3e-07 $X=7130 $Y=49209 $D=636
M932 192 100 t_blb<4> vdd hvtpfet l=6e-08 w=3e-07 $X=7130 $Y=49719 $D=636
M933 t_blb<4> 100 192 vdd hvtpfet l=6e-08 w=3e-07 $X=7130 $Y=49979 $D=636
M934 b_blb_n<4> 103 b_blb<4> vdd hvtpfet l=6e-08 w=8e-07 $X=7133 $Y=-170 $D=636
M935 t_blb_n<4> 104 t_blb<4> vdd hvtpfet l=6e-08 w=8e-07 $X=7133 $Y=50503 $D=636
M936 316 59 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=7223 $Y=29008 $D=636
M937 vdd vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=7295 $Y=35893 $D=636
M938 vdd 103 b_blb_n<4> vdd hvtpfet l=6e-08 w=8e-07 $X=7393 $Y=-170 $D=636
M939 vdd 104 t_blb_n<4> vdd hvtpfet l=6e-08 w=8e-07 $X=7393 $Y=50503 $D=636
M940 b_blb_n<3> 109 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=7827 $Y=-170 $D=636
M941 t_blb_n<3> 110 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=7827 $Y=50503 $D=636
M942 vdd vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=7845 $Y=35893 $D=636
M943 192 111 b_blb<3> vdd hvtpfet l=6e-08 w=3e-07 $X=7850 $Y=1094 $D=636
M944 b_blb<3> 111 192 vdd hvtpfet l=6e-08 w=3e-07 $X=7850 $Y=1354 $D=636
M945 b_blb_n<3> 111 193 vdd hvtpfet l=6e-08 w=3e-07 $X=7850 $Y=1864 $D=636
M946 193 111 b_blb_n<3> vdd hvtpfet l=6e-08 w=3e-07 $X=7850 $Y=2124 $D=636
M947 t_blb_n<3> 112 193 vdd hvtpfet l=6e-08 w=3e-07 $X=7850 $Y=48949 $D=636
M948 193 112 t_blb_n<3> vdd hvtpfet l=6e-08 w=3e-07 $X=7850 $Y=49209 $D=636
M949 192 112 t_blb<3> vdd hvtpfet l=6e-08 w=3e-07 $X=7850 $Y=49719 $D=636
M950 t_blb<3> 112 192 vdd hvtpfet l=6e-08 w=3e-07 $X=7850 $Y=49979 $D=636
M951 140 clk_dqb vdd vdd hvtpfet l=6e-08 w=4e-07 $X=7895 $Y=21427 $D=636
M952 138 clk_dqb_n vdd vdd hvtpfet l=6e-08 w=4e-07 $X=7895 $Y=23694 $D=636
M953 122 121 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=7895 $Y=24394 $D=636
M954 148 122 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=7895 $Y=24904 $D=636
M955 vdd 108 323 vdd hvtpfet l=6e-08 w=6e-07 $X=7997 $Y=29008 $D=636
M956 b_blb<3> 109 b_blb_n<3> vdd hvtpfet l=6e-08 w=8e-07 $X=8087 $Y=-170 $D=636
M957 t_blb<3> 110 t_blb_n<3> vdd hvtpfet l=6e-08 w=8e-07 $X=8087 $Y=50503 $D=636
M958 667 111 114 vdd hvtpfet l=6e-08 w=8e-07 $X=8175 $Y=5556 $D=636
M959 111 b_cb<3> vdd vdd hvtpfet l=6e-08 w=4e-07 $X=8175 $Y=10611 $D=636
M960 109 111 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=8175 $Y=12911 $D=636
M961 110 112 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=8175 $Y=37822 $D=636
M962 112 t_cb<3> vdd vdd hvtpfet l=6e-08 w=4e-07 $X=8175 $Y=40122 $D=636
M963 668 112 115 vdd hvtpfet l=6e-08 w=8e-07 $X=8175 $Y=44777 $D=636
M964 14 t_tm_preb_n vdd vdd hvtpfet l=6e-08 w=5e-07 $X=8180 $Y=18290 $D=636
M965 108 116 vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=8290 $Y=35893 $D=636
M966 108 117 193 vdd hvtpfet l=1e-07 w=2e-07 $X=8325 $Y=36723 $D=636
M967 vdd 109 b_blb<3> vdd hvtpfet l=6e-08 w=8e-07 $X=8347 $Y=-170 $D=636
M968 vdd 110 t_blb<3> vdd hvtpfet l=6e-08 w=8e-07 $X=8347 $Y=50503 $D=636
M969 vdd 11 667 vdd hvtpfet l=6e-08 w=8e-07 $X=8435 $Y=5556 $D=636
M970 vdd b_mb<0> 111 vdd hvtpfet l=6e-08 w=4e-07 $X=8435 $Y=10611 $D=636
M971 vdd 13 109 vdd hvtpfet l=6e-08 w=4e-07 $X=8435 $Y=12911 $D=636
M972 vdd 14 110 vdd hvtpfet l=6e-08 w=4e-07 $X=8435 $Y=37822 $D=636
M973 vdd t_mb<0> 112 vdd hvtpfet l=6e-08 w=4e-07 $X=8435 $Y=40122 $D=636
M974 vdd 11 668 vdd hvtpfet l=6e-08 w=8e-07 $X=8435 $Y=44777 $D=636
M975 vdd t_tm_preb_n 14 vdd hvtpfet l=6e-08 w=5e-07 $X=8440 $Y=18290 $D=636
M976 vdd saeb_n 117 vdd hvtpfet l=6e-08 w=6e-07 $X=8507 $Y=29008 $D=636
M977 193 117 108 vdd hvtpfet l=1e-07 w=2e-07 $X=8625 $Y=36723 $D=636
M978 ddqb 108 vdd vdd hvtpfet l=7e-08 w=3.2e-07 $X=8630 $Y=32628 $D=636
M979 vdd 116 108 vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=8630 $Y=35893 $D=636
M980 669 20 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=8695 $Y=5556 $D=636
M981 127 b_ma<0> vdd vdd hvtpfet l=6e-08 w=4e-07 $X=8695 $Y=10611 $D=636
M982 132 22 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=8695 $Y=12911 $D=636
M983 133 23 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=8695 $Y=37822 $D=636
M984 128 t_ma<0> vdd vdd hvtpfet l=6e-08 w=4e-07 $X=8695 $Y=40122 $D=636
M985 670 20 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=8695 $Y=44777 $D=636
M986 13 b_tm_preb_n vdd vdd hvtpfet l=6e-08 w=5e-07 $X=8700 $Y=18290 $D=636
M987 137 142 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=8767 $Y=29008 $D=636
M988 b_bla_n<3> 132 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=8783 $Y=-170 $D=636
M989 t_bla_n<3> 133 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=8783 $Y=50503 $D=636
M990 vdd 126 195 vdd hvtpfet l=6e-08 w=6e-07 $X=8907 $Y=27488 $D=636
M991 vdd 108 ddqb vdd hvtpfet l=7e-08 w=3.2e-07 $X=8920 $Y=32628 $D=636
M992 108 117 193 vdd hvtpfet l=1e-07 w=2e-07 $X=8925 $Y=36723 $D=636
M993 124 127 669 vdd hvtpfet l=6e-08 w=8e-07 $X=8955 $Y=5556 $D=636
M994 vdd b_ca<3> 127 vdd hvtpfet l=6e-08 w=4e-07 $X=8955 $Y=10611 $D=636
M995 vdd 127 132 vdd hvtpfet l=6e-08 w=4e-07 $X=8955 $Y=12911 $D=636
M996 vdd 128 133 vdd hvtpfet l=6e-08 w=4e-07 $X=8955 $Y=37822 $D=636
M997 vdd t_ca<3> 128 vdd hvtpfet l=6e-08 w=4e-07 $X=8955 $Y=40122 $D=636
M998 125 128 670 vdd hvtpfet l=6e-08 w=8e-07 $X=8955 $Y=44777 $D=636
M999 vdd b_tm_preb_n 13 vdd hvtpfet l=6e-08 w=5e-07 $X=8960 $Y=18290 $D=636
M1000 116 108 vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=8970 $Y=35893 $D=636
M1001 221 127 b_bla<3> vdd hvtpfet l=6e-08 w=3e-07 $X=9040 $Y=1094 $D=636
M1002 b_bla<3> 127 221 vdd hvtpfet l=6e-08 w=3e-07 $X=9040 $Y=1354 $D=636
M1003 b_bla_n<3> 127 222 vdd hvtpfet l=6e-08 w=3e-07 $X=9040 $Y=1864 $D=636
M1004 222 127 b_bla_n<3> vdd hvtpfet l=6e-08 w=3e-07 $X=9040 $Y=2124 $D=636
M1005 t_bla_n<3> 128 222 vdd hvtpfet l=6e-08 w=3e-07 $X=9040 $Y=48949 $D=636
M1006 222 128 t_bla_n<3> vdd hvtpfet l=6e-08 w=3e-07 $X=9040 $Y=49209 $D=636
M1007 221 128 t_bla<3> vdd hvtpfet l=6e-08 w=3e-07 $X=9040 $Y=49719 $D=636
M1008 t_bla<3> 128 221 vdd hvtpfet l=6e-08 w=3e-07 $X=9040 $Y=49979 $D=636
M1009 b_bla<3> 132 b_bla_n<3> vdd hvtpfet l=6e-08 w=8e-07 $X=9043 $Y=-170 $D=636
M1010 t_bla<3> 133 t_bla_n<3> vdd hvtpfet l=6e-08 w=8e-07 $X=9043 $Y=50503 $D=636
M1011 108 sa_preb_n vdd vdd hvtpfet l=1e-07 w=6e-07 $X=9200 $Y=32628 $D=636
M1012 193 117 108 vdd hvtpfet l=1e-07 w=2e-07 $X=9225 $Y=36723 $D=636
M1013 vdd 132 b_bla<3> vdd hvtpfet l=6e-08 w=8e-07 $X=9303 $Y=-170 $D=636
M1014 vdd 133 t_bla<3> vdd hvtpfet l=6e-08 w=8e-07 $X=9303 $Y=50503 $D=636
M1015 vdd 108 116 vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=9310 $Y=35893 $D=636
M1016 11 lweb vdd vdd hvtpfet l=6e-08 w=8e-07 $X=9427 $Y=27288 $D=636
M1017 vdd 139 150 vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=9445 $Y=15085 $D=636
M1018 vdd db 143 vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=9445 $Y=16115 $D=636
M1019 359 vdd vdd vdd hvtpfet l=6e-08 w=6e-07 $X=9470 $Y=18290 $D=636
M1020 116 sa_preb_n 108 vdd hvtpfet l=1e-07 w=6e-07 $X=9500 $Y=32628 $D=636
M1021 108 116 vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=9650 $Y=35893 $D=636
M1022 671 saeb_n vdd vdd hvtpfet l=6e-08 w=6e-07 $X=9677 $Y=29008 $D=636
M1023 vdd lweb 11 vdd hvtpfet l=6e-08 w=8e-07 $X=9687 $Y=27288 $D=636
M1024 vdd vdd 359 vdd hvtpfet l=6e-08 w=6e-07 $X=9730 $Y=18290 $D=636
M1025 b_bla<2> 146 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=9737 $Y=-170 $D=636
M1026 t_bla<2> 147 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=9737 $Y=50503 $D=636
M1027 221 144 b_bla<2> vdd hvtpfet l=6e-08 w=3e-07 $X=9760 $Y=1094 $D=636
M1028 b_bla<2> 144 221 vdd hvtpfet l=6e-08 w=3e-07 $X=9760 $Y=1354 $D=636
M1029 b_bla_n<2> 144 222 vdd hvtpfet l=6e-08 w=3e-07 $X=9760 $Y=1864 $D=636
M1030 222 144 b_bla_n<2> vdd hvtpfet l=6e-08 w=3e-07 $X=9760 $Y=2124 $D=636
M1031 t_bla_n<2> 145 222 vdd hvtpfet l=6e-08 w=3e-07 $X=9760 $Y=48949 $D=636
M1032 222 145 t_bla_n<2> vdd hvtpfet l=6e-08 w=3e-07 $X=9760 $Y=49209 $D=636
M1033 221 145 t_bla<2> vdd hvtpfet l=6e-08 w=3e-07 $X=9760 $Y=49719 $D=636
M1034 t_bla<2> 145 221 vdd hvtpfet l=6e-08 w=3e-07 $X=9760 $Y=49979 $D=636
M1035 116 117 192 vdd hvtpfet l=1e-07 w=2e-07 $X=9775 $Y=36723 $D=636
M1036 139 152 vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=9785 $Y=15085 $D=636
M1037 151 143 vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=9785 $Y=16115 $D=636
M1038 vdd sa_preb_n 116 vdd hvtpfet l=1e-07 w=6e-07 $X=9800 $Y=32628 $D=636
M1039 142 116 671 vdd hvtpfet l=6e-08 w=6e-07 $X=9867 $Y=29008 $D=636
M1040 11 148 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=9947 $Y=27288 $D=636
M1041 359 vdd vdd vdd hvtpfet l=6e-08 w=6e-07 $X=9990 $Y=18290 $D=636
M1042 vdd 116 108 vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=9990 $Y=35893 $D=636
M1043 b_bla_n<2> 146 b_bla<2> vdd hvtpfet l=6e-08 w=8e-07 $X=9997 $Y=-170 $D=636
M1044 t_bla_n<2> 147 t_bla<2> vdd hvtpfet l=6e-08 w=8e-07 $X=9997 $Y=50503 $D=636
M1045 192 117 116 vdd hvtpfet l=1e-07 w=2e-07 $X=10075 $Y=36723 $D=636
M1046 676 144 153 vdd hvtpfet l=6e-08 w=8e-07 $X=10085 $Y=5556 $D=636
M1047 144 b_ca<2> vdd vdd hvtpfet l=6e-08 w=4e-07 $X=10085 $Y=10611 $D=636
M1048 146 144 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=10085 $Y=12911 $D=636
M1049 147 145 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=10085 $Y=37822 $D=636
M1050 145 t_ca<2> vdd vdd hvtpfet l=6e-08 w=4e-07 $X=10085 $Y=40122 $D=636
M1051 677 145 154 vdd hvtpfet l=6e-08 w=8e-07 $X=10085 $Y=44777 $D=636
M1052 ddqb_n 116 vdd vdd hvtpfet l=7e-08 w=3.2e-07 $X=10110 $Y=32628 $D=636
M1053 678 137 142 vdd hvtpfet l=6e-08 w=6e-07 $X=10127 $Y=29008 $D=636
M1054 vdd 148 11 vdd hvtpfet l=6e-08 w=8e-07 $X=10207 $Y=27288 $D=636
M1055 vdd vdd 359 vdd hvtpfet l=6e-08 w=6e-07 $X=10250 $Y=18290 $D=636
M1056 vdd 146 b_bla_n<2> vdd hvtpfet l=6e-08 w=8e-07 $X=10257 $Y=-170 $D=636
M1057 vdd 147 t_bla_n<2> vdd hvtpfet l=6e-08 w=8e-07 $X=10257 $Y=50503 $D=636
M1058 qb 137 vdd vdd hvtpfet l=6e-08 w=9e-07 $X=10262 $Y=19812 $D=636
M1059 qb 137 vdd vdd hvtpfet l=6e-08 w=9e-07 $X=10262 $Y=20072 $D=636
M1060 vdd 117 678 vdd hvtpfet l=6e-08 w=6e-07 $X=10317 $Y=29008 $D=636
M1061 679 149 vdd vdd hvtpfet l=6e-08 w=4.8e-07 $X=10327 $Y=21012 $D=636
M1062 679 138 126 vdd hvtpfet l=6e-08 w=4.8e-07 $X=10327 $Y=21202 $D=636
M1063 680 165 126 vdd hvtpfet l=6e-08 w=2.1e-07 $X=10327 $Y=21477 $D=636
M1064 680 140 vdd vdd hvtpfet l=6e-08 w=2.1e-07 $X=10327 $Y=21667 $D=636
M1065 vdd 126 165 vdd hvtpfet l=6e-08 w=3.2e-07 $X=10327 $Y=21942 $D=636
M1066 156 126 vdd vdd hvtpfet l=6e-08 w=4.8e-07 $X=10327 $Y=22762 $D=636
M1067 681 150 vdd vdd hvtpfet l=6e-08 w=4.8e-07 $X=10327 $Y=23729 $D=636
M1068 681 138 121 vdd hvtpfet l=6e-08 w=4.8e-07 $X=10327 $Y=23919 $D=636
M1069 682 166 121 vdd hvtpfet l=6e-08 w=2.1e-07 $X=10327 $Y=24194 $D=636
M1070 682 140 vdd vdd hvtpfet l=6e-08 w=2.1e-07 $X=10327 $Y=24384 $D=636
M1071 vdd 121 166 vdd hvtpfet l=6e-08 w=3.2e-07 $X=10327 $Y=24659 $D=636
M1072 116 108 vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=10330 $Y=35893 $D=636
M1073 vdd 20 676 vdd hvtpfet l=6e-08 w=8e-07 $X=10345 $Y=5556 $D=636
M1074 vdd b_ma<0> 144 vdd hvtpfet l=6e-08 w=4e-07 $X=10345 $Y=10611 $D=636
M1075 vdd 22 146 vdd hvtpfet l=6e-08 w=4e-07 $X=10345 $Y=12911 $D=636
M1076 vdd 23 147 vdd hvtpfet l=6e-08 w=4e-07 $X=10345 $Y=37822 $D=636
M1077 vdd t_ma<0> 145 vdd hvtpfet l=6e-08 w=4e-07 $X=10345 $Y=40122 $D=636
M1078 vdd 20 677 vdd hvtpfet l=6e-08 w=8e-07 $X=10345 $Y=44777 $D=636
M1079 vdd 155 152 vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=10375 $Y=15085 $D=636
M1080 vdd 151 164 vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=10375 $Y=16115 $D=636
M1081 116 117 192 vdd hvtpfet l=1e-07 w=2e-07 $X=10375 $Y=36723 $D=636
M1082 vdd 116 ddqb_n vdd hvtpfet l=7e-08 w=3.2e-07 $X=10400 $Y=32628 $D=636
M1083 359 vdd vdd vdd hvtpfet l=6e-08 w=6e-07 $X=10510 $Y=18290 $D=636
M1084 683 11 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=10605 $Y=5556 $D=636
M1085 157 b_mb<0> vdd vdd hvtpfet l=6e-08 w=4e-07 $X=10605 $Y=10611 $D=636
M1086 162 13 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=10605 $Y=12911 $D=636
M1087 163 14 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=10605 $Y=37822 $D=636
M1088 158 t_mb<0> vdd vdd hvtpfet l=6e-08 w=4e-07 $X=10605 $Y=40122 $D=636
M1089 684 11 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=10605 $Y=44777 $D=636
M1090 vdd 108 116 vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=10670 $Y=35893 $D=636
M1091 192 117 116 vdd hvtpfet l=1e-07 w=2e-07 $X=10675 $Y=36723 $D=636
M1092 b_blb<2> 162 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=10693 $Y=-170 $D=636
M1093 t_blb<2> 163 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=10693 $Y=50503 $D=636
M1094 155 bwenb vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=10715 $Y=15085 $D=636
M1095 149 164 vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=10715 $Y=16115 $D=636
M1096 213 156 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=10717 $Y=27488 $D=636
M1097 vdd vdd 359 vdd hvtpfet l=6e-08 w=6e-07 $X=10770 $Y=18290 $D=636
M1098 370 vdd vdd vdd hvtpfet l=6e-08 w=6e-07 $X=10827 $Y=29008 $D=636
M1099 159 157 683 vdd hvtpfet l=6e-08 w=8e-07 $X=10865 $Y=5556 $D=636
M1100 vdd b_cb<2> 157 vdd hvtpfet l=6e-08 w=4e-07 $X=10865 $Y=10611 $D=636
M1101 vdd 157 162 vdd hvtpfet l=6e-08 w=4e-07 $X=10865 $Y=12911 $D=636
M1102 vdd 158 163 vdd hvtpfet l=6e-08 w=4e-07 $X=10865 $Y=37822 $D=636
M1103 vdd t_cb<2> 158 vdd hvtpfet l=6e-08 w=4e-07 $X=10865 $Y=40122 $D=636
M1104 160 158 684 vdd hvtpfet l=6e-08 w=8e-07 $X=10865 $Y=44777 $D=636
M1105 192 157 b_blb<2> vdd hvtpfet l=6e-08 w=3e-07 $X=10950 $Y=1094 $D=636
M1106 b_blb<2> 157 192 vdd hvtpfet l=6e-08 w=3e-07 $X=10950 $Y=1354 $D=636
M1107 b_blb_n<2> 157 193 vdd hvtpfet l=6e-08 w=3e-07 $X=10950 $Y=1864 $D=636
M1108 193 157 b_blb_n<2> vdd hvtpfet l=6e-08 w=3e-07 $X=10950 $Y=2124 $D=636
M1109 t_blb_n<2> 158 193 vdd hvtpfet l=6e-08 w=3e-07 $X=10950 $Y=48949 $D=636
M1110 193 158 t_blb_n<2> vdd hvtpfet l=6e-08 w=3e-07 $X=10950 $Y=49209 $D=636
M1111 192 158 t_blb<2> vdd hvtpfet l=6e-08 w=3e-07 $X=10950 $Y=49719 $D=636
M1112 t_blb<2> 158 192 vdd hvtpfet l=6e-08 w=3e-07 $X=10950 $Y=49979 $D=636
M1113 b_blb_n<2> 162 b_blb<2> vdd hvtpfet l=6e-08 w=8e-07 $X=10953 $Y=-170 $D=636
M1114 t_blb_n<2> 163 t_blb<2> vdd hvtpfet l=6e-08 w=8e-07 $X=10953 $Y=50503 $D=636
M1115 vdd vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=11115 $Y=35893 $D=636
M1116 vdd 162 b_blb_n<2> vdd hvtpfet l=6e-08 w=8e-07 $X=11213 $Y=-170 $D=636
M1117 vdd 163 t_blb_n<2> vdd hvtpfet l=6e-08 w=8e-07 $X=11213 $Y=50503 $D=636
M1118 b_blb_n<1> 167 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=11647 $Y=-170 $D=636
M1119 t_blb_n<1> 168 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=11647 $Y=50503 $D=636
M1120 vdd vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=11665 $Y=35893 $D=636
M1121 192 169 b_blb<1> vdd hvtpfet l=6e-08 w=3e-07 $X=11670 $Y=1094 $D=636
M1122 b_blb<1> 169 192 vdd hvtpfet l=6e-08 w=3e-07 $X=11670 $Y=1354 $D=636
M1123 b_blb_n<1> 169 193 vdd hvtpfet l=6e-08 w=3e-07 $X=11670 $Y=1864 $D=636
M1124 193 169 b_blb_n<1> vdd hvtpfet l=6e-08 w=3e-07 $X=11670 $Y=2124 $D=636
M1125 t_blb_n<1> 170 193 vdd hvtpfet l=6e-08 w=3e-07 $X=11670 $Y=48949 $D=636
M1126 193 170 t_blb_n<1> vdd hvtpfet l=6e-08 w=3e-07 $X=11670 $Y=49209 $D=636
M1127 192 170 t_blb<1> vdd hvtpfet l=6e-08 w=3e-07 $X=11670 $Y=49719 $D=636
M1128 t_blb<1> 170 192 vdd hvtpfet l=6e-08 w=3e-07 $X=11670 $Y=49979 $D=636
M1129 b_blb<1> 167 b_blb_n<1> vdd hvtpfet l=6e-08 w=8e-07 $X=11907 $Y=-170 $D=636
M1130 t_blb<1> 168 t_blb_n<1> vdd hvtpfet l=6e-08 w=8e-07 $X=11907 $Y=50503 $D=636
M1131 689 169 171 vdd hvtpfet l=6e-08 w=8e-07 $X=11995 $Y=5556 $D=636
M1132 169 b_cb<1> vdd vdd hvtpfet l=6e-08 w=4e-07 $X=11995 $Y=10611 $D=636
M1133 167 169 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=11995 $Y=12911 $D=636
M1134 168 170 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=11995 $Y=37822 $D=636
M1135 170 t_cb<1> vdd vdd hvtpfet l=6e-08 w=4e-07 $X=11995 $Y=40122 $D=636
M1136 690 170 172 vdd hvtpfet l=6e-08 w=8e-07 $X=11995 $Y=44777 $D=636
M1137 384 vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=12065 $Y=15090 $D=636
M1138 385 vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=12065 $Y=16110 $D=636
M1139 402 vdd vdd vdd hvtpfet l=6e-08 w=6e-07 $X=12090 $Y=18290 $D=636
M1140 vdd vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=12110 $Y=35893 $D=636
M1141 vdd vdd 381 vdd hvtpfet l=6e-08 w=6e-07 $X=12143 $Y=27488 $D=636
M1142 vdd vdd vdd vdd hvtpfet l=1e-07 w=2e-07 $X=12145 $Y=36723 $D=636
M1143 vdd vdd vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=12154 $Y=19812 $D=636
M1144 vdd vdd vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=12154 $Y=20072 $D=636
M1145 vdd vdd vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=12154 $Y=21162 $D=636
M1146 vdd vdd vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=12154 $Y=21422 $D=636
M1147 vdd vdd vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=12154 $Y=21682 $D=636
M1148 vdd vdd vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=12154 $Y=21942 $D=636
M1149 vdd vdd vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=12154 $Y=22762 $D=636
M1150 vdd vdd vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=12154 $Y=23879 $D=636
M1151 vdd vdd vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=12154 $Y=24139 $D=636
M1152 vdd vdd vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=12154 $Y=24399 $D=636
M1153 vdd vdd vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=12154 $Y=24659 $D=636
M1154 vdd 167 b_blb<1> vdd hvtpfet l=6e-08 w=8e-07 $X=12167 $Y=-170 $D=636
M1155 vdd 168 t_blb<1> vdd hvtpfet l=6e-08 w=8e-07 $X=12167 $Y=50503 $D=636
M1156 vdd 11 689 vdd hvtpfet l=6e-08 w=8e-07 $X=12255 $Y=5556 $D=636
M1157 vdd b_mb<0> 169 vdd hvtpfet l=6e-08 w=4e-07 $X=12255 $Y=10611 $D=636
M1158 vdd 13 167 vdd hvtpfet l=6e-08 w=4e-07 $X=12255 $Y=12911 $D=636
M1159 vdd 14 168 vdd hvtpfet l=6e-08 w=4e-07 $X=12255 $Y=37822 $D=636
M1160 vdd t_mb<0> 170 vdd hvtpfet l=6e-08 w=4e-07 $X=12255 $Y=40122 $D=636
M1161 vdd 11 690 vdd hvtpfet l=6e-08 w=8e-07 $X=12255 $Y=44777 $D=636
M1162 vdd vdd 402 vdd hvtpfet l=6e-08 w=6e-07 $X=12350 $Y=18290 $D=636
M1163 vdd vdd vdd vdd hvtpfet l=6e-08 w=6e-07 $X=12403 $Y=29008 $D=636
M1164 vdd vdd 384 vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=12405 $Y=15090 $D=636
M1165 vdd vdd 385 vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=12405 $Y=16110 $D=636
M1166 vdd vdd vdd vdd hvtpfet l=1e-07 w=2e-07 $X=12445 $Y=36723 $D=636
M1167 vdd vdd vdd vdd hvtpfet l=7e-08 w=3.2e-07 $X=12450 $Y=32628 $D=636
M1168 vdd vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=12450 $Y=35893 $D=636
M1169 691 20 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=12515 $Y=5556 $D=636
M1170 175 b_ma<0> vdd vdd hvtpfet l=6e-08 w=4e-07 $X=12515 $Y=10611 $D=636
M1171 177 22 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=12515 $Y=12911 $D=636
M1172 178 23 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=12515 $Y=37822 $D=636
M1173 176 t_ma<0> vdd vdd hvtpfet l=6e-08 w=4e-07 $X=12515 $Y=40122 $D=636
M1174 692 20 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=12515 $Y=44777 $D=636
M1175 b_bla_n<1> 177 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=12603 $Y=-170 $D=636
M1176 t_bla_n<1> 178 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=12603 $Y=50503 $D=636
M1177 402 vdd vdd vdd hvtpfet l=6e-08 w=6e-07 $X=12610 $Y=18290 $D=636
M1178 403 vdd vdd vdd hvtpfet l=6e-08 w=8e-07 $X=12653 $Y=27288 $D=636
M1179 vdd vdd vdd vdd hvtpfet l=6e-08 w=6e-07 $X=12663 $Y=29008 $D=636
M1180 vdd vdd vdd vdd hvtpfet l=7e-08 w=3.2e-07 $X=12740 $Y=32628 $D=636
M1181 vdd vdd vdd vdd hvtpfet l=1e-07 w=2e-07 $X=12745 $Y=36723 $D=636
M1182 173 175 691 vdd hvtpfet l=6e-08 w=8e-07 $X=12775 $Y=5556 $D=636
M1183 vdd b_ca<1> 175 vdd hvtpfet l=6e-08 w=4e-07 $X=12775 $Y=10611 $D=636
M1184 vdd 175 177 vdd hvtpfet l=6e-08 w=4e-07 $X=12775 $Y=12911 $D=636
M1185 vdd 176 178 vdd hvtpfet l=6e-08 w=4e-07 $X=12775 $Y=37822 $D=636
M1186 vdd t_ca<1> 176 vdd hvtpfet l=6e-08 w=4e-07 $X=12775 $Y=40122 $D=636
M1187 174 176 692 vdd hvtpfet l=6e-08 w=8e-07 $X=12775 $Y=44777 $D=636
M1188 vdd vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=12790 $Y=35893 $D=636
M1189 221 175 b_bla<1> vdd hvtpfet l=6e-08 w=3e-07 $X=12860 $Y=1094 $D=636
M1190 b_bla<1> 175 221 vdd hvtpfet l=6e-08 w=3e-07 $X=12860 $Y=1354 $D=636
M1191 b_bla_n<1> 175 222 vdd hvtpfet l=6e-08 w=3e-07 $X=12860 $Y=1864 $D=636
M1192 222 175 b_bla_n<1> vdd hvtpfet l=6e-08 w=3e-07 $X=12860 $Y=2124 $D=636
M1193 t_bla_n<1> 176 222 vdd hvtpfet l=6e-08 w=3e-07 $X=12860 $Y=48949 $D=636
M1194 222 176 t_bla_n<1> vdd hvtpfet l=6e-08 w=3e-07 $X=12860 $Y=49209 $D=636
M1195 221 176 t_bla<1> vdd hvtpfet l=6e-08 w=3e-07 $X=12860 $Y=49719 $D=636
M1196 t_bla<1> 176 221 vdd hvtpfet l=6e-08 w=3e-07 $X=12860 $Y=49979 $D=636
M1197 b_bla<1> 177 b_bla_n<1> vdd hvtpfet l=6e-08 w=8e-07 $X=12863 $Y=-170 $D=636
M1198 t_bla<1> 178 t_bla_n<1> vdd hvtpfet l=6e-08 w=8e-07 $X=12863 $Y=50503 $D=636
M1199 vdd vdd 402 vdd hvtpfet l=6e-08 w=6e-07 $X=12870 $Y=18290 $D=636
M1200 vdd vdd 403 vdd hvtpfet l=6e-08 w=8e-07 $X=12913 $Y=27288 $D=636
M1201 vdd vdd vdd vdd hvtpfet l=6e-08 w=6e-07 $X=12923 $Y=29008 $D=636
M1202 400 vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=12995 $Y=15090 $D=636
M1203 401 vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=12995 $Y=16110 $D=636
M1204 vdd vdd vdd vdd hvtpfet l=1e-07 w=6e-07 $X=13020 $Y=32628 $D=636
M1205 vdd vdd vdd vdd hvtpfet l=1e-07 w=2e-07 $X=13045 $Y=36723 $D=636
M1206 vdd 177 b_bla<1> vdd hvtpfet l=6e-08 w=8e-07 $X=13123 $Y=-170 $D=636
M1207 vdd 178 t_bla<1> vdd hvtpfet l=6e-08 w=8e-07 $X=13123 $Y=50503 $D=636
M1208 402 vdd vdd vdd hvtpfet l=6e-08 w=6e-07 $X=13130 $Y=18290 $D=636
M1209 vdd vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=13130 $Y=35893 $D=636
M1210 403 vdd vdd vdd hvtpfet l=6e-08 w=8e-07 $X=13173 $Y=27288 $D=636
M1211 vdd vdd vdd vdd hvtpfet l=6e-08 w=6e-07 $X=13183 $Y=29008 $D=636
M1212 vdd vdd vdd vdd hvtpfet l=1e-07 w=6e-07 $X=13320 $Y=32628 $D=636
M1213 vdd vdd 400 vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=13335 $Y=15090 $D=636
M1214 vdd vdd 401 vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=13335 $Y=16110 $D=636
M1215 vdd vdd 402 vdd hvtpfet l=6e-08 w=6e-07 $X=13390 $Y=18290 $D=636
M1216 vdd vdd 403 vdd hvtpfet l=6e-08 w=8e-07 $X=13433 $Y=27288 $D=636
M1217 vdd vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=13470 $Y=35893 $D=636
M1218 b_bla<0> 181 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=13557 $Y=-170 $D=636
M1219 t_bla<0> 182 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=13557 $Y=50503 $D=636
M1220 221 179 b_bla<0> vdd hvtpfet l=6e-08 w=3e-07 $X=13580 $Y=1094 $D=636
M1221 b_bla<0> 179 221 vdd hvtpfet l=6e-08 w=3e-07 $X=13580 $Y=1354 $D=636
M1222 b_bla_n<0> 179 222 vdd hvtpfet l=6e-08 w=3e-07 $X=13580 $Y=1864 $D=636
M1223 222 179 b_bla_n<0> vdd hvtpfet l=6e-08 w=3e-07 $X=13580 $Y=2124 $D=636
M1224 t_bla_n<0> 180 222 vdd hvtpfet l=6e-08 w=3e-07 $X=13580 $Y=48949 $D=636
M1225 222 180 t_bla_n<0> vdd hvtpfet l=6e-08 w=3e-07 $X=13580 $Y=49209 $D=636
M1226 221 180 t_bla<0> vdd hvtpfet l=6e-08 w=3e-07 $X=13580 $Y=49719 $D=636
M1227 t_bla<0> 180 221 vdd hvtpfet l=6e-08 w=3e-07 $X=13580 $Y=49979 $D=636
M1228 vdd vdd vdd vdd hvtpfet l=1e-07 w=2e-07 $X=13595 $Y=36723 $D=636
M1229 vdd vdd vdd vdd hvtpfet l=1e-07 w=6e-07 $X=13620 $Y=32628 $D=636
M1230 vdd vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=13810 $Y=35893 $D=636
M1231 b_bla_n<0> 181 b_bla<0> vdd hvtpfet l=6e-08 w=8e-07 $X=13817 $Y=-170 $D=636
M1232 t_bla_n<0> 182 t_bla<0> vdd hvtpfet l=6e-08 w=8e-07 $X=13817 $Y=50503 $D=636
M1233 vdd vdd vdd vdd hvtpfet l=1e-07 w=2e-07 $X=13895 $Y=36723 $D=636
M1234 426 vdd vdd vdd hvtpfet l=6e-08 w=5e-07 $X=13900 $Y=18290 $D=636
M1235 697 179 183 vdd hvtpfet l=6e-08 w=8e-07 $X=13905 $Y=5556 $D=636
M1236 179 b_ca<0> vdd vdd hvtpfet l=6e-08 w=4e-07 $X=13905 $Y=10611 $D=636
M1237 181 179 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=13905 $Y=12911 $D=636
M1238 182 180 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=13905 $Y=37822 $D=636
M1239 180 t_ca<0> vdd vdd hvtpfet l=6e-08 w=4e-07 $X=13905 $Y=40122 $D=636
M1240 698 180 184 vdd hvtpfet l=6e-08 w=8e-07 $X=13905 $Y=44777 $D=636
M1241 vdd vdd vdd vdd hvtpfet l=7e-08 w=3.2e-07 $X=13930 $Y=32628 $D=636
M1242 415 vdd vdd vdd hvtpfet l=6e-08 w=6e-07 $X=13953 $Y=27488 $D=636
M1243 vdd 181 b_bla_n<0> vdd hvtpfet l=6e-08 w=8e-07 $X=14077 $Y=-170 $D=636
M1244 vdd 182 t_bla_n<0> vdd hvtpfet l=6e-08 w=8e-07 $X=14077 $Y=50503 $D=636
M1245 vdd vdd vdd vdd hvtpfet l=6e-08 w=6e-07 $X=14093 $Y=29008 $D=636
M1246 vdd vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=14150 $Y=35893 $D=636
M1247 vdd vdd 426 vdd hvtpfet l=6e-08 w=5e-07 $X=14160 $Y=18290 $D=636
M1248 vdd 20 697 vdd hvtpfet l=6e-08 w=8e-07 $X=14165 $Y=5556 $D=636
M1249 vdd b_ma<0> 179 vdd hvtpfet l=6e-08 w=4e-07 $X=14165 $Y=10611 $D=636
M1250 vdd 22 181 vdd hvtpfet l=6e-08 w=4e-07 $X=14165 $Y=12911 $D=636
M1251 vdd 23 182 vdd hvtpfet l=6e-08 w=4e-07 $X=14165 $Y=37822 $D=636
M1252 vdd t_ma<0> 180 vdd hvtpfet l=6e-08 w=4e-07 $X=14165 $Y=40122 $D=636
M1253 vdd 20 698 vdd hvtpfet l=6e-08 w=8e-07 $X=14165 $Y=44777 $D=636
M1254 vdd vdd vdd vdd hvtpfet l=1e-07 w=2e-07 $X=14195 $Y=36723 $D=636
M1255 vdd vdd vdd vdd hvtpfet l=7e-08 w=3.2e-07 $X=14220 $Y=32628 $D=636
M1256 vdd vdd vdd vdd hvtpfet l=6e-08 w=6e-07 $X=14353 $Y=29008 $D=636
M1257 426 vdd vdd vdd hvtpfet l=6e-08 w=5e-07 $X=14420 $Y=18290 $D=636
M1258 699 11 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=14425 $Y=5556 $D=636
M1259 185 b_mb<0> vdd vdd hvtpfet l=6e-08 w=4e-07 $X=14425 $Y=10611 $D=636
M1260 189 13 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=14425 $Y=12911 $D=636
M1261 190 14 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=14425 $Y=37822 $D=636
M1262 186 t_mb<0> vdd vdd hvtpfet l=6e-08 w=4e-07 $X=14425 $Y=40122 $D=636
M1263 700 11 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=14425 $Y=44777 $D=636
M1264 vdd vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=14490 $Y=35893 $D=636
M1265 vdd vdd vdd vdd hvtpfet l=1e-07 w=2e-07 $X=14495 $Y=36723 $D=636
M1266 b_blb<0> 189 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=14513 $Y=-170 $D=636
M1267 t_blb<0> 190 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=14513 $Y=50503 $D=636
M1268 416 vdd vdd vdd hvtpfet l=6e-08 w=4e-07 $X=14625 $Y=21427 $D=636
M1269 417 vdd vdd vdd hvtpfet l=6e-08 w=4e-07 $X=14625 $Y=23694 $D=636
M1270 418 vdd vdd vdd hvtpfet l=6e-08 w=4e-07 $X=14625 $Y=24394 $D=636
M1271 419 vdd vdd vdd hvtpfet l=6e-08 w=4e-07 $X=14625 $Y=24904 $D=636
M1272 vdd vdd 426 vdd hvtpfet l=6e-08 w=5e-07 $X=14680 $Y=18290 $D=636
M1273 187 185 699 vdd hvtpfet l=6e-08 w=8e-07 $X=14685 $Y=5556 $D=636
M1274 vdd b_cb<0> 185 vdd hvtpfet l=6e-08 w=4e-07 $X=14685 $Y=10611 $D=636
M1275 vdd 185 189 vdd hvtpfet l=6e-08 w=4e-07 $X=14685 $Y=12911 $D=636
M1276 vdd 186 190 vdd hvtpfet l=6e-08 w=4e-07 $X=14685 $Y=37822 $D=636
M1277 vdd t_cb<0> 186 vdd hvtpfet l=6e-08 w=4e-07 $X=14685 $Y=40122 $D=636
M1278 188 186 700 vdd hvtpfet l=6e-08 w=8e-07 $X=14685 $Y=44777 $D=636
M1279 192 185 b_blb<0> vdd hvtpfet l=6e-08 w=3e-07 $X=14770 $Y=1094 $D=636
M1280 b_blb<0> 185 192 vdd hvtpfet l=6e-08 w=3e-07 $X=14770 $Y=1354 $D=636
M1281 b_blb_n<0> 185 193 vdd hvtpfet l=6e-08 w=3e-07 $X=14770 $Y=1864 $D=636
M1282 193 185 b_blb_n<0> vdd hvtpfet l=6e-08 w=3e-07 $X=14770 $Y=2124 $D=636
M1283 t_blb_n<0> 186 193 vdd hvtpfet l=6e-08 w=3e-07 $X=14770 $Y=48949 $D=636
M1284 193 186 t_blb_n<0> vdd hvtpfet l=6e-08 w=3e-07 $X=14770 $Y=49209 $D=636
M1285 192 186 t_blb<0> vdd hvtpfet l=6e-08 w=3e-07 $X=14770 $Y=49719 $D=636
M1286 t_blb<0> 186 192 vdd hvtpfet l=6e-08 w=3e-07 $X=14770 $Y=49979 $D=636
M1287 b_blb_n<0> 189 b_blb<0> vdd hvtpfet l=6e-08 w=8e-07 $X=14773 $Y=-170 $D=636
M1288 t_blb_n<0> 190 t_blb<0> vdd hvtpfet l=6e-08 w=8e-07 $X=14773 $Y=50503 $D=636
M1289 vdd vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=14935 $Y=35893 $D=636
M1290 vdd 189 b_blb_n<0> vdd hvtpfet l=6e-08 w=8e-07 $X=15033 $Y=-170 $D=636
M1291 vdd 190 t_blb_n<0> vdd hvtpfet l=6e-08 w=8e-07 $X=15033 $Y=50503 $D=636
.ends

************************************************************************
* Library Name: XMC55_DPS
* Cell Name:    xmc55_dps_localc8io_dummy
************************************************************************
.SUBCKT xmc55_dps_localc8io_dummy b_dbl b_dwl b_tie_low dbl_pd_n<3> 
+ dbl_pd_n<2> dbl_pd_n<1> dbl_pd_n<0> stclk t_dbl t_dwl t_tie_low vdd vss
** N=889 EP=13 IP=0 FDC=76
M0 vss 2 17 vss hvtnfet l=6e-08 w=2e-07 $X=265 $Y=2781 $D=616
M1 vss 3 18 vss hvtnfet l=6e-08 w=2e-07 $X=265 $Y=48152 $D=616
M2 28 t_dbl vss vss hvtnfet l=6e-08 w=4e-07 $X=340 $Y=26568 $D=616
M3 vss 8 stclk vss hvtnfet l=6e-08 w=3e-07 $X=340 $Y=29928 $D=616
M4 49 b_dwl vss vss hvtnfet l=6e-08 w=4e-07 $X=535 $Y=2781 $D=616
M5 50 t_dwl vss vss hvtnfet l=6e-08 w=4e-07 $X=535 $Y=47952 $D=616
M6 b_tie_low 15 vss vss hvtnfet l=7e-08 w=3.2e-07 $X=540 $Y=4916 $D=616
M7 t_tie_low 16 vss vss hvtnfet l=7e-08 w=3.2e-07 $X=540 $Y=45897 $D=616
M8 8 b_dbl 28 vss hvtnfet l=6e-08 w=4e-07 $X=600 $Y=26568 $D=616
M9 vss dbl_pd_n<2> 12 vss hvtnfet l=6e-08 w=3e-07 $X=630 $Y=19039 $D=616
M10 vss dbl_pd_n<1> 14 vss hvtnfet l=6e-08 w=3e-07 $X=630 $Y=21399 $D=616
M11 vss dbl_pd_n<0> 13 vss hvtnfet l=6e-08 w=3e-07 $X=630 $Y=22329 $D=616
M12 vss dbl_pd_n<3> 21 vss hvtnfet l=6e-08 w=3e-07 $X=630 $Y=24794 $D=616
M13 2 21 49 vss hvtnfet l=6e-08 w=4e-07 $X=795 $Y=2781 $D=616
M14 3 21 50 vss hvtnfet l=6e-08 w=4e-07 $X=795 $Y=47952 $D=616
M15 vdd vdd vdd vdd hvtpfet l=6e-08 w=8e-07 $X=187 $Y=-170 $D=636
M16 vdd vdd vdd vdd hvtpfet l=6e-08 w=8e-07 $X=187 $Y=50503 $D=636
M17 vdd 2 17 vdd hvtpfet l=6e-08 w=4e-07 $X=265 $Y=2061 $D=636
M18 vdd 3 18 vdd hvtpfet l=6e-08 w=4e-07 $X=265 $Y=48672 $D=636
M19 8 t_dbl vdd vdd hvtpfet l=6e-08 w=4e-07 $X=340 $Y=27288 $D=636
M20 vdd 8 stclk vdd hvtpfet l=6e-08 w=6e-07 $X=340 $Y=29008 $D=636
M21 b_dbl vdd vdd vdd hvtpfet l=6e-08 w=8e-07 $X=447 $Y=-170 $D=636
M22 t_dbl vdd vdd vdd hvtpfet l=6e-08 w=8e-07 $X=447 $Y=50503 $D=636
M23 2 b_dwl vdd vdd hvtpfet l=6e-08 w=4e-07 $X=535 $Y=2061 $D=636
M24 3 t_dwl vdd vdd hvtpfet l=6e-08 w=4e-07 $X=535 $Y=48672 $D=636
M25 15 15 vdd vdd hvtpfet l=7e-08 w=6.4e-07 $X=540 $Y=5556 $D=636
M26 16 16 vdd vdd hvtpfet l=7e-08 w=6.4e-07 $X=540 $Y=44937 $D=636
M27 vdd b_dbl 8 vdd hvtpfet l=6e-08 w=4e-07 $X=600 $Y=27288 $D=636
M28 vdd dbl_pd_n<2> 12 vdd hvtpfet l=6e-08 w=5e-07 $X=630 $Y=19659 $D=636
M29 vdd dbl_pd_n<1> 14 vdd hvtpfet l=6e-08 w=5e-07 $X=630 $Y=20579 $D=636
M30 vdd dbl_pd_n<0> 13 vdd hvtpfet l=6e-08 w=5e-07 $X=630 $Y=22949 $D=636
M31 vdd dbl_pd_n<3> 21 vdd hvtpfet l=6e-08 w=5e-07 $X=630 $Y=23974 $D=636
M32 vdd b_dwl b_dbl vdd hvtpfet l=6e-08 w=8e-07 $X=707 $Y=-170 $D=636
M33 vdd t_dwl t_dbl vdd hvtpfet l=6e-08 w=8e-07 $X=707 $Y=50503 $D=636
M34 vdd 21 2 vdd hvtpfet l=6e-08 w=4e-07 $X=795 $Y=2061 $D=636
M35 vdd 21 3 vdd hvtpfet l=6e-08 w=4e-07 $X=795 $Y=48672 $D=636
M36 vss t_tie_low 29 vss srpddnfet l=6e-08 w=3.15e-07 $X=670 $Y=7281 $D=778
M37 vss t_tie_low 30 vss srpddnfet l=6e-08 w=3.15e-07 $X=670 $Y=7876 $D=778
M38 vss t_tie_low 31 vss srpddnfet l=6e-08 w=3.15e-07 $X=670 $Y=9246 $D=778
M39 vss 12 32 vss srpddnfet l=6e-08 w=3.15e-07 $X=670 $Y=10871 $D=778
M40 vss 12 33 vss srpddnfet l=6e-08 w=3.15e-07 $X=670 $Y=11466 $D=778
M41 vss 12 34 vss srpddnfet l=6e-08 w=3.15e-07 $X=670 $Y=13091 $D=778
M42 vss 12 35 vss srpddnfet l=6e-08 w=3.15e-07 $X=670 $Y=13686 $D=778
M43 vss 13 36 vss srpddnfet l=6e-08 w=3.15e-07 $X=670 $Y=15311 $D=778
M44 vss 14 37 vss srpddnfet l=6e-08 w=3.15e-07 $X=670 $Y=16681 $D=778
M45 vss 14 38 vss srpddnfet l=6e-08 w=3.15e-07 $X=670 $Y=17276 $D=778
M46 vss 14 39 vss srpddnfet l=6e-08 w=3.15e-07 $X=670 $Y=33542 $D=778
M47 vss 14 40 vss srpddnfet l=6e-08 w=3.15e-07 $X=670 $Y=34137 $D=778
M48 vss 13 41 vss srpddnfet l=6e-08 w=3.15e-07 $X=670 $Y=35507 $D=778
M49 vss 12 42 vss srpddnfet l=6e-08 w=3.15e-07 $X=670 $Y=37132 $D=778
M50 vss 12 43 vss srpddnfet l=6e-08 w=3.15e-07 $X=670 $Y=37727 $D=778
M51 vss 12 44 vss srpddnfet l=6e-08 w=3.15e-07 $X=670 $Y=39352 $D=778
M52 vss 12 45 vss srpddnfet l=6e-08 w=3.15e-07 $X=670 $Y=39947 $D=778
M53 vss t_tie_low 46 vss srpddnfet l=6e-08 w=3.15e-07 $X=670 $Y=41572 $D=778
M54 vss t_tie_low 47 vss srpddnfet l=6e-08 w=3.15e-07 $X=670 $Y=42942 $D=778
M55 vss t_tie_low 48 vss srpddnfet l=6e-08 w=3.15e-07 $X=670 $Y=43537 $D=778
M56 b_dbl 17 29 vss srpgdnfet l=7.5e-08 w=1.05e-07 $X=655 $Y=6816 $D=780
M57 b_dbl 17 30 vss srpgdnfet l=7.5e-08 w=1.05e-07 $X=655 $Y=8551 $D=780
M58 b_dbl 17 31 vss srpgdnfet l=7.5e-08 w=1.05e-07 $X=655 $Y=9921 $D=780
M59 b_dbl 17 32 vss srpgdnfet l=7.5e-08 w=1.05e-07 $X=655 $Y=10406 $D=780
M60 b_dbl 17 33 vss srpgdnfet l=7.5e-08 w=1.05e-07 $X=655 $Y=12141 $D=780
M61 b_dbl 17 34 vss srpgdnfet l=7.5e-08 w=1.05e-07 $X=655 $Y=12626 $D=780
M62 b_dbl 17 35 vss srpgdnfet l=7.5e-08 w=1.05e-07 $X=655 $Y=14361 $D=780
M63 b_dbl 17 36 vss srpgdnfet l=7.5e-08 w=1.05e-07 $X=655 $Y=14846 $D=780
M64 b_dbl 17 37 vss srpgdnfet l=7.5e-08 w=1.05e-07 $X=655 $Y=16216 $D=780
M65 b_dbl 17 38 vss srpgdnfet l=7.5e-08 w=1.05e-07 $X=655 $Y=17951 $D=780
M66 t_dbl 18 39 vss srpgdnfet l=7.5e-08 w=1.05e-07 $X=655 $Y=33077 $D=780
M67 t_dbl 18 40 vss srpgdnfet l=7.5e-08 w=1.05e-07 $X=655 $Y=34812 $D=780
M68 t_dbl 18 41 vss srpgdnfet l=7.5e-08 w=1.05e-07 $X=655 $Y=36182 $D=780
M69 t_dbl 18 42 vss srpgdnfet l=7.5e-08 w=1.05e-07 $X=655 $Y=36667 $D=780
M70 t_dbl 18 43 vss srpgdnfet l=7.5e-08 w=1.05e-07 $X=655 $Y=38402 $D=780
M71 t_dbl 18 44 vss srpgdnfet l=7.5e-08 w=1.05e-07 $X=655 $Y=38887 $D=780
M72 t_dbl 18 45 vss srpgdnfet l=7.5e-08 w=1.05e-07 $X=655 $Y=40622 $D=780
M73 t_dbl 18 46 vss srpgdnfet l=7.5e-08 w=1.05e-07 $X=655 $Y=41107 $D=780
M74 t_dbl 18 47 vss srpgdnfet l=7.5e-08 w=1.05e-07 $X=655 $Y=42477 $D=780
M75 t_dbl 18 48 vss srpgdnfet l=7.5e-08 w=1.05e-07 $X=655 $Y=44212 $D=780
.ends

************************************************************************
* Library Name: XMC55_DPS
* Cell Name:    xmc55_dps_localc8io_edge
************************************************************************
.SUBCKT xmc55_dps_localc8io_edge tie_low vdd vss
** N=1093 EP=3 IP=0 FDC=59
M0 vss vss vss vss hvtnfet l=6e-08 w=4e-07 $X=970 $Y=2941 $D=616
M1 vss vss vss vss hvtnfet l=6e-08 w=4e-07 $X=970 $Y=3201 $D=616
M2 vss vss vss vss hvtnfet l=6e-08 w=4e-07 $X=970 $Y=3881 $D=616
M3 vss vss vss vss hvtnfet l=6e-08 w=4e-07 $X=970 $Y=4141 $D=616
M4 vss vss vss vss hvtnfet l=6e-08 w=4e-07 $X=970 $Y=46932 $D=616
M5 vss vss vss vss hvtnfet l=6e-08 w=4e-07 $X=970 $Y=47192 $D=616
M6 vss vss vss vss hvtnfet l=6e-08 w=4e-07 $X=970 $Y=47872 $D=616
M7 vss vss vss vss hvtnfet l=6e-08 w=4e-07 $X=970 $Y=48132 $D=616
M8 18 tie_low vss vss hvtnfet l=6e-08 w=2.1e-07 $X=1025 $Y=14555 $D=616
M9 19 tie_low vss vss hvtnfet l=6e-08 w=2.1e-07 $X=1025 $Y=16755 $D=616
M10 20 tie_low vss vss hvtnfet l=6e-08 w=2.1e-07 $X=1025 $Y=17760 $D=616
M11 5 5 vss vss hvtnfet l=6e-08 w=3.2e-07 $X=1025 $Y=26624 $D=616
M12 vss 2 tie_low vss hvtnfet l=6e-08 w=2.1e-07 $X=1025 $Y=33548 $D=616
M13 vss tie_low 10 vss hvtnfet l=6e-08 w=4e-07 $X=1130 $Y=4836 $D=616
M14 vss tie_low 11 vss hvtnfet l=6e-08 w=4e-07 $X=1130 $Y=11331 $D=616
M15 vss tie_low 12 vss hvtnfet l=6e-08 w=4e-07 $X=1130 $Y=12191 $D=616
M16 vss tie_low 13 vss hvtnfet l=6e-08 w=4e-07 $X=1130 $Y=38542 $D=616
M17 vss tie_low 14 vss hvtnfet l=6e-08 w=4e-07 $X=1130 $Y=39402 $D=616
M18 vss tie_low 15 vss hvtnfet l=6e-08 w=4e-07 $X=1130 $Y=45897 $D=616
M19 vss 5 5 vss hvtnfet l=6e-08 w=3.2e-07 $X=1285 $Y=26624 $D=616
M20 vdd vdd vdd vdd hvtpfet l=6e-08 w=3e-07 $X=975 $Y=19812 $D=636
M21 vdd vdd vdd vdd hvtpfet l=6e-08 w=3e-07 $X=975 $Y=20072 $D=636
M22 vdd vdd vdd vdd hvtpfet l=6e-08 w=3e-07 $X=975 $Y=20902 $D=636
M23 vdd vdd vdd vdd hvtpfet l=6e-08 w=3e-07 $X=975 $Y=21162 $D=636
M24 vdd vdd vdd vdd hvtpfet l=6e-08 w=3e-07 $X=975 $Y=21422 $D=636
M25 vdd vdd vdd vdd hvtpfet l=6e-08 w=3e-07 $X=975 $Y=21682 $D=636
M26 vdd vdd vdd vdd hvtpfet l=6e-08 w=3e-07 $X=975 $Y=21942 $D=636
M27 vdd vdd vdd vdd hvtpfet l=6e-08 w=3e-07 $X=975 $Y=22762 $D=636
M28 vdd vdd vdd vdd hvtpfet l=6e-08 w=3e-07 $X=975 $Y=23729 $D=636
M29 vdd vdd vdd vdd hvtpfet l=6e-08 w=3e-07 $X=975 $Y=23989 $D=636
M30 vdd vdd vdd vdd hvtpfet l=6e-08 w=3e-07 $X=975 $Y=24249 $D=636
M31 vdd vdd vdd vdd hvtpfet l=6e-08 w=3e-07 $X=975 $Y=24509 $D=636
M32 vdd vdd vdd vdd hvtpfet l=6e-08 w=3e-07 $X=975 $Y=24769 $D=636
M33 18 tie_low vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=1025 $Y=15085 $D=636
M34 19 tie_low vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=1025 $Y=16115 $D=636
M35 20 tie_low vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=1025 $Y=18290 $D=636
M36 21 5 2 vdd hvtpfet l=6e-08 w=4.8e-07 $X=1025 $Y=27313 $D=636
M37 22 5 2 vdd hvtpfet l=6e-08 w=4.8e-07 $X=1025 $Y=29008 $D=636
M38 vdd 2 tie_low vdd hvtpfet l=6e-08 w=3.2e-07 $X=1025 $Y=32908 $D=636
M39 vdd vdd vdd vdd hvtpfet l=6e-08 w=3e-07 $X=1070 $Y=1094 $D=636
M40 vdd vdd vdd vdd hvtpfet l=6e-08 w=3e-07 $X=1070 $Y=1354 $D=636
M41 vdd vdd vdd vdd hvtpfet l=6e-08 w=3e-07 $X=1070 $Y=1864 $D=636
M42 vdd vdd vdd vdd hvtpfet l=6e-08 w=3e-07 $X=1070 $Y=2124 $D=636
M43 vdd vdd vdd vdd hvtpfet l=6e-08 w=3e-07 $X=1070 $Y=48949 $D=636
M44 vdd vdd vdd vdd hvtpfet l=6e-08 w=3e-07 $X=1070 $Y=49209 $D=636
M45 vdd vdd vdd vdd hvtpfet l=6e-08 w=3e-07 $X=1070 $Y=49719 $D=636
M46 vdd vdd vdd vdd hvtpfet l=6e-08 w=3e-07 $X=1070 $Y=49979 $D=636
M47 vdd vdd vdd vdd hvtpfet l=6e-08 w=8e-07 $X=1073 $Y=-170 $D=636
M48 vdd vdd vdd vdd hvtpfet l=6e-08 w=8e-07 $X=1073 $Y=50503 $D=636
M49 vdd tie_low 10 vdd hvtpfet l=6e-08 w=8e-07 $X=1130 $Y=5556 $D=636
M50 vdd tie_low 11 vdd hvtpfet l=6e-08 w=4e-07 $X=1130 $Y=10611 $D=636
M51 vdd tie_low 12 vdd hvtpfet l=6e-08 w=4e-07 $X=1130 $Y=12911 $D=636
M52 vdd tie_low 13 vdd hvtpfet l=6e-08 w=4e-07 $X=1130 $Y=37822 $D=636
M53 vdd tie_low 14 vdd hvtpfet l=6e-08 w=4e-07 $X=1130 $Y=40122 $D=636
M54 vdd tie_low 15 vdd hvtpfet l=6e-08 w=8e-07 $X=1130 $Y=44777 $D=636
M55 vdd 5 21 vdd hvtpfet l=6e-08 w=4.8e-07 $X=1285 $Y=27313 $D=636
M56 vdd 5 22 vdd hvtpfet l=6e-08 w=4.8e-07 $X=1285 $Y=29008 $D=636
M57 vdd vdd vdd vdd hvtpfet l=6e-08 w=8e-07 $X=1333 $Y=-170 $D=636
M58 vdd vdd vdd vdd hvtpfet l=6e-08 w=8e-07 $X=1333 $Y=50503 $D=636
.ends

************************************************************************
* Library Name: XMC55_DPS
* Cell Name:    xmc55_dps_collar_dq_8_bw
************************************************************************
.SUBCKT xmc55_dps_collar_dq_8_bw bwena bwena_int bwenb bwenb_int da da_int db 
+ db_int qa qa_int qb qb_int vdd vss
** N=649 EP=14 IP=0 FDC=76
D0 vss bwena diodenx AREA=7.04e-14 $X=4187 $Y=130 $D=2
D1 vss da diodenx AREA=7.04e-14 $X=6092 $Y=130 $D=2
D2 vss db diodenx AREA=7.04e-14 $X=8010 $Y=130 $D=2
D3 vss bwenb diodenx AREA=7.04e-14 $X=9915 $Y=130 $D=2
M4 12 vdd vss vss hvtnfet l=6e-08 w=6e-07 $X=580 $Y=1420 $D=616
M5 13 vdd vss vss hvtnfet l=6e-08 w=9e-07 $X=1090 $Y=1120 $D=616
M6 vss vdd 13 vss hvtnfet l=6e-08 w=9e-07 $X=1350 $Y=1120 $D=616
M7 14 vdd vss vss hvtnfet l=6e-08 w=9e-07 $X=1610 $Y=1120 $D=616
M8 vss vdd 14 vss hvtnfet l=6e-08 w=9e-07 $X=1870 $Y=1120 $D=616
M9 vss vdd 15 vss hvtnfet l=6e-08 w=6e-07 $X=2380 $Y=1420 $D=616
M10 16 vdd vss vss hvtnfet l=6e-08 w=6e-07 $X=2890 $Y=1420 $D=616
M11 17 vdd vss vss hvtnfet l=6e-08 w=9e-07 $X=3400 $Y=1120 $D=616
M12 vss vdd 17 vss hvtnfet l=6e-08 w=9e-07 $X=3660 $Y=1120 $D=616
M13 3 bwena vss vss hvtnfet l=6e-08 w=6e-07 $X=4400 $Y=1420 $D=616
M14 bwena_int 3 vss vss hvtnfet l=6e-08 w=9e-07 $X=4910 $Y=1120 $D=616
M15 vss 3 bwena_int vss hvtnfet l=6e-08 w=9e-07 $X=5170 $Y=1120 $D=616
M16 qa qa_int vss vss hvtnfet l=6e-08 w=9e-07 $X=5430 $Y=1120 $D=616
M17 vss qa_int qa vss hvtnfet l=6e-08 w=9e-07 $X=5690 $Y=1120 $D=616
M18 vss vdd 20 vss hvtnfet l=6e-08 w=6e-07 $X=6200 $Y=1420 $D=616
M19 6 da vss vss hvtnfet l=6e-08 w=6e-07 $X=6710 $Y=1420 $D=616
M20 da_int 6 vss vss hvtnfet l=6e-08 w=9e-07 $X=7220 $Y=1120 $D=616
M21 vss 6 da_int vss hvtnfet l=6e-08 w=9e-07 $X=7480 $Y=1120 $D=616
M22 db_int 7 vss vss hvtnfet l=6e-08 w=9e-07 $X=7740 $Y=1120 $D=616
M23 vss 7 db_int vss hvtnfet l=6e-08 w=9e-07 $X=8000 $Y=1120 $D=616
M24 vss db 7 vss hvtnfet l=6e-08 w=6e-07 $X=8510 $Y=1420 $D=616
M25 24 vdd vss vss hvtnfet l=6e-08 w=6e-07 $X=9020 $Y=1420 $D=616
M26 qb qb_int vss vss hvtnfet l=6e-08 w=9e-07 $X=9530 $Y=1120 $D=616
M27 vss qb_int qb vss hvtnfet l=6e-08 w=9e-07 $X=9790 $Y=1120 $D=616
M28 bwenb_int 10 vss vss hvtnfet l=6e-08 w=9e-07 $X=10050 $Y=1120 $D=616
M29 vss 10 bwenb_int vss hvtnfet l=6e-08 w=9e-07 $X=10310 $Y=1120 $D=616
M30 vss bwenb 10 vss hvtnfet l=6e-08 w=6e-07 $X=10820 $Y=1420 $D=616
M31 26 vdd vss vss hvtnfet l=6e-08 w=9e-07 $X=11560 $Y=1120 $D=616
M32 vss vdd 26 vss hvtnfet l=6e-08 w=9e-07 $X=11820 $Y=1120 $D=616
M33 vss vdd 27 vss hvtnfet l=6e-08 w=6e-07 $X=12330 $Y=1420 $D=616
M34 28 vdd vss vss hvtnfet l=6e-08 w=6e-07 $X=12840 $Y=1420 $D=616
M35 29 vdd vss vss hvtnfet l=6e-08 w=9e-07 $X=13350 $Y=1120 $D=616
M36 vss vdd 29 vss hvtnfet l=6e-08 w=9e-07 $X=13610 $Y=1120 $D=616
M37 30 vdd vss vss hvtnfet l=6e-08 w=9e-07 $X=13870 $Y=1120 $D=616
M38 vss vdd 30 vss hvtnfet l=6e-08 w=9e-07 $X=14130 $Y=1120 $D=616
M39 vss vdd 31 vss hvtnfet l=6e-08 w=6e-07 $X=14640 $Y=1420 $D=616
M40 12 vdd vdd vdd hvtpfet l=6e-08 w=1.2e-06 $X=580 $Y=2685 $D=636
M41 13 vdd vdd vdd hvtpfet l=6e-08 w=1.8e-06 $X=1090 $Y=2340 $D=636
M42 vdd vdd 13 vdd hvtpfet l=6e-08 w=1.8e-06 $X=1350 $Y=2340 $D=636
M43 14 vdd vdd vdd hvtpfet l=6e-08 w=1.8e-06 $X=1610 $Y=2340 $D=636
M44 vdd vdd 14 vdd hvtpfet l=6e-08 w=1.8e-06 $X=1870 $Y=2340 $D=636
M45 vdd vdd 15 vdd hvtpfet l=6e-08 w=1.2e-06 $X=2380 $Y=2685 $D=636
M46 16 vdd vdd vdd hvtpfet l=6e-08 w=1.2e-06 $X=2890 $Y=2685 $D=636
M47 17 vdd vdd vdd hvtpfet l=6e-08 w=1.8e-06 $X=3400 $Y=2340 $D=636
M48 vdd vdd 17 vdd hvtpfet l=6e-08 w=1.8e-06 $X=3660 $Y=2340 $D=636
M49 3 bwena vdd vdd hvtpfet l=6e-08 w=1.2e-06 $X=4400 $Y=2685 $D=636
M50 bwena_int 3 vdd vdd hvtpfet l=6e-08 w=1.8e-06 $X=4910 $Y=2340 $D=636
M51 vdd 3 bwena_int vdd hvtpfet l=6e-08 w=1.8e-06 $X=5170 $Y=2340 $D=636
M52 qa qa_int vdd vdd hvtpfet l=6e-08 w=1.8e-06 $X=5430 $Y=2340 $D=636
M53 vdd qa_int qa vdd hvtpfet l=6e-08 w=1.8e-06 $X=5690 $Y=2340 $D=636
M54 vdd vdd 20 vdd hvtpfet l=6e-08 w=1.2e-06 $X=6200 $Y=2685 $D=636
M55 6 da vdd vdd hvtpfet l=6e-08 w=1.2e-06 $X=6710 $Y=2685 $D=636
M56 da_int 6 vdd vdd hvtpfet l=6e-08 w=1.8e-06 $X=7220 $Y=2340 $D=636
M57 vdd 6 da_int vdd hvtpfet l=6e-08 w=1.8e-06 $X=7480 $Y=2340 $D=636
M58 db_int 7 vdd vdd hvtpfet l=6e-08 w=1.8e-06 $X=7740 $Y=2340 $D=636
M59 vdd 7 db_int vdd hvtpfet l=6e-08 w=1.8e-06 $X=8000 $Y=2340 $D=636
M60 vdd db 7 vdd hvtpfet l=6e-08 w=1.2e-06 $X=8510 $Y=2685 $D=636
M61 24 vdd vdd vdd hvtpfet l=6e-08 w=1.2e-06 $X=9020 $Y=2685 $D=636
M62 qb qb_int vdd vdd hvtpfet l=6e-08 w=1.8e-06 $X=9530 $Y=2340 $D=636
M63 vdd qb_int qb vdd hvtpfet l=6e-08 w=1.8e-06 $X=9790 $Y=2340 $D=636
M64 bwenb_int 10 vdd vdd hvtpfet l=6e-08 w=1.8e-06 $X=10050 $Y=2340 $D=636
M65 vdd 10 bwenb_int vdd hvtpfet l=6e-08 w=1.8e-06 $X=10310 $Y=2340 $D=636
M66 vdd bwenb 10 vdd hvtpfet l=6e-08 w=1.2e-06 $X=10820 $Y=2685 $D=636
M67 26 vdd vdd vdd hvtpfet l=6e-08 w=1.8e-06 $X=11560 $Y=2340 $D=636
M68 vdd vdd 26 vdd hvtpfet l=6e-08 w=1.8e-06 $X=11820 $Y=2340 $D=636
M69 vdd vdd 27 vdd hvtpfet l=6e-08 w=1.2e-06 $X=12330 $Y=2685 $D=636
M70 28 vdd vdd vdd hvtpfet l=6e-08 w=1.2e-06 $X=12840 $Y=2685 $D=636
M71 29 vdd vdd vdd hvtpfet l=6e-08 w=1.8e-06 $X=13350 $Y=2340 $D=636
M72 vdd vdd 29 vdd hvtpfet l=6e-08 w=1.8e-06 $X=13610 $Y=2340 $D=636
M73 30 vdd vdd vdd hvtpfet l=6e-08 w=1.8e-06 $X=13870 $Y=2340 $D=636
M74 vdd vdd 30 vdd hvtpfet l=6e-08 w=1.8e-06 $X=14130 $Y=2340 $D=636
M75 vdd vdd 31 vdd hvtpfet l=6e-08 w=1.2e-06 $X=14640 $Y=2685 $D=636
.ends

************************************************************************
* Library Name: XMC55_DPS
* Cell Name:    xmc55_dps_local_ctrl4
************************************************************************
.SUBCKT xmc55_dps_local_ctrl4 aa<12> aa<11> aa<10> aa<9> aa<8> aa<7> aa<6> 
+ aa<5> aa<4> aa<3> aa<2> aa<1> aa<0> ab<12> ab<11> ab<10> ab<9> ab<8> ab<7> 
+ ab<6> ab<5> ab<4> ab<3> ab<2> ab<1> ab<0> b_pxaa<3> b_pxaa<2> b_pxaa<1> 
+ b_pxaa<0> b_pxab<3> b_pxab<2> b_pxab<1> b_pxab<0> b_pxba_n<7> b_pxba_n<6> 
+ b_pxba_n<5> b_pxba_n<4> b_pxba_n<3> b_pxba_n<2> b_pxba_n<1> b_pxba_n<0> 
+ b_pxbb_n<7> b_pxbb_n<6> b_pxbb_n<5> b_pxbb_n<4> b_pxbb_n<3> b_pxbb_n<2> 
+ b_pxbb_n<1> b_pxbb_n<0> b_pxca_n<7> b_pxca_n<6> b_pxca_n<5> b_pxca_n<4> 
+ b_pxca_n<3> b_pxca_n<2> b_pxca_n<1> b_pxca_n<0> b_pxcb_n<7> b_pxcb_n<6> 
+ b_pxcb_n<5> b_pxcb_n<4> b_pxcb_n<3> b_pxcb_n<2> b_pxcb_n<1> b_pxcb_n<0> cena 
+ cenb clka clkb dbl_pd_n<3> dbl_pd_n<2> dbl_pd_n<1> dbl_pd_n<0> ddqa ddqa_n 
+ ddqb ddqb_n dwla<1> dwla<0> dwlb<1> dwlb<0> l_clk_dqa l_clk_dqa_n l_clk_dqb 
+ l_clk_dqb_n l_lwea l_lweb l_sa_prea_n l_sa_preb_n l_saea_n l_saeb_n lb_ca<3> 
+ lb_ca<2> lb_ca<1> lb_ca<0> lb_cb<3> lb_cb<2> lb_cb<1> lb_cb<0> lb_ma<3> 
+ lb_ma<2> lb_ma<1> lb_ma<0> lb_mb<3> lb_mb<2> lb_mb<1> lb_mb<0> lb_tm_prea_n 
+ lb_tm_preb_n lt_ca<3> lt_ca<2> lt_ca<1> lt_ca<0> lt_cb<3> lt_cb<2> lt_cb<1> 
+ lt_cb<0> lt_ma<3> lt_ma<2> lt_ma<1> lt_ma<0> lt_mb<3> lt_mb<2> lt_mb<1> 
+ lt_mb<0> lt_tm_prea_n lt_tm_preb_n r_clk_dqa r_clk_dqa_n r_clk_dqb 
+ r_clk_dqb_n r_lwea r_lweb r_sa_prea_n r_sa_preb_n r_saea_n r_saeb_n rb_ca<3> 
+ rb_ca<2> rb_ca<1> rb_ca<0> rb_cb<3> rb_cb<2> rb_cb<1> rb_cb<0> rb_ma<3> 
+ rb_ma<2> rb_ma<1> rb_ma<0> rb_mb<3> rb_mb<2> rb_mb<1> rb_mb<0> rb_tm_prea_n 
+ rb_tm_preb_n rt_ca<3> rt_ca<2> rt_ca<1> rt_ca<0> rt_cb<3> rt_cb<2> rt_cb<1> 
+ rt_cb<0> rt_ma<3> rt_ma<2> rt_ma<1> rt_ma<0> rt_mb<3> rt_mb<2> rt_mb<1> 
+ rt_mb<0> rt_tm_prea_n rt_tm_preb_n stclka stclkb t_pxaa<3> t_pxaa<2> 
+ t_pxaa<1> t_pxaa<0> t_pxab<3> t_pxab<2> t_pxab<1> t_pxab<0> t_pxba_n<7> 
+ t_pxba_n<6> t_pxba_n<5> t_pxba_n<4> t_pxba_n<3> t_pxba_n<2> t_pxba_n<1> 
+ t_pxba_n<0> t_pxbb_n<7> t_pxbb_n<6> t_pxbb_n<5> t_pxbb_n<4> t_pxbb_n<3> 
+ t_pxbb_n<2> t_pxbb_n<1> t_pxbb_n<0> t_pxca_n<7> t_pxca_n<6> t_pxca_n<5> 
+ t_pxca_n<4> t_pxca_n<3> t_pxca_n<2> t_pxca_n<1> t_pxca_n<0> t_pxcb_n<7> 
+ t_pxcb_n<6> t_pxcb_n<5> t_pxcb_n<4> t_pxcb_n<3> t_pxcb_n<2> t_pxcb_n<1> 
+ t_pxcb_n<0> tm<9> tm<8> tm<7> tm<6> tm<5> tm<4> tm<3> tm<2> tm<1> tm<0> vdd 
+ vss wena wenb
** N=19591 EP=230 IP=0 FDC=3266
M0 vss 5 15 vss hvtnfet l=6e-08 w=6e-07 $X=965 $Y=37277 $D=616
M1 11 1 vss vss hvtnfet l=6e-08 w=6e-07 $X=1225 $Y=336 $D=616
M2 12 2 vss vss hvtnfet l=6e-08 w=6e-07 $X=1225 $Y=5566 $D=616
M3 13 3 vss vss hvtnfet l=6e-08 w=6e-07 $X=1225 $Y=6796 $D=616
M4 14 4 vss vss hvtnfet l=6e-08 w=6e-07 $X=1225 $Y=12026 $D=616
M5 lb_tm_preb_n 20 vss vss hvtnfet l=6e-08 w=1.287e-06 $X=1225 $Y=13280 $D=616
M6 lt_tm_preb_n 21 vss vss hvtnfet l=6e-08 w=1.287e-06 $X=1225 $Y=20124 $D=616
M7 vss 8 l_clk_dqb vss hvtnfet l=6e-08 w=1.26e-06 $X=1225 $Y=22041 $D=616
M8 vss 9 l_clk_dqb_n vss hvtnfet l=6e-08 w=1.26e-06 $X=1225 $Y=29007 $D=616
M9 l_lweb 10 vss vss hvtnfet l=6e-08 w=1.287e-06 $X=1225 $Y=30897 $D=616
M10 15 5 vss vss hvtnfet l=6e-08 w=6e-07 $X=1225 $Y=37277 $D=616
M11 16 4 vss vss hvtnfet l=6e-08 w=6e-07 $X=1225 $Y=38507 $D=616
M12 17 3 vss vss hvtnfet l=6e-08 w=6e-07 $X=1225 $Y=43737 $D=616
M13 18 6 vss vss hvtnfet l=6e-08 w=6e-07 $X=1225 $Y=44967 $D=616
M14 19 7 vss vss hvtnfet l=6e-08 w=6e-07 $X=1225 $Y=50197 $D=616
M15 vss 20 lb_tm_preb_n vss hvtnfet l=6e-08 w=1.287e-06 $X=1485 $Y=13280 $D=616
M16 vss 21 lt_tm_preb_n vss hvtnfet l=6e-08 w=1.287e-06 $X=1485 $Y=20124 $D=616
M17 l_clk_dqb 8 vss vss hvtnfet l=6e-08 w=1.26e-06 $X=1485 $Y=22041 $D=616
M18 l_clk_dqb_n 9 vss vss hvtnfet l=6e-08 w=1.26e-06 $X=1485 $Y=29007 $D=616
M19 vss 10 l_lweb vss hvtnfet l=6e-08 w=1.287e-06 $X=1485 $Y=30897 $D=616
M20 lb_cb<0> 11 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=1735 $Y=328 $D=616
M21 lb_cb<2> 12 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=1735 $Y=5316 $D=616
M22 lb_mb<0> 13 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=1735 $Y=6788 $D=616
M23 lb_mb<2> 14 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=1735 $Y=11776 $D=616
M24 l_saeb_n 15 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=1735 $Y=37027 $D=616
M25 lt_mb<2> 16 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=1735 $Y=38499 $D=616
M26 lt_mb<0> 17 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=1735 $Y=43487 $D=616
M27 lt_cb<2> 18 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=1735 $Y=44959 $D=616
M28 lt_cb<0> 19 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=1735 $Y=49947 $D=616
M29 vss 8 l_clk_dqb vss hvtnfet l=6e-08 w=1.26e-06 $X=1745 $Y=22041 $D=616
M30 vss 9 l_clk_dqb_n vss hvtnfet l=6e-08 w=1.26e-06 $X=1745 $Y=29007 $D=616
M31 vss 11 lb_cb<0> vss hvtnfet l=6e-08 w=8.58e-07 $X=1995 $Y=328 $D=616
M32 vss 12 lb_cb<2> vss hvtnfet l=6e-08 w=8.58e-07 $X=1995 $Y=5316 $D=616
M33 vss 13 lb_mb<0> vss hvtnfet l=6e-08 w=8.58e-07 $X=1995 $Y=6788 $D=616
M34 vss 14 lb_mb<2> vss hvtnfet l=6e-08 w=8.58e-07 $X=1995 $Y=11776 $D=616
M35 vss 24 20 vss hvtnfet l=6e-08 w=6e-07 $X=1995 $Y=13282 $D=616
M36 vss 25 21 vss hvtnfet l=6e-08 w=6e-07 $X=1995 $Y=20809 $D=616
M37 vss 15 l_saeb_n vss hvtnfet l=6e-08 w=8.58e-07 $X=1995 $Y=37027 $D=616
M38 vss 16 lt_mb<2> vss hvtnfet l=6e-08 w=8.58e-07 $X=1995 $Y=38499 $D=616
M39 vss 17 lt_mb<0> vss hvtnfet l=6e-08 w=8.58e-07 $X=1995 $Y=43487 $D=616
M40 vss 18 lt_cb<2> vss hvtnfet l=6e-08 w=8.58e-07 $X=1995 $Y=44959 $D=616
M41 vss 19 lt_cb<0> vss hvtnfet l=6e-08 w=8.58e-07 $X=1995 $Y=49947 $D=616
M42 8 clkb vss vss hvtnfet l=6e-08 w=1.05e-06 $X=2005 $Y=22251 $D=616
M43 9 23 vss vss hvtnfet l=6e-08 w=1.05e-06 $X=2005 $Y=29007 $D=616
M44 lb_cb<0> 11 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=2255 $Y=328 $D=616
M45 lb_cb<2> 12 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=2255 $Y=5316 $D=616
M46 lb_mb<0> 13 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=2255 $Y=6788 $D=616
M47 lb_mb<2> 14 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=2255 $Y=11776 $D=616
M48 l_saeb_n 15 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=2255 $Y=37027 $D=616
M49 lt_mb<2> 16 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=2255 $Y=38499 $D=616
M50 lt_mb<0> 17 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=2255 $Y=43487 $D=616
M51 lt_cb<2> 18 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=2255 $Y=44959 $D=616
M52 lt_cb<0> 19 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=2255 $Y=49947 $D=616
M53 vss 15 l_saeb_n vss hvtnfet l=6e-08 w=8.58e-07 $X=2515 $Y=37027 $D=616
M54 vss 34 lb_cb<1> vss hvtnfet l=6e-08 w=8.58e-07 $X=2765 $Y=328 $D=616
M55 vss 35 lb_cb<3> vss hvtnfet l=6e-08 w=8.58e-07 $X=2765 $Y=5316 $D=616
M56 vss 36 lb_mb<1> vss hvtnfet l=6e-08 w=8.58e-07 $X=2765 $Y=6788 $D=616
M57 vss 37 lb_mb<3> vss hvtnfet l=6e-08 w=8.58e-07 $X=2765 $Y=11776 $D=616
M58 vss 39 lt_mb<3> vss hvtnfet l=6e-08 w=8.58e-07 $X=2765 $Y=38499 $D=616
M59 vss 40 lt_mb<1> vss hvtnfet l=6e-08 w=8.58e-07 $X=2765 $Y=43487 $D=616
M60 vss 41 lt_cb<3> vss hvtnfet l=6e-08 w=8.58e-07 $X=2765 $Y=44959 $D=616
M61 vss 42 lt_cb<1> vss hvtnfet l=6e-08 w=8.58e-07 $X=2765 $Y=49947 $D=616
M62 l_saeb_n 15 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=2775 $Y=37027 $D=616
M63 909 26 vss vss hvtnfet l=6e-08 w=1.8e-07 $X=2821 $Y=17143 $D=616
M64 26 28 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=2821 $Y=17812 $D=616
M65 4 29 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=2821 $Y=18983 $D=616
M66 910 4 vss vss hvtnfet l=6e-08 w=1.8e-07 $X=2821 $Y=19609 $D=616
M67 911 27 vss vss hvtnfet l=6e-08 w=1.8e-07 $X=2821 $Y=24063 $D=616
M68 27 30 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=2821 $Y=24732 $D=616
M69 3 31 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=2821 $Y=25903 $D=616
M70 912 3 vss vss hvtnfet l=6e-08 w=1.8e-07 $X=2821 $Y=26529 $D=616
M71 lb_cb<1> 34 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=3025 $Y=328 $D=616
M72 lb_cb<3> 35 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=3025 $Y=5316 $D=616
M73 lb_mb<1> 36 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=3025 $Y=6788 $D=616
M74 lb_mb<3> 37 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=3025 $Y=11776 $D=616
M75 lt_mb<3> 39 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=3025 $Y=38499 $D=616
M76 lt_mb<1> 40 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=3025 $Y=43487 $D=616
M77 lt_cb<3> 41 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=3025 $Y=44959 $D=616
M78 lt_cb<1> 42 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=3025 $Y=49947 $D=616
M79 28 33 909 vss hvtnfet l=6e-08 w=1.8e-07 $X=3081 $Y=17143 $D=616
M80 vss 28 26 vss hvtnfet l=6e-08 w=1.37e-07 $X=3081 $Y=17812 $D=616
M81 vss 29 4 vss hvtnfet l=6e-08 w=1.37e-07 $X=3081 $Y=18983 $D=616
M82 29 33 910 vss hvtnfet l=6e-08 w=1.8e-07 $X=3081 $Y=19609 $D=616
M83 30 33 911 vss hvtnfet l=6e-08 w=1.8e-07 $X=3081 $Y=24063 $D=616
M84 vss 30 27 vss hvtnfet l=6e-08 w=1.37e-07 $X=3081 $Y=24732 $D=616
M85 vss 31 3 vss hvtnfet l=6e-08 w=1.37e-07 $X=3081 $Y=25903 $D=616
M86 31 33 912 vss hvtnfet l=6e-08 w=1.8e-07 $X=3081 $Y=26529 $D=616
M87 vss 34 lb_cb<1> vss hvtnfet l=6e-08 w=8.58e-07 $X=3285 $Y=328 $D=616
M88 vss 35 lb_cb<3> vss hvtnfet l=6e-08 w=8.58e-07 $X=3285 $Y=5316 $D=616
M89 vss 36 lb_mb<1> vss hvtnfet l=6e-08 w=8.58e-07 $X=3285 $Y=6788 $D=616
M90 vss 37 lb_mb<3> vss hvtnfet l=6e-08 w=8.58e-07 $X=3285 $Y=11776 $D=616
M91 vss 51 l_sa_preb_n vss hvtnfet l=6e-08 w=8.58e-07 $X=3285 $Y=37027 $D=616
M92 vss 39 lt_mb<3> vss hvtnfet l=6e-08 w=8.58e-07 $X=3285 $Y=38499 $D=616
M93 vss 40 lt_mb<1> vss hvtnfet l=6e-08 w=8.58e-07 $X=3285 $Y=43487 $D=616
M94 vss 41 lt_cb<3> vss hvtnfet l=6e-08 w=8.58e-07 $X=3285 $Y=44959 $D=616
M95 vss 42 lt_cb<1> vss hvtnfet l=6e-08 w=8.58e-07 $X=3285 $Y=49947 $D=616
M96 vss ab<2> 44 vss hvtnfet l=6e-08 w=2.74e-07 $X=3396 $Y=13476 $D=616
M97 l_sa_preb_n 51 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=3545 $Y=37027 $D=616
M98 913 43 vss vss hvtnfet l=6e-08 w=8.23e-07 $X=3591 $Y=17143 $D=616
M99 914 43 vss vss hvtnfet l=6e-08 w=8.23e-07 $X=3591 $Y=18966 $D=616
M100 915 43 vss vss hvtnfet l=6e-08 w=8.23e-07 $X=3591 $Y=24063 $D=616
M101 916 43 vss vss hvtnfet l=6e-08 w=8.23e-07 $X=3591 $Y=25886 $D=616
M102 52 stclkb vss vss hvtnfet l=6e-08 w=2.74e-07 $X=3705 $Y=30668 $D=616
M103 vss 47 34 vss hvtnfet l=6e-08 w=6e-07 $X=3795 $Y=336 $D=616
M104 vss 48 35 vss hvtnfet l=6e-08 w=6e-07 $X=3795 $Y=5566 $D=616
M105 vss 27 36 vss hvtnfet l=6e-08 w=6e-07 $X=3795 $Y=6796 $D=616
M106 vss 26 37 vss hvtnfet l=6e-08 w=6e-07 $X=3795 $Y=12026 $D=616
M107 vss 26 39 vss hvtnfet l=6e-08 w=6e-07 $X=3795 $Y=38507 $D=616
M108 vss 27 40 vss hvtnfet l=6e-08 w=6e-07 $X=3795 $Y=43737 $D=616
M109 vss 49 41 vss hvtnfet l=6e-08 w=6e-07 $X=3795 $Y=44967 $D=616
M110 vss 50 42 vss hvtnfet l=6e-08 w=6e-07 $X=3795 $Y=50197 $D=616
M111 vss 51 l_sa_preb_n vss hvtnfet l=6e-08 w=8.58e-07 $X=3805 $Y=37027 $D=616
M112 917 45 913 vss hvtnfet l=6e-08 w=5.49e-07 $X=3861 $Y=17143 $D=616
M113 918 45 914 vss hvtnfet l=6e-08 w=5.49e-07 $X=3861 $Y=19240 $D=616
M114 919 46 915 vss hvtnfet l=6e-08 w=5.49e-07 $X=3861 $Y=24063 $D=616
M115 920 46 916 vss hvtnfet l=6e-08 w=5.49e-07 $X=3861 $Y=26160 $D=616
M116 53 44 vss vss hvtnfet l=6e-08 w=2.74e-07 $X=3906 $Y=13476 $D=616
M117 vss clkb 43 vss hvtnfet l=6e-08 w=6e-07 $X=4066 $Y=32403 $D=616
M118 28 53 917 vss hvtnfet l=6e-08 w=5.49e-07 $X=4121 $Y=17143 $D=616
M119 29 44 918 vss hvtnfet l=6e-08 w=5.49e-07 $X=4121 $Y=19240 $D=616
M120 30 53 919 vss hvtnfet l=6e-08 w=5.49e-07 $X=4121 $Y=24063 $D=616
M121 31 44 920 vss hvtnfet l=6e-08 w=5.49e-07 $X=4121 $Y=26160 $D=616
M122 vss 52 59 vss hvtnfet l=6e-08 w=5.49e-07 $X=4215 $Y=30668 $D=616
M123 vss 55 51 vss hvtnfet l=6e-08 w=6e-07 $X=4315 $Y=37277 $D=616
M124 43 clkb vss vss hvtnfet l=6e-08 w=6e-07 $X=4326 $Y=32403 $D=616
M125 vss ab<3> 46 vss hvtnfet l=6e-08 w=2.74e-07 $X=4416 $Y=13476 $D=616
M126 59 56 vss vss hvtnfet l=6e-08 w=5.49e-07 $X=4475 $Y=30668 $D=616
M127 b_pxab<0> 60 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=4550 $Y=336 $D=616
M128 60 61 vss vss hvtnfet l=6e-08 w=5e-07 $X=4550 $Y=6701 $D=616
M129 61 62 vss vss hvtnfet l=6e-08 w=3e-07 $X=4550 $Y=7831 $D=616
M130 921 57 vss vss hvtnfet l=6e-08 w=4.11e-07 $X=4550 $Y=11276 $D=616
M131 922 57 vss vss hvtnfet l=6e-08 w=4.11e-07 $X=4550 $Y=39446 $D=616
M132 64 63 vss vss hvtnfet l=6e-08 w=3e-07 $X=4550 $Y=43002 $D=616
M133 65 64 vss vss hvtnfet l=6e-08 w=5e-07 $X=4550 $Y=43932 $D=616
M134 t_pxab<0> 65 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=4550 $Y=49512 $D=616
M135 vss 60 b_pxab<0> vss hvtnfet l=6e-08 w=1.285e-06 $X=4810 $Y=336 $D=616
M136 vss 61 60 vss hvtnfet l=6e-08 w=5e-07 $X=4810 $Y=6701 $D=616
M137 vss 62 61 vss hvtnfet l=6e-08 w=3e-07 $X=4810 $Y=7831 $D=616
M138 62 24 921 vss hvtnfet l=6e-08 w=4.11e-07 $X=4810 $Y=11276 $D=616
M139 63 25 922 vss hvtnfet l=6e-08 w=4.11e-07 $X=4810 $Y=39446 $D=616
M140 vss 63 64 vss hvtnfet l=6e-08 w=3e-07 $X=4810 $Y=43002 $D=616
M141 vss 64 65 vss hvtnfet l=6e-08 w=5e-07 $X=4810 $Y=43932 $D=616
M142 vss 65 t_pxab<0> vss hvtnfet l=6e-08 w=1.285e-06 $X=4810 $Y=49512 $D=616
M143 45 46 vss vss hvtnfet l=6e-08 w=2.74e-07 $X=4926 $Y=13476 $D=616
M144 vss 66 586 vss hvtnfet l=1.4e-07 w=3.2e-07 $X=4939 $Y=37127 $D=616
M145 vss 59 56 vss hvtnfet l=6e-08 w=5.49e-07 $X=4985 $Y=30668 $D=616
M146 vss 58 587 vss hvtnfet l=6e-08 w=3.2e-07 $X=5069 $Y=32828 $D=616
M147 923 67 vss vss hvtnfet l=6e-08 w=1.8e-07 $X=5141 $Y=17143 $D=616
M148 67 73 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=5141 $Y=17812 $D=616
M149 68 74 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=5141 $Y=18983 $D=616
M150 924 68 vss vss hvtnfet l=6e-08 w=1.8e-07 $X=5141 $Y=19609 $D=616
M151 925 69 vss vss hvtnfet l=6e-08 w=1.8e-07 $X=5141 $Y=24063 $D=616
M152 69 75 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=5141 $Y=24732 $D=616
M153 57 76 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=5141 $Y=25903 $D=616
M154 926 57 vss vss hvtnfet l=6e-08 w=1.8e-07 $X=5141 $Y=26529 $D=616
M155 56 70 vss vss hvtnfet l=6e-08 w=5.49e-07 $X=5245 $Y=30668 $D=616
M156 66 71 vss vss hvtnfet l=1.4e-07 w=3.2e-07 $X=5279 $Y=37127 $D=616
M157 b_pxab<1> 78 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=5320 $Y=336 $D=616
M158 78 79 vss vss hvtnfet l=6e-08 w=5e-07 $X=5320 $Y=6701 $D=616
M159 79 80 vss vss hvtnfet l=6e-08 w=3e-07 $X=5320 $Y=7831 $D=616
M160 927 24 80 vss hvtnfet l=6e-08 w=4.11e-07 $X=5320 $Y=11276 $D=616
M161 928 25 81 vss hvtnfet l=6e-08 w=4.11e-07 $X=5320 $Y=39446 $D=616
M162 82 81 vss vss hvtnfet l=6e-08 w=3e-07 $X=5320 $Y=43002 $D=616
M163 83 82 vss vss hvtnfet l=6e-08 w=5e-07 $X=5320 $Y=43932 $D=616
M164 t_pxab<1> 83 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=5320 $Y=49512 $D=616
M165 73 33 923 vss hvtnfet l=6e-08 w=1.8e-07 $X=5401 $Y=17143 $D=616
M166 vss 73 67 vss hvtnfet l=6e-08 w=1.37e-07 $X=5401 $Y=17812 $D=616
M167 vss 74 68 vss hvtnfet l=6e-08 w=1.37e-07 $X=5401 $Y=18983 $D=616
M168 74 33 924 vss hvtnfet l=6e-08 w=1.8e-07 $X=5401 $Y=19609 $D=616
M169 75 33 925 vss hvtnfet l=6e-08 w=1.8e-07 $X=5401 $Y=24063 $D=616
M170 vss 75 69 vss hvtnfet l=6e-08 w=1.37e-07 $X=5401 $Y=24732 $D=616
M171 vss 76 57 vss hvtnfet l=6e-08 w=1.37e-07 $X=5401 $Y=25903 $D=616
M172 76 33 926 vss hvtnfet l=6e-08 w=1.8e-07 $X=5401 $Y=26529 $D=616
M173 929 72 vss vss hvtnfet l=6e-08 w=6.4e-07 $X=5579 $Y=32508 $D=616
M174 vss 78 b_pxab<1> vss hvtnfet l=6e-08 w=1.285e-06 $X=5580 $Y=336 $D=616
M175 vss 79 78 vss hvtnfet l=6e-08 w=5e-07 $X=5580 $Y=6701 $D=616
M176 vss 80 79 vss hvtnfet l=6e-08 w=3e-07 $X=5580 $Y=7831 $D=616
M177 vss 69 927 vss hvtnfet l=6e-08 w=4.11e-07 $X=5580 $Y=11276 $D=616
M178 vss 69 928 vss hvtnfet l=6e-08 w=4.11e-07 $X=5580 $Y=39446 $D=616
M179 vss 81 82 vss hvtnfet l=6e-08 w=3e-07 $X=5580 $Y=43002 $D=616
M180 vss 82 83 vss hvtnfet l=6e-08 w=5e-07 $X=5580 $Y=43932 $D=616
M181 vss 83 t_pxab<1> vss hvtnfet l=6e-08 w=1.285e-06 $X=5580 $Y=49512 $D=616
M182 vss ab<5> 86 vss hvtnfet l=6e-08 w=2.74e-07 $X=5716 $Y=13476 $D=616
M183 5 85 929 vss hvtnfet l=6e-08 w=6.4e-07 $X=5839 $Y=32508 $D=616
M184 930 43 vss vss hvtnfet l=6e-08 w=8.23e-07 $X=5911 $Y=17143 $D=616
M185 931 43 vss vss hvtnfet l=6e-08 w=8.23e-07 $X=5911 $Y=18966 $D=616
M186 932 43 vss vss hvtnfet l=6e-08 w=8.23e-07 $X=5911 $Y=24063 $D=616
M187 933 43 vss vss hvtnfet l=6e-08 w=8.23e-07 $X=5911 $Y=25886 $D=616
M188 70 clkb vss vss hvtnfet l=6e-08 w=6e-07 $X=6015 $Y=30668 $D=616
M189 vss ddqb 71 vss hvtnfet l=6e-08 w=2.4e-07 $X=6079 $Y=37292 $D=616
M190 b_pxab<2> 90 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=6090 $Y=336 $D=616
M191 90 91 vss vss hvtnfet l=6e-08 w=5e-07 $X=6090 $Y=6701 $D=616
M192 91 92 vss vss hvtnfet l=6e-08 w=3e-07 $X=6090 $Y=7831 $D=616
M193 934 68 vss vss hvtnfet l=6e-08 w=4.11e-07 $X=6090 $Y=11276 $D=616
M194 935 68 vss vss hvtnfet l=6e-08 w=4.11e-07 $X=6090 $Y=39446 $D=616
M195 94 93 vss vss hvtnfet l=6e-08 w=3e-07 $X=6090 $Y=43002 $D=616
M196 95 94 vss vss hvtnfet l=6e-08 w=5e-07 $X=6090 $Y=43932 $D=616
M197 t_pxab<2> 95 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=6090 $Y=49512 $D=616
M198 936 87 930 vss hvtnfet l=6e-08 w=5.49e-07 $X=6181 $Y=17143 $D=616
M199 937 87 931 vss hvtnfet l=6e-08 w=5.49e-07 $X=6181 $Y=19240 $D=616
M200 938 88 932 vss hvtnfet l=6e-08 w=5.49e-07 $X=6181 $Y=24063 $D=616
M201 939 88 933 vss hvtnfet l=6e-08 w=5.49e-07 $X=6181 $Y=26160 $D=616
M202 97 86 vss vss hvtnfet l=6e-08 w=2.74e-07 $X=6226 $Y=13476 $D=616
M203 71 ddqb_n vss vss hvtnfet l=6e-08 w=2.4e-07 $X=6339 $Y=37292 $D=616
M204 vss 90 b_pxab<2> vss hvtnfet l=6e-08 w=1.285e-06 $X=6350 $Y=336 $D=616
M205 vss 91 90 vss hvtnfet l=6e-08 w=5e-07 $X=6350 $Y=6701 $D=616
M206 vss 92 91 vss hvtnfet l=6e-08 w=3e-07 $X=6350 $Y=7831 $D=616
M207 92 24 934 vss hvtnfet l=6e-08 w=4.11e-07 $X=6350 $Y=11276 $D=616
M208 93 25 935 vss hvtnfet l=6e-08 w=4.11e-07 $X=6350 $Y=39446 $D=616
M209 vss 93 94 vss hvtnfet l=6e-08 w=3e-07 $X=6350 $Y=43002 $D=616
M210 vss 94 95 vss hvtnfet l=6e-08 w=5e-07 $X=6350 $Y=43932 $D=616
M211 vss 95 t_pxab<2> vss hvtnfet l=6e-08 w=1.285e-06 $X=6350 $Y=49512 $D=616
M212 73 97 936 vss hvtnfet l=6e-08 w=5.49e-07 $X=6441 $Y=17143 $D=616
M213 74 86 937 vss hvtnfet l=6e-08 w=5.49e-07 $X=6441 $Y=19240 $D=616
M214 75 97 938 vss hvtnfet l=6e-08 w=5.49e-07 $X=6441 $Y=24063 $D=616
M215 76 86 939 vss hvtnfet l=6e-08 w=5.49e-07 $X=6441 $Y=26160 $D=616
M216 85 89 vss vss hvtnfet l=6e-08 w=3.2e-07 $X=6524 $Y=32828 $D=616
M217 142 clkb 595 vss hvtnfet l=6e-08 w=8e-07 $X=6525 $Y=30668 $D=616
M218 vss ab<6> 88 vss hvtnfet l=6e-08 w=2.74e-07 $X=6736 $Y=13476 $D=616
M219 595 clkb 142 vss hvtnfet l=6e-08 w=8e-07 $X=6785 $Y=30668 $D=616
M220 b_pxab<3> 99 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=6860 $Y=336 $D=616
M221 99 100 vss vss hvtnfet l=6e-08 w=5e-07 $X=6860 $Y=6701 $D=616
M222 100 101 vss vss hvtnfet l=6e-08 w=3e-07 $X=6860 $Y=7831 $D=616
M223 940 24 101 vss hvtnfet l=6e-08 w=4.11e-07 $X=6860 $Y=11276 $D=616
M224 941 25 102 vss hvtnfet l=6e-08 w=4.11e-07 $X=6860 $Y=39446 $D=616
M225 103 102 vss vss hvtnfet l=6e-08 w=3e-07 $X=6860 $Y=43002 $D=616
M226 104 103 vss vss hvtnfet l=6e-08 w=5e-07 $X=6860 $Y=43932 $D=616
M227 t_pxab<3> 104 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=6860 $Y=49512 $D=616
M228 109 85 vss vss hvtnfet l=6e-08 w=3.2e-07 $X=7034 $Y=32828 $D=616
M229 89 58 vss vss hvtnfet l=6e-08 w=3.2e-07 $X=7069 $Y=37292 $D=616
M230 vss 99 b_pxab<3> vss hvtnfet l=6e-08 w=1.285e-06 $X=7120 $Y=336 $D=616
M231 vss 100 99 vss hvtnfet l=6e-08 w=5e-07 $X=7120 $Y=6701 $D=616
M232 vss 101 100 vss hvtnfet l=6e-08 w=3e-07 $X=7120 $Y=7831 $D=616
M233 vss 67 940 vss hvtnfet l=6e-08 w=4.11e-07 $X=7120 $Y=11276 $D=616
M234 vss 67 941 vss hvtnfet l=6e-08 w=4.11e-07 $X=7120 $Y=39446 $D=616
M235 vss 102 103 vss hvtnfet l=6e-08 w=3e-07 $X=7120 $Y=43002 $D=616
M236 vss 103 104 vss hvtnfet l=6e-08 w=5e-07 $X=7120 $Y=43932 $D=616
M237 vss 104 t_pxab<3> vss hvtnfet l=6e-08 w=1.285e-06 $X=7120 $Y=49512 $D=616
M238 87 88 vss vss hvtnfet l=6e-08 w=2.74e-07 $X=7246 $Y=13476 $D=616
M239 595 59 vss vss hvtnfet l=6e-08 w=8e-07 $X=7295 $Y=30668 $D=616
M240 942 105 vss vss hvtnfet l=6e-08 w=1.8e-07 $X=7461 $Y=17143 $D=616
M241 943 106 vss vss hvtnfet l=6e-08 w=1.8e-07 $X=7461 $Y=19609 $D=616
M242 944 107 vss vss hvtnfet l=6e-08 w=1.8e-07 $X=7461 $Y=24063 $D=616
M243 945 108 vss vss hvtnfet l=6e-08 w=1.8e-07 $X=7461 $Y=26529 $D=616
M244 105 111 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=7476 $Y=17812 $D=616
M245 106 112 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=7476 $Y=18983 $D=616
M246 107 113 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=7476 $Y=24732 $D=616
M247 108 114 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=7476 $Y=25903 $D=616
M248 vss 59 595 vss hvtnfet l=6e-08 w=8e-07 $X=7555 $Y=30668 $D=616
M249 vss 110 89 vss hvtnfet l=1.2e-07 w=1.5e-07 $X=7579 $Y=37297 $D=616
M250 vss 109 119 vss hvtnfet l=2.5e-07 w=3.5e-07 $X=7604 $Y=32613 $D=616
M251 b_pxbb_n<0> 115 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=7630 $Y=336 $D=616
M252 115 116 vss vss hvtnfet l=6e-08 w=5e-07 $X=7630 $Y=6701 $D=616
M253 116 107 vss vss hvtnfet l=6e-08 w=3e-07 $X=7630 $Y=7831 $D=616
M254 117 107 vss vss hvtnfet l=6e-08 w=3e-07 $X=7630 $Y=43002 $D=616
M255 118 117 vss vss hvtnfet l=6e-08 w=5e-07 $X=7630 $Y=43932 $D=616
M256 t_pxbb_n<0> 118 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=7630 $Y=49512 $D=616
M257 111 33 942 vss hvtnfet l=6e-08 w=1.8e-07 $X=7721 $Y=17143 $D=616
M258 112 33 943 vss hvtnfet l=6e-08 w=1.8e-07 $X=7721 $Y=19609 $D=616
M259 113 33 944 vss hvtnfet l=6e-08 w=1.8e-07 $X=7721 $Y=24063 $D=616
M260 114 33 945 vss hvtnfet l=6e-08 w=1.8e-07 $X=7721 $Y=26529 $D=616
M261 vss 111 105 vss hvtnfet l=6e-08 w=1.37e-07 $X=7736 $Y=17812 $D=616
M262 vss 112 106 vss hvtnfet l=6e-08 w=1.37e-07 $X=7736 $Y=18983 $D=616
M263 vss 113 107 vss hvtnfet l=6e-08 w=1.37e-07 $X=7736 $Y=24732 $D=616
M264 vss 114 108 vss hvtnfet l=6e-08 w=1.37e-07 $X=7736 $Y=25903 $D=616
M265 vss 115 b_pxbb_n<0> vss hvtnfet l=6e-08 w=1.285e-06 $X=7890 $Y=336 $D=616
M266 vss 116 115 vss hvtnfet l=6e-08 w=5e-07 $X=7890 $Y=6701 $D=616
M267 vss 107 116 vss hvtnfet l=6e-08 w=3e-07 $X=7890 $Y=7831 $D=616
M268 vss 107 117 vss hvtnfet l=6e-08 w=3e-07 $X=7890 $Y=43002 $D=616
M269 vss 117 118 vss hvtnfet l=6e-08 w=5e-07 $X=7890 $Y=43932 $D=616
M270 vss 118 t_pxbb_n<0> vss hvtnfet l=6e-08 w=1.285e-06 $X=7890 $Y=49512 $D=616
M271 120 119 vss vss hvtnfet l=6e-08 w=3.5e-07 $X=8054 $Y=32613 $D=616
M272 110 89 vss vss hvtnfet l=6e-08 w=3e-07 $X=8149 $Y=37257 $D=616
M273 946 43 vss vss hvtnfet l=6e-08 w=8.23e-07 $X=8231 $Y=17143 $D=616
M274 947 43 vss vss hvtnfet l=6e-08 w=8.23e-07 $X=8231 $Y=18966 $D=616
M275 948 43 vss vss hvtnfet l=6e-08 w=8.23e-07 $X=8231 $Y=24063 $D=616
M276 949 43 vss vss hvtnfet l=6e-08 w=8.23e-07 $X=8231 $Y=25886 $D=616
M277 b_pxbb_n<1> 125 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=8400 $Y=336 $D=616
M278 125 126 vss vss hvtnfet l=6e-08 w=5e-07 $X=8400 $Y=6701 $D=616
M279 126 108 vss vss hvtnfet l=6e-08 w=3e-07 $X=8400 $Y=7831 $D=616
M280 127 108 vss vss hvtnfet l=6e-08 w=3e-07 $X=8400 $Y=43002 $D=616
M281 128 127 vss vss hvtnfet l=6e-08 w=5e-07 $X=8400 $Y=43932 $D=616
M282 t_pxbb_n<1> 128 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=8400 $Y=49512 $D=616
M283 vss 122 121 vss hvtnfet l=6e-08 w=2.74e-07 $X=8466 $Y=13476 $D=616
M284 950 121 946 vss hvtnfet l=6e-08 w=5.49e-07 $X=8501 $Y=17417 $D=616
M285 951 121 947 vss hvtnfet l=6e-08 w=5.49e-07 $X=8501 $Y=18966 $D=616
M286 952 122 948 vss hvtnfet l=6e-08 w=5.49e-07 $X=8501 $Y=24337 $D=616
M287 953 122 949 vss hvtnfet l=6e-08 w=5.49e-07 $X=8501 $Y=25886 $D=616
M288 123 123 vss vss hvtnfet l=6e-08 w=2e-07 $X=8594 $Y=11546 $D=616
M289 954 120 55 vss hvtnfet l=6e-08 w=6.4e-07 $X=8619 $Y=32508 $D=616
M290 dwlb<0> 124 vss vss hvtnfet l=6e-08 w=3e-07 $X=8659 $Y=31098 $D=616
M291 25 124 vss vss hvtnfet l=6e-08 w=3e-07 $X=8659 $Y=37457 $D=616
M292 vss 125 b_pxbb_n<1> vss hvtnfet l=6e-08 w=1.285e-06 $X=8660 $Y=336 $D=616
M293 vss 126 125 vss hvtnfet l=6e-08 w=5e-07 $X=8660 $Y=6701 $D=616
M294 vss 108 126 vss hvtnfet l=6e-08 w=3e-07 $X=8660 $Y=7831 $D=616
M295 vss 108 127 vss hvtnfet l=6e-08 w=3e-07 $X=8660 $Y=43002 $D=616
M296 vss 127 128 vss hvtnfet l=6e-08 w=5e-07 $X=8660 $Y=43932 $D=616
M297 vss 128 t_pxbb_n<1> vss hvtnfet l=6e-08 w=1.285e-06 $X=8660 $Y=49512 $D=616
M298 955 129 950 vss hvtnfet l=6e-08 w=5.49e-07 $X=8761 $Y=17417 $D=616
M299 956 129 951 vss hvtnfet l=6e-08 w=5.49e-07 $X=8761 $Y=18966 $D=616
M300 957 129 952 vss hvtnfet l=6e-08 w=5.49e-07 $X=8761 $Y=24337 $D=616
M301 958 129 953 vss hvtnfet l=6e-08 w=5.49e-07 $X=8761 $Y=25886 $D=616
M302 vss 131 123 vss hvtnfet l=6e-08 w=2e-07 $X=8854 $Y=11546 $D=616
M303 vss vdd 954 vss hvtnfet l=6e-08 w=6.4e-07 $X=8879 $Y=32508 $D=616
M304 vss 124 dwlb<0> vss hvtnfet l=6e-08 w=3e-07 $X=8919 $Y=31098 $D=616
M305 vss 124 25 vss hvtnfet l=6e-08 w=3e-07 $X=8919 $Y=37457 $D=616
M306 122 ab<9> vss vss hvtnfet l=6e-08 w=2.74e-07 $X=8976 $Y=13476 $D=616
M307 111 132 955 vss hvtnfet l=6e-08 w=5.49e-07 $X=9021 $Y=17417 $D=616
M308 112 133 956 vss hvtnfet l=6e-08 w=5.49e-07 $X=9021 $Y=18966 $D=616
M309 113 132 957 vss hvtnfet l=6e-08 w=5.49e-07 $X=9021 $Y=24337 $D=616
M310 114 133 958 vss hvtnfet l=6e-08 w=5.49e-07 $X=9021 $Y=25886 $D=616
M311 b_pxbb_n<2> 135 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=9170 $Y=336 $D=616
M312 135 136 vss vss hvtnfet l=6e-08 w=5e-07 $X=9170 $Y=6701 $D=616
M313 136 137 vss vss hvtnfet l=6e-08 w=3e-07 $X=9170 $Y=7831 $D=616
M314 138 137 vss vss hvtnfet l=6e-08 w=3e-07 $X=9170 $Y=43002 $D=616
M315 139 138 vss vss hvtnfet l=6e-08 w=5e-07 $X=9170 $Y=43932 $D=616
M316 t_pxbb_n<2> 139 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=9170 $Y=49512 $D=616
M317 dwlb<0> 142 vss vss hvtnfet l=6e-08 w=3e-07 $X=9429 $Y=31098 $D=616
M318 25 143 vss vss hvtnfet l=6e-08 w=3e-07 $X=9429 $Y=37457 $D=616
M319 vss 135 b_pxbb_n<2> vss hvtnfet l=6e-08 w=1.285e-06 $X=9430 $Y=336 $D=616
M320 vss 136 135 vss hvtnfet l=6e-08 w=5e-07 $X=9430 $Y=6701 $D=616
M321 vss 137 136 vss hvtnfet l=6e-08 w=3e-07 $X=9430 $Y=7831 $D=616
M322 vss 137 138 vss hvtnfet l=6e-08 w=3e-07 $X=9430 $Y=43002 $D=616
M323 vss 138 139 vss hvtnfet l=6e-08 w=5e-07 $X=9430 $Y=43932 $D=616
M324 vss 139 t_pxbb_n<2> vss hvtnfet l=6e-08 w=1.285e-06 $X=9430 $Y=49512 $D=616
M325 vss 140 1 vss hvtnfet l=6e-08 w=2e-07 $X=9586 $Y=11276 $D=616
M326 vss 141 7 vss hvtnfet l=6e-08 w=2e-07 $X=9586 $Y=39657 $D=616
M327 vss 142 dwlb<0> vss hvtnfet l=6e-08 w=3e-07 $X=9689 $Y=31098 $D=616
M328 vss 143 25 vss hvtnfet l=6e-08 w=3e-07 $X=9689 $Y=37457 $D=616
M329 b_pxbb_n<3> 146 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=9940 $Y=336 $D=616
M330 146 147 vss vss hvtnfet l=6e-08 w=5e-07 $X=9940 $Y=6701 $D=616
M331 147 148 vss vss hvtnfet l=6e-08 w=3e-07 $X=9940 $Y=7831 $D=616
M332 149 148 vss vss hvtnfet l=6e-08 w=3e-07 $X=9940 $Y=43002 $D=616
M333 150 149 vss vss hvtnfet l=6e-08 w=5e-07 $X=9940 $Y=43932 $D=616
M334 t_pxbb_n<3> 150 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=9940 $Y=49512 $D=616
M335 vss ab<8> 129 vss hvtnfet l=6e-08 w=2.74e-07 $X=9986 $Y=13476 $D=616
M336 959 145 vss vss hvtnfet l=6e-08 w=4.11e-07 $X=10096 $Y=11276 $D=616
M337 960 145 vss vss hvtnfet l=6e-08 w=4.11e-07 $X=10096 $Y=39446 $D=616
M338 dwlb<1> 142 vss vss hvtnfet l=6e-08 w=3e-07 $X=10199 $Y=31098 $D=616
M339 24 143 vss vss hvtnfet l=6e-08 w=3e-07 $X=10199 $Y=37457 $D=616
M340 vss 146 b_pxbb_n<3> vss hvtnfet l=6e-08 w=1.285e-06 $X=10200 $Y=336 $D=616
M341 vss 147 146 vss hvtnfet l=6e-08 w=5e-07 $X=10200 $Y=6701 $D=616
M342 vss 148 147 vss hvtnfet l=6e-08 w=3e-07 $X=10200 $Y=7831 $D=616
M343 vss 148 149 vss hvtnfet l=6e-08 w=3e-07 $X=10200 $Y=43002 $D=616
M344 vss 149 150 vss hvtnfet l=6e-08 w=5e-07 $X=10200 $Y=43932 $D=616
M345 vss 150 t_pxbb_n<3> vss hvtnfet l=6e-08 w=1.285e-06 $X=10200 $Y=49512 $D=616
M346 160 129 vss vss hvtnfet l=6e-08 w=2.74e-07 $X=10246 $Y=13476 $D=616
M347 140 dwlb<1> 959 vss hvtnfet l=6e-08 w=4.11e-07 $X=10356 $Y=11276 $D=616
M348 141 dwlb<0> 960 vss hvtnfet l=6e-08 w=4.11e-07 $X=10356 $Y=39446 $D=616
M349 vss 153 124 vss hvtnfet l=6e-08 w=4e-07 $X=10406 $Y=32543 $D=616
M350 vss 142 dwlb<1> vss hvtnfet l=6e-08 w=3e-07 $X=10459 $Y=31098 $D=616
M351 vss 143 24 vss hvtnfet l=6e-08 w=3e-07 $X=10459 $Y=37457 $D=616
M352 b_pxbb_n<4> 156 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=10710 $Y=336 $D=616
M353 156 157 vss vss hvtnfet l=6e-08 w=5e-07 $X=10710 $Y=6701 $D=616
M354 157 105 vss vss hvtnfet l=6e-08 w=3e-07 $X=10710 $Y=7831 $D=616
M355 158 105 vss vss hvtnfet l=6e-08 w=3e-07 $X=10710 $Y=43002 $D=616
M356 159 158 vss vss hvtnfet l=6e-08 w=5e-07 $X=10710 $Y=43932 $D=616
M357 t_pxbb_n<4> 159 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=10710 $Y=49512 $D=616
M358 vss 132 133 vss hvtnfet l=6e-08 w=2.74e-07 $X=10846 $Y=13476 $D=616
M359 961 132 168 vss hvtnfet l=6e-08 w=5.49e-07 $X=10861 $Y=17417 $D=616
M360 962 133 169 vss hvtnfet l=6e-08 w=5.49e-07 $X=10861 $Y=18966 $D=616
M361 963 132 170 vss hvtnfet l=6e-08 w=5.49e-07 $X=10861 $Y=24337 $D=616
M362 964 133 171 vss hvtnfet l=6e-08 w=5.49e-07 $X=10861 $Y=25886 $D=616
M363 965 dwlb<1> 162 vss hvtnfet l=6e-08 w=4.11e-07 $X=10866 $Y=11276 $D=616
M364 966 dwlb<0> 163 vss hvtnfet l=6e-08 w=4.11e-07 $X=10866 $Y=39446 $D=616
M365 dwlb<1> 153 vss vss hvtnfet l=6e-08 w=3e-07 $X=10969 $Y=31098 $D=616
M366 24 153 vss vss hvtnfet l=6e-08 w=3e-07 $X=10969 $Y=37457 $D=616
M367 vss 156 b_pxbb_n<4> vss hvtnfet l=6e-08 w=1.285e-06 $X=10970 $Y=336 $D=616
M368 vss 157 156 vss hvtnfet l=6e-08 w=5e-07 $X=10970 $Y=6701 $D=616
M369 vss 105 157 vss hvtnfet l=6e-08 w=3e-07 $X=10970 $Y=7831 $D=616
M370 vss 105 158 vss hvtnfet l=6e-08 w=3e-07 $X=10970 $Y=43002 $D=616
M371 vss 158 159 vss hvtnfet l=6e-08 w=5e-07 $X=10970 $Y=43932 $D=616
M372 vss 159 t_pxbb_n<4> vss hvtnfet l=6e-08 w=1.285e-06 $X=10970 $Y=49512 $D=616
M373 132 ab<7> vss vss hvtnfet l=6e-08 w=2.74e-07 $X=11106 $Y=13476 $D=616
M374 153 154 vss vss hvtnfet l=6e-08 w=5e-07 $X=11106 $Y=32443 $D=616
M375 967 160 961 vss hvtnfet l=6e-08 w=5.49e-07 $X=11121 $Y=17417 $D=616
M376 968 160 962 vss hvtnfet l=6e-08 w=5.49e-07 $X=11121 $Y=18966 $D=616
M377 969 160 963 vss hvtnfet l=6e-08 w=5.49e-07 $X=11121 $Y=24337 $D=616
M378 970 160 964 vss hvtnfet l=6e-08 w=5.49e-07 $X=11121 $Y=25886 $D=616
M379 vss 155 965 vss hvtnfet l=6e-08 w=4.11e-07 $X=11126 $Y=11276 $D=616
M380 vss 155 966 vss hvtnfet l=6e-08 w=4.11e-07 $X=11126 $Y=39446 $D=616
M381 vss 153 dwlb<1> vss hvtnfet l=6e-08 w=3e-07 $X=11229 $Y=31098 $D=616
M382 vss 153 24 vss hvtnfet l=6e-08 w=3e-07 $X=11229 $Y=37457 $D=616
M383 971 121 967 vss hvtnfet l=6e-08 w=5.49e-07 $X=11381 $Y=17417 $D=616
M384 972 121 968 vss hvtnfet l=6e-08 w=5.49e-07 $X=11381 $Y=18966 $D=616
M385 973 122 969 vss hvtnfet l=6e-08 w=5.49e-07 $X=11381 $Y=24337 $D=616
M386 974 122 970 vss hvtnfet l=6e-08 w=5.49e-07 $X=11381 $Y=25886 $D=616
M387 b_pxbb_n<5> 164 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=11480 $Y=336 $D=616
M388 164 165 vss vss hvtnfet l=6e-08 w=5e-07 $X=11480 $Y=6701 $D=616
M389 165 106 vss vss hvtnfet l=6e-08 w=3e-07 $X=11480 $Y=7831 $D=616
M390 166 106 vss vss hvtnfet l=6e-08 w=3e-07 $X=11480 $Y=43002 $D=616
M391 167 166 vss vss hvtnfet l=6e-08 w=5e-07 $X=11480 $Y=43932 $D=616
M392 t_pxbb_n<5> 167 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=11480 $Y=49512 $D=616
M393 47 162 vss vss hvtnfet l=6e-08 w=2e-07 $X=11636 $Y=11276 $D=616
M394 50 163 vss vss hvtnfet l=6e-08 w=2e-07 $X=11636 $Y=39657 $D=616
M395 vss 43 971 vss hvtnfet l=6e-08 w=8.23e-07 $X=11651 $Y=17143 $D=616
M396 vss 43 972 vss hvtnfet l=6e-08 w=8.23e-07 $X=11651 $Y=18966 $D=616
M397 vss 43 973 vss hvtnfet l=6e-08 w=8.23e-07 $X=11651 $Y=24063 $D=616
M398 vss 43 974 vss hvtnfet l=6e-08 w=8.23e-07 $X=11651 $Y=25886 $D=616
M399 172 142 vss vss hvtnfet l=6e-08 w=2e-07 $X=11739 $Y=31098 $D=616
M400 vss 164 b_pxbb_n<5> vss hvtnfet l=6e-08 w=1.285e-06 $X=11740 $Y=336 $D=616
M401 vss 165 164 vss hvtnfet l=6e-08 w=5e-07 $X=11740 $Y=6701 $D=616
M402 vss 106 165 vss hvtnfet l=6e-08 w=3e-07 $X=11740 $Y=7831 $D=616
M403 vss 106 166 vss hvtnfet l=6e-08 w=3e-07 $X=11740 $Y=43002 $D=616
M404 vss 166 167 vss hvtnfet l=6e-08 w=5e-07 $X=11740 $Y=43932 $D=616
M405 vss 167 t_pxbb_n<5> vss hvtnfet l=6e-08 w=1.285e-06 $X=11740 $Y=49512 $D=616
M406 vss tm<0> dbl_pd_n<0> vss hvtnfet l=6e-08 w=2.14e-07 $X=11746 $Y=13361 $D=616
M407 dbl_pd_n<0> tm<0> vss vss hvtnfet l=6e-08 w=2.14e-07 $X=12006 $Y=13361 $D=616
M408 179 173 vss vss hvtnfet l=6e-08 w=2e-07 $X=12086 $Y=32533 $D=616
M409 vss 174 2 vss hvtnfet l=6e-08 w=2e-07 $X=12146 $Y=11276 $D=616
M410 177 168 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=12146 $Y=17812 $D=616
M411 178 169 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=12146 $Y=18983 $D=616
M412 137 170 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=12146 $Y=24732 $D=616
M413 148 171 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=12146 $Y=25903 $D=616
M414 vss 175 6 vss hvtnfet l=6e-08 w=2e-07 $X=12146 $Y=39657 $D=616
M415 975 33 168 vss hvtnfet l=6e-08 w=1.8e-07 $X=12161 $Y=17143 $D=616
M416 976 33 169 vss hvtnfet l=6e-08 w=1.8e-07 $X=12161 $Y=19609 $D=616
M417 977 33 170 vss hvtnfet l=6e-08 w=1.8e-07 $X=12161 $Y=24063 $D=616
M418 978 33 171 vss hvtnfet l=6e-08 w=1.8e-07 $X=12161 $Y=26529 $D=616
M419 vss 172 143 vss hvtnfet l=6e-08 w=6e-07 $X=12193 $Y=37037 $D=616
M420 b_pxbb_n<6> 180 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=12250 $Y=336 $D=616
M421 180 181 vss vss hvtnfet l=6e-08 w=5e-07 $X=12250 $Y=6701 $D=616
M422 181 177 vss vss hvtnfet l=6e-08 w=3e-07 $X=12250 $Y=7831 $D=616
M423 182 177 vss vss hvtnfet l=6e-08 w=3e-07 $X=12250 $Y=43002 $D=616
M424 183 182 vss vss hvtnfet l=6e-08 w=5e-07 $X=12250 $Y=43932 $D=616
M425 t_pxbb_n<6> 183 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=12250 $Y=49512 $D=616
M426 vss tm<0> dbl_pd_n<0> vss hvtnfet l=6e-08 w=2.14e-07 $X=12266 $Y=13361 $D=616
M427 vss 142 184 vss hvtnfet l=2.5e-07 w=3.5e-07 $X=12309 $Y=30853 $D=616
M428 vss 168 177 vss hvtnfet l=6e-08 w=1.37e-07 $X=12406 $Y=17812 $D=616
M429 vss 169 178 vss hvtnfet l=6e-08 w=1.37e-07 $X=12406 $Y=18983 $D=616
M430 vss 170 137 vss hvtnfet l=6e-08 w=1.37e-07 $X=12406 $Y=24732 $D=616
M431 vss 171 148 vss hvtnfet l=6e-08 w=1.37e-07 $X=12406 $Y=25903 $D=616
M432 vss 177 975 vss hvtnfet l=6e-08 w=1.8e-07 $X=12421 $Y=17143 $D=616
M433 vss 178 976 vss hvtnfet l=6e-08 w=1.8e-07 $X=12421 $Y=19609 $D=616
M434 vss 137 977 vss hvtnfet l=6e-08 w=1.8e-07 $X=12421 $Y=24063 $D=616
M435 vss 148 978 vss hvtnfet l=6e-08 w=1.8e-07 $X=12421 $Y=26529 $D=616
M436 vss 180 b_pxbb_n<6> vss hvtnfet l=6e-08 w=1.285e-06 $X=12510 $Y=336 $D=616
M437 vss 181 180 vss hvtnfet l=6e-08 w=5e-07 $X=12510 $Y=6701 $D=616
M438 vss 177 181 vss hvtnfet l=6e-08 w=3e-07 $X=12510 $Y=7831 $D=616
M439 vss 177 182 vss hvtnfet l=6e-08 w=3e-07 $X=12510 $Y=43002 $D=616
M440 vss 182 183 vss hvtnfet l=6e-08 w=5e-07 $X=12510 $Y=43932 $D=616
M441 vss 183 t_pxbb_n<6> vss hvtnfet l=6e-08 w=1.285e-06 $X=12510 $Y=49512 $D=616
M442 vss 179 186 vss hvtnfet l=6e-08 w=2e-07 $X=12596 $Y=32533 $D=616
M443 979 185 vss vss hvtnfet l=6e-08 w=4.11e-07 $X=12656 $Y=11276 $D=616
M444 980 185 vss vss hvtnfet l=6e-08 w=4.11e-07 $X=12656 $Y=39446 $D=616
M445 191 184 vss vss hvtnfet l=6e-08 w=3.5e-07 $X=12759 $Y=30853 $D=616
M446 vss 131 dbl_pd_n<2> vss hvtnfet l=6e-08 w=2.14e-07 $X=12776 $Y=13361 $D=616
M447 186 191 vss vss hvtnfet l=6e-08 w=2e-07 $X=12856 $Y=32533 $D=616
M448 174 dwlb<1> 979 vss hvtnfet l=6e-08 w=4.11e-07 $X=12916 $Y=11276 $D=616
M449 175 dwlb<0> 980 vss hvtnfet l=6e-08 w=4.11e-07 $X=12916 $Y=39446 $D=616
M450 981 187 vss vss hvtnfet l=6e-08 w=1.8e-07 $X=12931 $Y=17143 $D=616
M451 982 188 vss vss hvtnfet l=6e-08 w=1.8e-07 $X=12931 $Y=19609 $D=616
M452 983 189 vss vss hvtnfet l=6e-08 w=1.8e-07 $X=12931 $Y=24063 $D=616
M453 984 190 vss vss hvtnfet l=6e-08 w=1.8e-07 $X=12931 $Y=26529 $D=616
M454 187 192 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=12946 $Y=17812 $D=616
M455 188 193 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=12946 $Y=18983 $D=616
M456 189 194 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=12946 $Y=24732 $D=616
M457 190 195 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=12946 $Y=25903 $D=616
M458 vss 186 143 vss hvtnfet l=6e-08 w=6e-07 $X=12973 $Y=37037 $D=616
M459 b_pxbb_n<7> 196 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=13020 $Y=336 $D=616
M460 196 197 vss vss hvtnfet l=6e-08 w=5e-07 $X=13020 $Y=6701 $D=616
M461 197 178 vss vss hvtnfet l=6e-08 w=3e-07 $X=13020 $Y=7831 $D=616
M462 198 178 vss vss hvtnfet l=6e-08 w=3e-07 $X=13020 $Y=43002 $D=616
M463 199 198 vss vss hvtnfet l=6e-08 w=5e-07 $X=13020 $Y=43932 $D=616
M464 t_pxbb_n<7> 199 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=13020 $Y=49512 $D=616
M465 dbl_pd_n<2> 131 vss vss hvtnfet l=6e-08 w=2.14e-07 $X=13036 $Y=13361 $D=616
M466 192 33 981 vss hvtnfet l=6e-08 w=1.8e-07 $X=13191 $Y=17143 $D=616
M467 193 33 982 vss hvtnfet l=6e-08 w=1.8e-07 $X=13191 $Y=19609 $D=616
M468 194 33 983 vss hvtnfet l=6e-08 w=1.8e-07 $X=13191 $Y=24063 $D=616
M469 195 33 984 vss hvtnfet l=6e-08 w=1.8e-07 $X=13191 $Y=26529 $D=616
M470 vss 192 187 vss hvtnfet l=6e-08 w=1.37e-07 $X=13206 $Y=17812 $D=616
M471 vss 193 188 vss hvtnfet l=6e-08 w=1.37e-07 $X=13206 $Y=18983 $D=616
M472 vss 194 189 vss hvtnfet l=6e-08 w=1.37e-07 $X=13206 $Y=24732 $D=616
M473 vss 195 190 vss hvtnfet l=6e-08 w=1.37e-07 $X=13206 $Y=25903 $D=616
M474 vss 196 b_pxbb_n<7> vss hvtnfet l=6e-08 w=1.285e-06 $X=13280 $Y=336 $D=616
M475 vss 197 196 vss hvtnfet l=6e-08 w=5e-07 $X=13280 $Y=6701 $D=616
M476 vss 178 197 vss hvtnfet l=6e-08 w=3e-07 $X=13280 $Y=7831 $D=616
M477 vss 178 198 vss hvtnfet l=6e-08 w=3e-07 $X=13280 $Y=43002 $D=616
M478 vss 198 199 vss hvtnfet l=6e-08 w=5e-07 $X=13280 $Y=43932 $D=616
M479 vss 199 t_pxbb_n<7> vss hvtnfet l=6e-08 w=1.285e-06 $X=13280 $Y=49512 $D=616
M480 vss 131 dbl_pd_n<2> vss hvtnfet l=6e-08 w=2.14e-07 $X=13296 $Y=13361 $D=616
M481 vss 191 202 vss hvtnfet l=2.5e-07 w=3.5e-07 $X=13429 $Y=30853 $D=616
M482 vss tm<7> 203 vss hvtnfet l=6e-08 w=2e-07 $X=13432 $Y=32533 $D=616
M483 985 43 vss vss hvtnfet l=6e-08 w=8.23e-07 $X=13701 $Y=17143 $D=616
M484 986 43 vss vss hvtnfet l=6e-08 w=8.23e-07 $X=13701 $Y=18966 $D=616
M485 987 43 vss vss hvtnfet l=6e-08 w=8.23e-07 $X=13701 $Y=24063 $D=616
M486 988 43 vss vss hvtnfet l=6e-08 w=8.23e-07 $X=13701 $Y=25886 $D=616
M487 vss 200 143 vss hvtnfet l=6e-08 w=6e-07 $X=13753 $Y=37037 $D=616
M488 b_pxcb_n<0> 206 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=13790 $Y=336 $D=616
M489 206 207 vss vss hvtnfet l=6e-08 w=5e-07 $X=13790 $Y=6701 $D=616
M490 207 189 vss vss hvtnfet l=6e-08 w=3e-07 $X=13790 $Y=7831 $D=616
M491 208 189 vss vss hvtnfet l=6e-08 w=3e-07 $X=13790 $Y=43002 $D=616
M492 209 208 vss vss hvtnfet l=6e-08 w=5e-07 $X=13790 $Y=43932 $D=616
M493 t_pxcb_n<0> 209 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=13790 $Y=49512 $D=616
M494 211 202 vss vss hvtnfet l=6e-08 w=3.5e-07 $X=13879 $Y=30853 $D=616
M495 vss 205 204 vss hvtnfet l=6e-08 w=2.74e-07 $X=13936 $Y=13476 $D=616
M496 vss 203 200 vss hvtnfet l=6e-08 w=2e-07 $X=13942 $Y=32533 $D=616
M497 989 204 985 vss hvtnfet l=6e-08 w=5.49e-07 $X=13971 $Y=17417 $D=616
M498 990 204 986 vss hvtnfet l=6e-08 w=5.49e-07 $X=13971 $Y=18966 $D=616
M499 991 205 987 vss hvtnfet l=6e-08 w=5.49e-07 $X=13971 $Y=24337 $D=616
M500 992 205 988 vss hvtnfet l=6e-08 w=5.49e-07 $X=13971 $Y=25886 $D=616
M501 vss 206 b_pxcb_n<0> vss hvtnfet l=6e-08 w=1.285e-06 $X=14050 $Y=336 $D=616
M502 vss 207 206 vss hvtnfet l=6e-08 w=5e-07 $X=14050 $Y=6701 $D=616
M503 vss 189 207 vss hvtnfet l=6e-08 w=3e-07 $X=14050 $Y=7831 $D=616
M504 vss 189 208 vss hvtnfet l=6e-08 w=3e-07 $X=14050 $Y=43002 $D=616
M505 vss 208 209 vss hvtnfet l=6e-08 w=5e-07 $X=14050 $Y=43932 $D=616
M506 vss 209 t_pxcb_n<0> vss hvtnfet l=6e-08 w=1.285e-06 $X=14050 $Y=49512 $D=616
M507 200 211 vss vss hvtnfet l=6e-08 w=2e-07 $X=14202 $Y=32533 $D=616
M508 993 dwlb<1> 216 vss hvtnfet l=6e-08 w=4.11e-07 $X=14216 $Y=11276 $D=616
M509 994 dwlb<0> 217 vss hvtnfet l=6e-08 w=4.11e-07 $X=14216 $Y=39446 $D=616
M510 995 210 989 vss hvtnfet l=6e-08 w=5.49e-07 $X=14231 $Y=17417 $D=616
M511 996 210 990 vss hvtnfet l=6e-08 w=5.49e-07 $X=14231 $Y=18966 $D=616
M512 997 210 991 vss hvtnfet l=6e-08 w=5.49e-07 $X=14231 $Y=24337 $D=616
M513 998 210 992 vss hvtnfet l=6e-08 w=5.49e-07 $X=14231 $Y=25886 $D=616
M514 205 ab<12> vss vss hvtnfet l=6e-08 w=2.74e-07 $X=14446 $Y=13476 $D=616
M515 vss 212 993 vss hvtnfet l=6e-08 w=4.11e-07 $X=14476 $Y=11276 $D=616
M516 vss 212 994 vss hvtnfet l=6e-08 w=4.11e-07 $X=14476 $Y=39446 $D=616
M517 192 213 995 vss hvtnfet l=6e-08 w=5.49e-07 $X=14491 $Y=17417 $D=616
M518 193 214 996 vss hvtnfet l=6e-08 w=5.49e-07 $X=14491 $Y=18966 $D=616
M519 194 213 997 vss hvtnfet l=6e-08 w=5.49e-07 $X=14491 $Y=24337 $D=616
M520 195 214 998 vss hvtnfet l=6e-08 w=5.49e-07 $X=14491 $Y=25886 $D=616
M521 b_pxcb_n<1> 218 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=14560 $Y=336 $D=616
M522 218 219 vss vss hvtnfet l=6e-08 w=5e-07 $X=14560 $Y=6701 $D=616
M523 219 190 vss vss hvtnfet l=6e-08 w=3e-07 $X=14560 $Y=7831 $D=616
M524 220 190 vss vss hvtnfet l=6e-08 w=3e-07 $X=14560 $Y=43002 $D=616
M525 221 220 vss vss hvtnfet l=6e-08 w=5e-07 $X=14560 $Y=43932 $D=616
M526 t_pxcb_n<1> 221 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=14560 $Y=49512 $D=616
M527 vss 123 624 vss hvtnfet l=6e-08 w=6e-07 $X=14796 $Y=30668 $D=616
M528 vss 218 b_pxcb_n<1> vss hvtnfet l=6e-08 w=1.285e-06 $X=14820 $Y=336 $D=616
M529 vss 219 218 vss hvtnfet l=6e-08 w=5e-07 $X=14820 $Y=6701 $D=616
M530 vss 190 219 vss hvtnfet l=6e-08 w=3e-07 $X=14820 $Y=7831 $D=616
M531 vss 190 220 vss hvtnfet l=6e-08 w=3e-07 $X=14820 $Y=43002 $D=616
M532 vss 220 221 vss hvtnfet l=6e-08 w=5e-07 $X=14820 $Y=43932 $D=616
M533 vss 221 t_pxcb_n<1> vss hvtnfet l=6e-08 w=1.285e-06 $X=14820 $Y=49512 $D=616
M534 vss 72 58 vss hvtnfet l=6e-08 w=2e-07 $X=14872 $Y=37045 $D=616
M535 48 216 vss vss hvtnfet l=6e-08 w=2e-07 $X=14986 $Y=11276 $D=616
M536 49 217 vss vss hvtnfet l=6e-08 w=2e-07 $X=14986 $Y=39657 $D=616
M537 vss 43 33 vss hvtnfet l=6e-08 w=7e-07 $X=15316 $Y=30668 $D=616
M538 b_pxcb_n<2> 223 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=15330 $Y=336 $D=616
M539 223 224 vss vss hvtnfet l=6e-08 w=5e-07 $X=15330 $Y=6701 $D=616
M540 224 225 vss vss hvtnfet l=6e-08 w=3e-07 $X=15330 $Y=7831 $D=616
M541 226 225 vss vss hvtnfet l=6e-08 w=3e-07 $X=15330 $Y=43002 $D=616
M542 227 226 vss vss hvtnfet l=6e-08 w=5e-07 $X=15330 $Y=43932 $D=616
M543 t_pxcb_n<2> 227 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=15330 $Y=49512 $D=616
M544 629 229 vss vss hvtnfet l=6e-08 w=4e-07 $X=15382 $Y=37045 $D=616
M545 vss ab<11> 210 vss hvtnfet l=6e-08 w=2.74e-07 $X=15456 $Y=13476 $D=616
M546 33 43 vss vss hvtnfet l=6e-08 w=7e-07 $X=15576 $Y=30668 $D=616
M547 vss 223 b_pxcb_n<2> vss hvtnfet l=6e-08 w=1.285e-06 $X=15590 $Y=336 $D=616
M548 vss 224 223 vss hvtnfet l=6e-08 w=5e-07 $X=15590 $Y=6701 $D=616
M549 vss 225 224 vss hvtnfet l=6e-08 w=3e-07 $X=15590 $Y=7831 $D=616
M550 vss 225 226 vss hvtnfet l=6e-08 w=3e-07 $X=15590 $Y=43002 $D=616
M551 vss 226 227 vss hvtnfet l=6e-08 w=5e-07 $X=15590 $Y=43932 $D=616
M552 vss 227 t_pxcb_n<2> vss hvtnfet l=6e-08 w=1.285e-06 $X=15590 $Y=49512 $D=616
M553 vss 228 231 vss hvtnfet l=6e-08 w=2.1e-07 $X=15621 $Y=32688 $D=616
M554 72 172 629 vss hvtnfet l=6e-08 w=4e-07 $X=15642 $Y=37045 $D=616
M555 240 210 vss vss hvtnfet l=6e-08 w=2.74e-07 $X=15716 $Y=13476 $D=616
M556 631 tm<0> vss vss hvtnfet l=6e-08 w=2.74e-07 $X=15880 $Y=39358 $D=616
M557 630 131 vss vss hvtnfet l=6e-08 w=2.1e-07 $X=15881 $Y=32688 $D=616
M558 vss tm<3> 242 vss hvtnfet l=7e-08 w=3.2e-07 $X=16057 $Y=11276 $D=616
M559 b_pxcb_n<3> 235 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=16100 $Y=336 $D=616
M560 235 236 vss vss hvtnfet l=6e-08 w=5e-07 $X=16100 $Y=6701 $D=616
M561 236 237 vss vss hvtnfet l=6e-08 w=3e-07 $X=16100 $Y=7831 $D=616
M562 238 237 vss vss hvtnfet l=6e-08 w=3e-07 $X=16100 $Y=43002 $D=616
M563 239 238 vss vss hvtnfet l=6e-08 w=5e-07 $X=16100 $Y=43932 $D=616
M564 t_pxcb_n<3> 239 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=16100 $Y=49512 $D=616
M565 228 231 630 vss hvtnfet l=6e-08 w=2.1e-07 $X=16141 $Y=32688 $D=616
M566 vss 213 214 vss hvtnfet l=6e-08 w=2.74e-07 $X=16316 $Y=13476 $D=616
M567 635 232 vss vss hvtnfet l=6e-08 w=3.2e-07 $X=16322 $Y=37277 $D=616
M568 243 tm<4> vss vss hvtnfet l=7e-08 w=3.2e-07 $X=16327 $Y=11276 $D=616
M569 999 213 249 vss hvtnfet l=6e-08 w=5.49e-07 $X=16331 $Y=17417 $D=616
M570 1000 214 250 vss hvtnfet l=6e-08 w=5.49e-07 $X=16331 $Y=18966 $D=616
M571 1001 213 251 vss hvtnfet l=6e-08 w=5.49e-07 $X=16331 $Y=24337 $D=616
M572 1002 214 252 vss hvtnfet l=6e-08 w=5.49e-07 $X=16331 $Y=25886 $D=616
M573 vss 123 644 vss hvtnfet l=6e-08 w=6e-07 $X=16346 $Y=30668 $D=616
M574 vss 235 b_pxcb_n<3> vss hvtnfet l=6e-08 w=1.285e-06 $X=16360 $Y=336 $D=616
M575 vss 236 235 vss hvtnfet l=6e-08 w=5e-07 $X=16360 $Y=6701 $D=616
M576 vss 237 236 vss hvtnfet l=6e-08 w=3e-07 $X=16360 $Y=7831 $D=616
M577 vss 237 238 vss hvtnfet l=6e-08 w=3e-07 $X=16360 $Y=43002 $D=616
M578 vss 238 239 vss hvtnfet l=6e-08 w=5e-07 $X=16360 $Y=43932 $D=616
M579 vss 239 t_pxcb_n<3> vss hvtnfet l=6e-08 w=1.285e-06 $X=16360 $Y=49512 $D=616
M580 636 123 228 vss hvtnfet l=6e-08 w=3.2e-07 $X=16401 $Y=32578 $D=616
M581 213 ab<10> vss vss hvtnfet l=6e-08 w=2.74e-07 $X=16576 $Y=13476 $D=616
M582 229 142 635 vss hvtnfet l=6e-08 w=3.2e-07 $X=16582 $Y=37277 $D=616
M583 1003 240 999 vss hvtnfet l=6e-08 w=5.49e-07 $X=16591 $Y=17417 $D=616
M584 1004 240 1000 vss hvtnfet l=6e-08 w=5.49e-07 $X=16591 $Y=18966 $D=616
M585 1005 240 1001 vss hvtnfet l=6e-08 w=5.49e-07 $X=16591 $Y=24337 $D=616
M586 1006 240 1002 vss hvtnfet l=6e-08 w=5.49e-07 $X=16591 $Y=25886 $D=616
M587 644 123 vss vss hvtnfet l=6e-08 w=6e-07 $X=16606 $Y=30668 $D=616
M588 vss 123 636 vss hvtnfet l=6e-08 w=3.2e-07 $X=16661 $Y=32578 $D=616
M589 637 tm<6> vss vss hvtnfet l=6e-08 w=2.74e-07 $X=16680 $Y=39358 $D=616
M590 638 244 229 vss hvtnfet l=6e-08 w=2.1e-07 $X=16842 $Y=37277 $D=616
M591 vss 243 643 vss hvtnfet l=6e-08 w=4.8e-07 $X=16847 $Y=11276 $D=616
M592 1007 204 1003 vss hvtnfet l=6e-08 w=5.49e-07 $X=16851 $Y=17417 $D=616
M593 1008 204 1004 vss hvtnfet l=6e-08 w=5.49e-07 $X=16851 $Y=18966 $D=616
M594 1009 205 1005 vss hvtnfet l=6e-08 w=5.49e-07 $X=16851 $Y=24337 $D=616
M595 1010 205 1006 vss hvtnfet l=6e-08 w=5.49e-07 $X=16851 $Y=25886 $D=616
M596 642 123 644 vss hvtnfet l=6e-08 w=6e-07 $X=16866 $Y=30668 $D=616
M597 b_pxcb_n<4> 245 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=16870 $Y=336 $D=616
M598 245 246 vss vss hvtnfet l=6e-08 w=5e-07 $X=16870 $Y=6701 $D=616
M599 246 187 vss vss hvtnfet l=6e-08 w=3e-07 $X=16870 $Y=7831 $D=616
M600 247 187 vss vss hvtnfet l=6e-08 w=3e-07 $X=16870 $Y=43002 $D=616
M601 248 247 vss vss hvtnfet l=6e-08 w=5e-07 $X=16870 $Y=43932 $D=616
M602 t_pxcb_n<4> 248 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=16870 $Y=49512 $D=616
M603 vss 172 638 vss hvtnfet l=6e-08 w=2.1e-07 $X=17102 $Y=37277 $D=616
M604 643 242 vss vss hvtnfet l=6e-08 w=4.8e-07 $X=17107 $Y=11276 $D=616
M605 vss 43 1007 vss hvtnfet l=6e-08 w=8.23e-07 $X=17121 $Y=17143 $D=616
M606 vss 43 1008 vss hvtnfet l=6e-08 w=8.23e-07 $X=17121 $Y=18966 $D=616
M607 vss 43 1009 vss hvtnfet l=6e-08 w=8.23e-07 $X=17121 $Y=24063 $D=616
M608 vss 43 1010 vss hvtnfet l=6e-08 w=8.23e-07 $X=17121 $Y=25886 $D=616
M609 644 123 642 vss hvtnfet l=6e-08 w=6e-07 $X=17126 $Y=30668 $D=616
M610 vss 245 b_pxcb_n<4> vss hvtnfet l=6e-08 w=1.285e-06 $X=17130 $Y=336 $D=616
M611 vss 246 245 vss hvtnfet l=6e-08 w=5e-07 $X=17130 $Y=6701 $D=616
M612 vss 187 246 vss hvtnfet l=6e-08 w=3e-07 $X=17130 $Y=7831 $D=616
M613 vss 187 247 vss hvtnfet l=6e-08 w=3e-07 $X=17130 $Y=43002 $D=616
M614 vss 247 248 vss hvtnfet l=6e-08 w=5e-07 $X=17130 $Y=43932 $D=616
M615 vss 248 t_pxcb_n<4> vss hvtnfet l=6e-08 w=1.285e-06 $X=17130 $Y=49512 $D=616
M616 244 229 vss vss hvtnfet l=6e-08 w=2.1e-07 $X=17362 $Y=37277 $D=616
M617 253 249 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=17616 $Y=17812 $D=616
M618 254 250 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=17616 $Y=18983 $D=616
M619 225 251 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=17616 $Y=24732 $D=616
M620 237 252 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=17616 $Y=25903 $D=616
M621 647 242 vss vss hvtnfet l=6e-08 w=4.8e-07 $X=17617 $Y=11276 $D=616
M622 1011 33 249 vss hvtnfet l=6e-08 w=1.8e-07 $X=17631 $Y=17143 $D=616
M623 1012 33 250 vss hvtnfet l=6e-08 w=1.8e-07 $X=17631 $Y=19609 $D=616
M624 1013 33 251 vss hvtnfet l=6e-08 w=1.8e-07 $X=17631 $Y=24063 $D=616
M625 1014 33 252 vss hvtnfet l=6e-08 w=1.8e-07 $X=17631 $Y=26529 $D=616
M626 b_pxcb_n<5> 255 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=17640 $Y=336 $D=616
M627 255 256 vss vss hvtnfet l=6e-08 w=5e-07 $X=17640 $Y=6701 $D=616
M628 256 188 vss vss hvtnfet l=6e-08 w=3e-07 $X=17640 $Y=7831 $D=616
M629 257 188 vss vss hvtnfet l=6e-08 w=3e-07 $X=17640 $Y=43002 $D=616
M630 258 257 vss vss hvtnfet l=6e-08 w=5e-07 $X=17640 $Y=43932 $D=616
M631 t_pxcb_n<5> 258 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=17640 $Y=49512 $D=616
M632 23 clkb vss vss hvtnfet l=6e-08 w=4.5e-07 $X=17646 $Y=30668 $D=616
M633 vss 249 253 vss hvtnfet l=6e-08 w=1.37e-07 $X=17876 $Y=17812 $D=616
M634 vss 250 254 vss hvtnfet l=6e-08 w=1.37e-07 $X=17876 $Y=18983 $D=616
M635 vss 251 225 vss hvtnfet l=6e-08 w=1.37e-07 $X=17876 $Y=24732 $D=616
M636 vss 252 237 vss hvtnfet l=6e-08 w=1.37e-07 $X=17876 $Y=25903 $D=616
M637 vss tm<4> 647 vss hvtnfet l=6e-08 w=4.8e-07 $X=17877 $Y=11276 $D=616
M638 vss 253 1011 vss hvtnfet l=6e-08 w=1.8e-07 $X=17891 $Y=17143 $D=616
M639 vss 254 1012 vss hvtnfet l=6e-08 w=1.8e-07 $X=17891 $Y=19609 $D=616
M640 vss 225 1013 vss hvtnfet l=6e-08 w=1.8e-07 $X=17891 $Y=24063 $D=616
M641 vss 237 1014 vss hvtnfet l=6e-08 w=1.8e-07 $X=17891 $Y=26529 $D=616
M642 vss 255 b_pxcb_n<5> vss hvtnfet l=6e-08 w=1.285e-06 $X=17900 $Y=336 $D=616
M643 vss 256 255 vss hvtnfet l=6e-08 w=5e-07 $X=17900 $Y=6701 $D=616
M644 vss 188 256 vss hvtnfet l=6e-08 w=3e-07 $X=17900 $Y=7831 $D=616
M645 vss 188 257 vss hvtnfet l=6e-08 w=3e-07 $X=17900 $Y=43002 $D=616
M646 vss 257 258 vss hvtnfet l=6e-08 w=5e-07 $X=17900 $Y=43932 $D=616
M647 vss 258 t_pxcb_n<5> vss hvtnfet l=6e-08 w=1.285e-06 $X=17900 $Y=49512 $D=616
M648 vss 260 273 vss hvtnfet l=6e-08 w=2.74e-07 $X=18106 $Y=13476 $D=616
M649 vss wenb 232 vss hvtnfet l=6e-08 w=2e-07 $X=18366 $Y=37147 $D=616
M650 648 tm<4> vss vss hvtnfet l=6e-08 w=4.8e-07 $X=18387 $Y=11276 $D=616
M651 b_pxcb_n<6> 265 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=18410 $Y=336 $D=616
M652 265 266 vss vss hvtnfet l=6e-08 w=5e-07 $X=18410 $Y=6701 $D=616
M653 266 253 vss vss hvtnfet l=6e-08 w=3e-07 $X=18410 $Y=7831 $D=616
M654 267 253 vss vss hvtnfet l=6e-08 w=3e-07 $X=18410 $Y=43002 $D=616
M655 268 267 vss vss hvtnfet l=6e-08 w=5e-07 $X=18410 $Y=43932 $D=616
M656 t_pxcb_n<6> 268 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=18410 $Y=49512 $D=616
M657 651 ab<4> vss vss hvtnfet l=6e-08 w=3.2e-07 $X=18460 $Y=30918 $D=616
M658 652 wenb vss vss hvtnfet l=6e-08 w=3.2e-07 $X=18460 $Y=32578 $D=616
M659 vss tm<2> 173 vss hvtnfet l=6e-08 w=2.74e-07 $X=18510 $Y=39358 $D=616
M660 260 ab<1> vss vss hvtnfet l=6e-08 w=2.74e-07 $X=18616 $Y=13476 $D=616
M661 232 264 vss vss hvtnfet l=6e-08 w=2e-07 $X=18626 $Y=37147 $D=616
M662 vss tm<3> 648 vss hvtnfet l=6e-08 w=4.8e-07 $X=18647 $Y=11276 $D=616
M663 vss 265 b_pxcb_n<6> vss hvtnfet l=6e-08 w=1.285e-06 $X=18670 $Y=336 $D=616
M664 vss 266 265 vss hvtnfet l=6e-08 w=5e-07 $X=18670 $Y=6701 $D=616
M665 vss 253 266 vss hvtnfet l=6e-08 w=3e-07 $X=18670 $Y=7831 $D=616
M666 vss 253 267 vss hvtnfet l=6e-08 w=3e-07 $X=18670 $Y=43002 $D=616
M667 vss 267 268 vss hvtnfet l=6e-08 w=5e-07 $X=18670 $Y=43932 $D=616
M668 vss 268 t_pxcb_n<6> vss hvtnfet l=6e-08 w=1.285e-06 $X=18670 $Y=49512 $D=616
M669 154 23 651 vss hvtnfet l=6e-08 w=3.2e-07 $X=18720 $Y=30918 $D=616
M670 274 23 652 vss hvtnfet l=6e-08 w=3.2e-07 $X=18720 $Y=32578 $D=616
M671 1015 269 280 vss hvtnfet l=6e-08 w=5.49e-07 $X=18911 $Y=17143 $D=616
M672 1016 270 281 vss hvtnfet l=6e-08 w=5.49e-07 $X=18911 $Y=19240 $D=616
M673 1017 269 282 vss hvtnfet l=6e-08 w=5.49e-07 $X=18911 $Y=24063 $D=616
M674 1018 270 283 vss hvtnfet l=6e-08 w=5.49e-07 $X=18911 $Y=26160 $D=616
M675 653 271 154 vss hvtnfet l=6e-08 w=2.1e-07 $X=18980 $Y=30918 $D=616
M676 654 272 274 vss hvtnfet l=6e-08 w=2.1e-07 $X=18980 $Y=32688 $D=616
M677 vss 270 269 vss hvtnfet l=6e-08 w=2.74e-07 $X=19126 $Y=13476 $D=616
M678 659 tm<3> vss vss hvtnfet l=6e-08 w=4.8e-07 $X=19157 $Y=11276 $D=616
M679 1019 273 1015 vss hvtnfet l=6e-08 w=5.49e-07 $X=19171 $Y=17143 $D=616
M680 1020 273 1016 vss hvtnfet l=6e-08 w=5.49e-07 $X=19171 $Y=19240 $D=616
M681 1021 260 1017 vss hvtnfet l=6e-08 w=5.49e-07 $X=19171 $Y=24063 $D=616
M682 1022 260 1018 vss hvtnfet l=6e-08 w=5.49e-07 $X=19171 $Y=26160 $D=616
M683 b_pxcb_n<7> 275 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=19180 $Y=336 $D=616
M684 275 276 vss vss hvtnfet l=6e-08 w=5e-07 $X=19180 $Y=6701 $D=616
M685 276 254 vss vss hvtnfet l=6e-08 w=3e-07 $X=19180 $Y=7831 $D=616
M686 277 254 vss vss hvtnfet l=6e-08 w=3e-07 $X=19180 $Y=43002 $D=616
M687 278 277 vss vss hvtnfet l=6e-08 w=5e-07 $X=19180 $Y=43932 $D=616
M688 t_pxcb_n<7> 278 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=19180 $Y=49512 $D=616
M689 vss clkb 653 vss hvtnfet l=6e-08 w=2.1e-07 $X=19240 $Y=30918 $D=616
M690 vss clkb 654 vss hvtnfet l=6e-08 w=2.1e-07 $X=19240 $Y=32688 $D=616
M691 vss 243 659 vss hvtnfet l=6e-08 w=4.8e-07 $X=19417 $Y=11276 $D=616
M692 vss 275 b_pxcb_n<7> vss hvtnfet l=6e-08 w=1.285e-06 $X=19440 $Y=336 $D=616
M693 vss 276 275 vss hvtnfet l=6e-08 w=5e-07 $X=19440 $Y=6701 $D=616
M694 vss 254 276 vss hvtnfet l=6e-08 w=3e-07 $X=19440 $Y=7831 $D=616
M695 vss 254 277 vss hvtnfet l=6e-08 w=3e-07 $X=19440 $Y=43002 $D=616
M696 vss 277 278 vss hvtnfet l=6e-08 w=5e-07 $X=19440 $Y=43932 $D=616
M697 vss 278 t_pxcb_n<7> vss hvtnfet l=6e-08 w=1.285e-06 $X=19440 $Y=49512 $D=616
M698 vss 43 1019 vss hvtnfet l=6e-08 w=8.23e-07 $X=19441 $Y=17143 $D=616
M699 vss 43 1020 vss hvtnfet l=6e-08 w=8.23e-07 $X=19441 $Y=18966 $D=616
M700 vss 43 1021 vss hvtnfet l=6e-08 w=8.23e-07 $X=19441 $Y=24063 $D=616
M701 vss 43 1022 vss hvtnfet l=6e-08 w=8.23e-07 $X=19441 $Y=25886 $D=616
M702 271 154 vss vss hvtnfet l=6e-08 w=2.1e-07 $X=19500 $Y=30918 $D=616
M703 272 274 vss vss hvtnfet l=6e-08 w=2.1e-07 $X=19500 $Y=32688 $D=616
M704 270 ab<0> vss vss hvtnfet l=6e-08 w=2.74e-07 $X=19636 $Y=13476 $D=616
M705 vss 15 r_saeb_n vss hvtnfet l=6e-08 w=8.58e-07 $X=19675 $Y=37027 $D=616
M706 r_saeb_n 15 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=19935 $Y=37027 $D=616
M707 1023 33 280 vss hvtnfet l=6e-08 w=1.8e-07 $X=19951 $Y=17143 $D=616
M708 212 280 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=19951 $Y=17812 $D=616
M709 185 281 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=19951 $Y=18983 $D=616
M710 1024 33 281 vss hvtnfet l=6e-08 w=1.8e-07 $X=19951 $Y=19609 $D=616
M711 1025 33 282 vss hvtnfet l=6e-08 w=1.8e-07 $X=19951 $Y=24063 $D=616
M712 155 282 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=19951 $Y=24732 $D=616
M713 145 283 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=19951 $Y=25903 $D=616
M714 1026 33 283 vss hvtnfet l=6e-08 w=1.8e-07 $X=19951 $Y=26529 $D=616
M715 vss 11 rb_cb<0> vss hvtnfet l=6e-08 w=8.58e-07 $X=20195 $Y=328 $D=616
M716 vss 12 rb_cb<2> vss hvtnfet l=6e-08 w=8.58e-07 $X=20195 $Y=5316 $D=616
M717 vss 13 rb_mb<0> vss hvtnfet l=6e-08 w=8.58e-07 $X=20195 $Y=6788 $D=616
M718 vss 14 rb_mb<2> vss hvtnfet l=6e-08 w=8.58e-07 $X=20195 $Y=11776 $D=616
M719 vss 15 r_saeb_n vss hvtnfet l=6e-08 w=8.58e-07 $X=20195 $Y=37027 $D=616
M720 vss 16 rt_mb<2> vss hvtnfet l=6e-08 w=8.58e-07 $X=20195 $Y=38499 $D=616
M721 vss 17 rt_mb<0> vss hvtnfet l=6e-08 w=8.58e-07 $X=20195 $Y=43487 $D=616
M722 vss 18 rt_cb<2> vss hvtnfet l=6e-08 w=8.58e-07 $X=20195 $Y=44959 $D=616
M723 vss 19 rt_cb<0> vss hvtnfet l=6e-08 w=8.58e-07 $X=20195 $Y=49947 $D=616
M724 vss 212 1023 vss hvtnfet l=6e-08 w=1.8e-07 $X=20211 $Y=17143 $D=616
M725 vss 280 212 vss hvtnfet l=6e-08 w=1.37e-07 $X=20211 $Y=17812 $D=616
M726 vss 281 185 vss hvtnfet l=6e-08 w=1.37e-07 $X=20211 $Y=18983 $D=616
M727 vss 185 1024 vss hvtnfet l=6e-08 w=1.8e-07 $X=20211 $Y=19609 $D=616
M728 vss 155 1025 vss hvtnfet l=6e-08 w=1.8e-07 $X=20211 $Y=24063 $D=616
M729 vss 282 155 vss hvtnfet l=6e-08 w=1.37e-07 $X=20211 $Y=24732 $D=616
M730 vss 283 145 vss hvtnfet l=6e-08 w=1.37e-07 $X=20211 $Y=25903 $D=616
M731 vss 145 1026 vss hvtnfet l=6e-08 w=1.8e-07 $X=20211 $Y=26529 $D=616
M732 rb_cb<0> 11 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=20455 $Y=328 $D=616
M733 rb_cb<2> 12 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=20455 $Y=5316 $D=616
M734 rb_mb<0> 13 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=20455 $Y=6788 $D=616
M735 rb_mb<2> 14 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=20455 $Y=11776 $D=616
M736 r_saeb_n 15 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=20455 $Y=37027 $D=616
M737 rt_mb<2> 16 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=20455 $Y=38499 $D=616
M738 rt_mb<0> 17 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=20455 $Y=43487 $D=616
M739 rt_cb<2> 18 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=20455 $Y=44959 $D=616
M740 rt_cb<0> 19 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=20455 $Y=49947 $D=616
M741 vss 11 rb_cb<0> vss hvtnfet l=6e-08 w=8.58e-07 $X=20715 $Y=328 $D=616
M742 vss 12 rb_cb<2> vss hvtnfet l=6e-08 w=8.58e-07 $X=20715 $Y=5316 $D=616
M743 vss 13 rb_mb<0> vss hvtnfet l=6e-08 w=8.58e-07 $X=20715 $Y=6788 $D=616
M744 vss 14 rb_mb<2> vss hvtnfet l=6e-08 w=8.58e-07 $X=20715 $Y=11776 $D=616
M745 vss 15 r_saeb_n vss hvtnfet l=6e-08 w=8.58e-07 $X=20715 $Y=37027 $D=616
M746 vss 16 rt_mb<2> vss hvtnfet l=6e-08 w=8.58e-07 $X=20715 $Y=38499 $D=616
M747 vss 17 rt_mb<0> vss hvtnfet l=6e-08 w=8.58e-07 $X=20715 $Y=43487 $D=616
M748 vss 18 rt_cb<2> vss hvtnfet l=6e-08 w=8.58e-07 $X=20715 $Y=44959 $D=616
M749 vss 19 rt_cb<0> vss hvtnfet l=6e-08 w=8.58e-07 $X=20715 $Y=49947 $D=616
M750 10 274 vss vss hvtnfet l=6e-08 w=6e-07 $X=20725 $Y=30899 $D=616
M751 rb_cb<1> 34 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=20975 $Y=328 $D=616
M752 rb_cb<3> 35 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=20975 $Y=5316 $D=616
M753 rb_mb<1> 36 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=20975 $Y=6788 $D=616
M754 rb_mb<3> 37 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=20975 $Y=11776 $D=616
M755 r_clk_dqb 8 vss vss hvtnfet l=6e-08 w=1.26e-06 $X=20975 $Y=22041 $D=616
M756 r_clk_dqb_n 9 vss vss hvtnfet l=6e-08 w=1.26e-06 $X=20975 $Y=29007 $D=616
M757 r_sa_preb_n 51 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=20975 $Y=37027 $D=616
M758 rt_mb<3> 39 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=20975 $Y=38499 $D=616
M759 rt_mb<1> 40 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=20975 $Y=43487 $D=616
M760 rt_cb<3> 41 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=20975 $Y=44959 $D=616
M761 rt_cb<1> 42 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=20975 $Y=49947 $D=616
M762 vss 34 rb_cb<1> vss hvtnfet l=6e-08 w=8.58e-07 $X=21235 $Y=328 $D=616
M763 vss 35 rb_cb<3> vss hvtnfet l=6e-08 w=8.58e-07 $X=21235 $Y=5316 $D=616
M764 vss 36 rb_mb<1> vss hvtnfet l=6e-08 w=8.58e-07 $X=21235 $Y=6788 $D=616
M765 vss 37 rb_mb<3> vss hvtnfet l=6e-08 w=8.58e-07 $X=21235 $Y=11776 $D=616
M766 rb_tm_preb_n 20 vss vss hvtnfet l=6e-08 w=1.287e-06 $X=21235 $Y=13280 $D=616
M767 rt_tm_preb_n 21 vss vss hvtnfet l=6e-08 w=1.287e-06 $X=21235 $Y=20124 $D=616
M768 vss 8 r_clk_dqb vss hvtnfet l=6e-08 w=1.26e-06 $X=21235 $Y=22041 $D=616
M769 vss 9 r_clk_dqb_n vss hvtnfet l=6e-08 w=1.26e-06 $X=21235 $Y=29007 $D=616
M770 r_lweb 10 vss vss hvtnfet l=6e-08 w=1.287e-06 $X=21235 $Y=30897 $D=616
M771 vss 51 r_sa_preb_n vss hvtnfet l=6e-08 w=8.58e-07 $X=21235 $Y=37027 $D=616
M772 vss 39 rt_mb<3> vss hvtnfet l=6e-08 w=8.58e-07 $X=21235 $Y=38499 $D=616
M773 vss 40 rt_mb<1> vss hvtnfet l=6e-08 w=8.58e-07 $X=21235 $Y=43487 $D=616
M774 vss 41 rt_cb<3> vss hvtnfet l=6e-08 w=8.58e-07 $X=21235 $Y=44959 $D=616
M775 vss 42 rt_cb<1> vss hvtnfet l=6e-08 w=8.58e-07 $X=21235 $Y=49947 $D=616
M776 rb_cb<1> 34 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=21495 $Y=328 $D=616
M777 rb_cb<3> 35 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=21495 $Y=5316 $D=616
M778 rb_mb<1> 36 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=21495 $Y=6788 $D=616
M779 rb_mb<3> 37 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=21495 $Y=11776 $D=616
M780 vss 20 rb_tm_preb_n vss hvtnfet l=6e-08 w=1.287e-06 $X=21495 $Y=13280 $D=616
M781 vss 21 rt_tm_preb_n vss hvtnfet l=6e-08 w=1.287e-06 $X=21495 $Y=20124 $D=616
M782 r_clk_dqb 8 vss vss hvtnfet l=6e-08 w=1.26e-06 $X=21495 $Y=22041 $D=616
M783 r_clk_dqb_n 9 vss vss hvtnfet l=6e-08 w=1.26e-06 $X=21495 $Y=29007 $D=616
M784 vss 10 r_lweb vss hvtnfet l=6e-08 w=1.287e-06 $X=21495 $Y=30897 $D=616
M785 r_sa_preb_n 51 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=21495 $Y=37027 $D=616
M786 rt_mb<3> 39 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=21495 $Y=38499 $D=616
M787 rt_mb<1> 40 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=21495 $Y=43487 $D=616
M788 rt_cb<3> 41 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=21495 $Y=44959 $D=616
M789 rt_cb<1> 42 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=21495 $Y=49947 $D=616
M790 vss 289 lb_ca<1> vss hvtnfet l=6e-08 w=8.58e-07 $X=22005 $Y=328 $D=616
M791 vss 290 lb_ca<3> vss hvtnfet l=6e-08 w=8.58e-07 $X=22005 $Y=5316 $D=616
M792 vss 291 lb_ma<1> vss hvtnfet l=6e-08 w=8.58e-07 $X=22005 $Y=6788 $D=616
M793 vss 292 lb_ma<3> vss hvtnfet l=6e-08 w=8.58e-07 $X=22005 $Y=11776 $D=616
M794 lb_tm_prea_n 285 vss vss hvtnfet l=6e-08 w=1.287e-06 $X=22005 $Y=13280 $D=616
M795 lt_tm_prea_n 286 vss vss hvtnfet l=6e-08 w=1.287e-06 $X=22005 $Y=20124 $D=616
M796 vss 287 l_clk_dqa vss hvtnfet l=6e-08 w=1.26e-06 $X=22005 $Y=22041 $D=616
M797 vss 288 l_clk_dqa_n vss hvtnfet l=6e-08 w=1.26e-06 $X=22005 $Y=29007 $D=616
M798 l_lwea 284 vss vss hvtnfet l=6e-08 w=1.287e-06 $X=22005 $Y=30897 $D=616
M799 vss 293 l_sa_prea_n vss hvtnfet l=6e-08 w=8.58e-07 $X=22005 $Y=37027 $D=616
M800 vss 294 lt_ma<3> vss hvtnfet l=6e-08 w=8.58e-07 $X=22005 $Y=38499 $D=616
M801 vss 295 lt_ma<1> vss hvtnfet l=6e-08 w=8.58e-07 $X=22005 $Y=43487 $D=616
M802 vss 296 lt_ca<3> vss hvtnfet l=6e-08 w=8.58e-07 $X=22005 $Y=44959 $D=616
M803 vss 297 lt_ca<1> vss hvtnfet l=6e-08 w=8.58e-07 $X=22005 $Y=49947 $D=616
M804 lb_ca<1> 289 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=22265 $Y=328 $D=616
M805 lb_ca<3> 290 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=22265 $Y=5316 $D=616
M806 lb_ma<1> 291 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=22265 $Y=6788 $D=616
M807 lb_ma<3> 292 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=22265 $Y=11776 $D=616
M808 vss 285 lb_tm_prea_n vss hvtnfet l=6e-08 w=1.287e-06 $X=22265 $Y=13280 $D=616
M809 vss 286 lt_tm_prea_n vss hvtnfet l=6e-08 w=1.287e-06 $X=22265 $Y=20124 $D=616
M810 l_clk_dqa 287 vss vss hvtnfet l=6e-08 w=1.26e-06 $X=22265 $Y=22041 $D=616
M811 l_clk_dqa_n 288 vss vss hvtnfet l=6e-08 w=1.26e-06 $X=22265 $Y=29007 $D=616
M812 vss 284 l_lwea vss hvtnfet l=6e-08 w=1.287e-06 $X=22265 $Y=30897 $D=616
M813 l_sa_prea_n 293 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=22265 $Y=37027 $D=616
M814 lt_ma<3> 294 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=22265 $Y=38499 $D=616
M815 lt_ma<1> 295 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=22265 $Y=43487 $D=616
M816 lt_ca<3> 296 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=22265 $Y=44959 $D=616
M817 lt_ca<1> 297 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=22265 $Y=49947 $D=616
M818 vss 289 lb_ca<1> vss hvtnfet l=6e-08 w=8.58e-07 $X=22525 $Y=328 $D=616
M819 vss 290 lb_ca<3> vss hvtnfet l=6e-08 w=8.58e-07 $X=22525 $Y=5316 $D=616
M820 vss 291 lb_ma<1> vss hvtnfet l=6e-08 w=8.58e-07 $X=22525 $Y=6788 $D=616
M821 vss 292 lb_ma<3> vss hvtnfet l=6e-08 w=8.58e-07 $X=22525 $Y=11776 $D=616
M822 vss 287 l_clk_dqa vss hvtnfet l=6e-08 w=1.26e-06 $X=22525 $Y=22041 $D=616
M823 vss 288 l_clk_dqa_n vss hvtnfet l=6e-08 w=1.26e-06 $X=22525 $Y=29007 $D=616
M824 vss 293 l_sa_prea_n vss hvtnfet l=6e-08 w=8.58e-07 $X=22525 $Y=37027 $D=616
M825 vss 294 lt_ma<3> vss hvtnfet l=6e-08 w=8.58e-07 $X=22525 $Y=38499 $D=616
M826 vss 295 lt_ma<1> vss hvtnfet l=6e-08 w=8.58e-07 $X=22525 $Y=43487 $D=616
M827 vss 296 lt_ca<3> vss hvtnfet l=6e-08 w=8.58e-07 $X=22525 $Y=44959 $D=616
M828 vss 297 lt_ca<1> vss hvtnfet l=6e-08 w=8.58e-07 $X=22525 $Y=49947 $D=616
M829 vss 298 284 vss hvtnfet l=6e-08 w=6e-07 $X=22775 $Y=30899 $D=616
M830 lb_ca<0> 299 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=22785 $Y=328 $D=616
M831 lb_ca<2> 300 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=22785 $Y=5316 $D=616
M832 lb_ma<0> 301 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=22785 $Y=6788 $D=616
M833 lb_ma<2> 302 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=22785 $Y=11776 $D=616
M834 l_saea_n 303 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=22785 $Y=37027 $D=616
M835 lt_ma<2> 304 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=22785 $Y=38499 $D=616
M836 lt_ma<0> 305 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=22785 $Y=43487 $D=616
M837 lt_ca<2> 306 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=22785 $Y=44959 $D=616
M838 lt_ca<0> 307 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=22785 $Y=49947 $D=616
M839 vss 299 lb_ca<0> vss hvtnfet l=6e-08 w=8.58e-07 $X=23045 $Y=328 $D=616
M840 vss 300 lb_ca<2> vss hvtnfet l=6e-08 w=8.58e-07 $X=23045 $Y=5316 $D=616
M841 vss 301 lb_ma<0> vss hvtnfet l=6e-08 w=8.58e-07 $X=23045 $Y=6788 $D=616
M842 vss 302 lb_ma<2> vss hvtnfet l=6e-08 w=8.58e-07 $X=23045 $Y=11776 $D=616
M843 vss 303 l_saea_n vss hvtnfet l=6e-08 w=8.58e-07 $X=23045 $Y=37027 $D=616
M844 vss 304 lt_ma<2> vss hvtnfet l=6e-08 w=8.58e-07 $X=23045 $Y=38499 $D=616
M845 vss 305 lt_ma<0> vss hvtnfet l=6e-08 w=8.58e-07 $X=23045 $Y=43487 $D=616
M846 vss 306 lt_ca<2> vss hvtnfet l=6e-08 w=8.58e-07 $X=23045 $Y=44959 $D=616
M847 vss 307 lt_ca<0> vss hvtnfet l=6e-08 w=8.58e-07 $X=23045 $Y=49947 $D=616
M848 1027 308 vss vss hvtnfet l=6e-08 w=1.8e-07 $X=23289 $Y=17143 $D=616
M849 308 312 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=23289 $Y=17812 $D=616
M850 309 313 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=23289 $Y=18983 $D=616
M851 1028 309 vss vss hvtnfet l=6e-08 w=1.8e-07 $X=23289 $Y=19609 $D=616
M852 1029 310 vss vss hvtnfet l=6e-08 w=1.8e-07 $X=23289 $Y=24063 $D=616
M853 310 314 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=23289 $Y=24732 $D=616
M854 311 315 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=23289 $Y=25903 $D=616
M855 1030 311 vss vss hvtnfet l=6e-08 w=1.8e-07 $X=23289 $Y=26529 $D=616
M856 lb_ca<0> 299 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=23305 $Y=328 $D=616
M857 lb_ca<2> 300 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=23305 $Y=5316 $D=616
M858 lb_ma<0> 301 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=23305 $Y=6788 $D=616
M859 lb_ma<2> 302 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=23305 $Y=11776 $D=616
M860 l_saea_n 303 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=23305 $Y=37027 $D=616
M861 lt_ma<2> 304 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=23305 $Y=38499 $D=616
M862 lt_ma<0> 305 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=23305 $Y=43487 $D=616
M863 lt_ca<2> 306 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=23305 $Y=44959 $D=616
M864 lt_ca<0> 307 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=23305 $Y=49947 $D=616
M865 312 317 1027 vss hvtnfet l=6e-08 w=1.8e-07 $X=23549 $Y=17143 $D=616
M866 vss 312 308 vss hvtnfet l=6e-08 w=1.37e-07 $X=23549 $Y=17812 $D=616
M867 vss 313 309 vss hvtnfet l=6e-08 w=1.37e-07 $X=23549 $Y=18983 $D=616
M868 313 317 1028 vss hvtnfet l=6e-08 w=1.8e-07 $X=23549 $Y=19609 $D=616
M869 314 317 1029 vss hvtnfet l=6e-08 w=1.8e-07 $X=23549 $Y=24063 $D=616
M870 vss 314 310 vss hvtnfet l=6e-08 w=1.37e-07 $X=23549 $Y=24732 $D=616
M871 vss 315 311 vss hvtnfet l=6e-08 w=1.37e-07 $X=23549 $Y=25903 $D=616
M872 315 317 1030 vss hvtnfet l=6e-08 w=1.8e-07 $X=23549 $Y=26529 $D=616
M873 vss 303 l_saea_n vss hvtnfet l=6e-08 w=8.58e-07 $X=23565 $Y=37027 $D=616
M874 l_saea_n 303 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=23825 $Y=37027 $D=616
M875 vss aa<0> 327 vss hvtnfet l=6e-08 w=2.74e-07 $X=23864 $Y=13476 $D=616
M876 vss 324 331 vss hvtnfet l=6e-08 w=2.1e-07 $X=24000 $Y=30918 $D=616
M877 vss 298 332 vss hvtnfet l=6e-08 w=2.1e-07 $X=24000 $Y=32688 $D=616
M878 1031 323 vss vss hvtnfet l=6e-08 w=8.23e-07 $X=24059 $Y=17143 $D=616
M879 1032 323 vss vss hvtnfet l=6e-08 w=8.23e-07 $X=24059 $Y=18966 $D=616
M880 1033 323 vss vss hvtnfet l=6e-08 w=8.23e-07 $X=24059 $Y=24063 $D=616
M881 1034 323 vss vss hvtnfet l=6e-08 w=8.23e-07 $X=24059 $Y=25886 $D=616
M882 b_pxca_n<7> 318 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=24060 $Y=336 $D=616
M883 318 319 vss vss hvtnfet l=6e-08 w=5e-07 $X=24060 $Y=6701 $D=616
M884 319 320 vss vss hvtnfet l=6e-08 w=3e-07 $X=24060 $Y=7831 $D=616
M885 321 320 vss vss hvtnfet l=6e-08 w=3e-07 $X=24060 $Y=43002 $D=616
M886 322 321 vss vss hvtnfet l=6e-08 w=5e-07 $X=24060 $Y=43932 $D=616
M887 t_pxca_n<7> 322 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=24060 $Y=49512 $D=616
M888 709 325 vss vss hvtnfet l=6e-08 w=4.8e-07 $X=24083 $Y=11276 $D=616
M889 710 clka vss vss hvtnfet l=6e-08 w=2.1e-07 $X=24260 $Y=30918 $D=616
M890 711 clka vss vss hvtnfet l=6e-08 w=2.1e-07 $X=24260 $Y=32688 $D=616
M891 vss 318 b_pxca_n<7> vss hvtnfet l=6e-08 w=1.285e-06 $X=24320 $Y=336 $D=616
M892 vss 319 318 vss hvtnfet l=6e-08 w=5e-07 $X=24320 $Y=6701 $D=616
M893 vss 320 319 vss hvtnfet l=6e-08 w=3e-07 $X=24320 $Y=7831 $D=616
M894 vss 320 321 vss hvtnfet l=6e-08 w=3e-07 $X=24320 $Y=43002 $D=616
M895 vss 321 322 vss hvtnfet l=6e-08 w=5e-07 $X=24320 $Y=43932 $D=616
M896 vss 322 t_pxca_n<7> vss hvtnfet l=6e-08 w=1.285e-06 $X=24320 $Y=49512 $D=616
M897 1035 328 1031 vss hvtnfet l=6e-08 w=5.49e-07 $X=24329 $Y=17143 $D=616
M898 1036 328 1032 vss hvtnfet l=6e-08 w=5.49e-07 $X=24329 $Y=19240 $D=616
M899 1037 329 1033 vss hvtnfet l=6e-08 w=5.49e-07 $X=24329 $Y=24063 $D=616
M900 1038 329 1034 vss hvtnfet l=6e-08 w=5.49e-07 $X=24329 $Y=26160 $D=616
M901 vss tm<8> 709 vss hvtnfet l=6e-08 w=4.8e-07 $X=24343 $Y=11276 $D=616
M902 334 327 vss vss hvtnfet l=6e-08 w=2.74e-07 $X=24374 $Y=13476 $D=616
M903 vss tm<5> 264 vss hvtnfet l=6e-08 w=2.74e-07 $X=24518 $Y=39358 $D=616
M904 324 331 710 vss hvtnfet l=6e-08 w=2.1e-07 $X=24520 $Y=30918 $D=616
M905 298 332 711 vss hvtnfet l=6e-08 w=2.1e-07 $X=24520 $Y=32688 $D=616
M906 312 334 1035 vss hvtnfet l=6e-08 w=5.49e-07 $X=24589 $Y=17143 $D=616
M907 313 327 1036 vss hvtnfet l=6e-08 w=5.49e-07 $X=24589 $Y=19240 $D=616
M908 314 334 1037 vss hvtnfet l=6e-08 w=5.49e-07 $X=24589 $Y=24063 $D=616
M909 315 327 1038 vss hvtnfet l=6e-08 w=5.49e-07 $X=24589 $Y=26160 $D=616
M910 714 340 324 vss hvtnfet l=6e-08 w=3.2e-07 $X=24780 $Y=30918 $D=616
M911 715 340 298 vss hvtnfet l=6e-08 w=3.2e-07 $X=24780 $Y=32578 $D=616
M912 b_pxca_n<6> 335 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=24830 $Y=336 $D=616
M913 335 336 vss vss hvtnfet l=6e-08 w=5e-07 $X=24830 $Y=6701 $D=616
M914 336 337 vss vss hvtnfet l=6e-08 w=3e-07 $X=24830 $Y=7831 $D=616
M915 338 337 vss vss hvtnfet l=6e-08 w=3e-07 $X=24830 $Y=43002 $D=616
M916 339 338 vss vss hvtnfet l=6e-08 w=5e-07 $X=24830 $Y=43932 $D=616
M917 t_pxca_n<6> 339 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=24830 $Y=49512 $D=616
M918 718 tm<8> vss vss hvtnfet l=6e-08 w=4.8e-07 $X=24853 $Y=11276 $D=616
M919 vss 264 376 vss hvtnfet l=6e-08 w=2e-07 $X=24874 $Y=37147 $D=616
M920 vss aa<1> 329 vss hvtnfet l=6e-08 w=2.74e-07 $X=24884 $Y=13476 $D=616
M921 vss aa<4> 714 vss hvtnfet l=6e-08 w=3.2e-07 $X=25040 $Y=30918 $D=616
M922 vss wena 715 vss hvtnfet l=6e-08 w=3.2e-07 $X=25040 $Y=32578 $D=616
M923 vss 335 b_pxca_n<6> vss hvtnfet l=6e-08 w=1.285e-06 $X=25090 $Y=336 $D=616
M924 vss 336 335 vss hvtnfet l=6e-08 w=5e-07 $X=25090 $Y=6701 $D=616
M925 vss 337 336 vss hvtnfet l=6e-08 w=3e-07 $X=25090 $Y=7831 $D=616
M926 vss 337 338 vss hvtnfet l=6e-08 w=3e-07 $X=25090 $Y=43002 $D=616
M927 vss 338 339 vss hvtnfet l=6e-08 w=5e-07 $X=25090 $Y=43932 $D=616
M928 vss 339 t_pxca_n<6> vss hvtnfet l=6e-08 w=1.285e-06 $X=25090 $Y=49512 $D=616
M929 vss tm<9> 718 vss hvtnfet l=6e-08 w=4.8e-07 $X=25113 $Y=11276 $D=616
M930 376 wena vss vss hvtnfet l=6e-08 w=2e-07 $X=25134 $Y=37147 $D=616
M931 328 329 vss vss hvtnfet l=6e-08 w=2.74e-07 $X=25394 $Y=13476 $D=616
M932 b_pxca_n<5> 345 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=25600 $Y=336 $D=616
M933 345 346 vss vss hvtnfet l=6e-08 w=5e-07 $X=25600 $Y=6701 $D=616
M934 346 347 vss vss hvtnfet l=6e-08 w=3e-07 $X=25600 $Y=7831 $D=616
M935 348 347 vss vss hvtnfet l=6e-08 w=3e-07 $X=25600 $Y=43002 $D=616
M936 349 348 vss vss hvtnfet l=6e-08 w=5e-07 $X=25600 $Y=43932 $D=616
M937 t_pxca_n<5> 349 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=25600 $Y=49512 $D=616
M938 1039 337 vss vss hvtnfet l=6e-08 w=1.8e-07 $X=25609 $Y=17143 $D=616
M939 1040 320 vss vss hvtnfet l=6e-08 w=1.8e-07 $X=25609 $Y=19609 $D=616
M940 1041 350 vss vss hvtnfet l=6e-08 w=1.8e-07 $X=25609 $Y=24063 $D=616
M941 1042 351 vss vss hvtnfet l=6e-08 w=1.8e-07 $X=25609 $Y=26529 $D=616
M942 721 tm<9> vss vss hvtnfet l=6e-08 w=4.8e-07 $X=25623 $Y=11276 $D=616
M943 337 352 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=25624 $Y=17812 $D=616
M944 320 353 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=25624 $Y=18983 $D=616
M945 350 354 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=25624 $Y=24732 $D=616
M946 351 355 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=25624 $Y=25903 $D=616
M947 vss clka 340 vss hvtnfet l=6e-08 w=4.5e-07 $X=25854 $Y=30668 $D=616
M948 vss 345 b_pxca_n<5> vss hvtnfet l=6e-08 w=1.285e-06 $X=25860 $Y=336 $D=616
M949 vss 346 345 vss hvtnfet l=6e-08 w=5e-07 $X=25860 $Y=6701 $D=616
M950 vss 347 346 vss hvtnfet l=6e-08 w=3e-07 $X=25860 $Y=7831 $D=616
M951 vss 347 348 vss hvtnfet l=6e-08 w=3e-07 $X=25860 $Y=43002 $D=616
M952 vss 348 349 vss hvtnfet l=6e-08 w=5e-07 $X=25860 $Y=43932 $D=616
M953 vss 349 t_pxca_n<5> vss hvtnfet l=6e-08 w=1.285e-06 $X=25860 $Y=49512 $D=616
M954 352 317 1039 vss hvtnfet l=6e-08 w=1.8e-07 $X=25869 $Y=17143 $D=616
M955 353 317 1040 vss hvtnfet l=6e-08 w=1.8e-07 $X=25869 $Y=19609 $D=616
M956 354 317 1041 vss hvtnfet l=6e-08 w=1.8e-07 $X=25869 $Y=24063 $D=616
M957 355 317 1042 vss hvtnfet l=6e-08 w=1.8e-07 $X=25869 $Y=26529 $D=616
M958 vss 366 721 vss hvtnfet l=6e-08 w=4.8e-07 $X=25883 $Y=11276 $D=616
M959 vss 352 337 vss hvtnfet l=6e-08 w=1.37e-07 $X=25884 $Y=17812 $D=616
M960 vss 353 320 vss hvtnfet l=6e-08 w=1.37e-07 $X=25884 $Y=18983 $D=616
M961 vss 354 350 vss hvtnfet l=6e-08 w=1.37e-07 $X=25884 $Y=24732 $D=616
M962 vss 355 351 vss hvtnfet l=6e-08 w=1.37e-07 $X=25884 $Y=25903 $D=616
M963 vss 356 363 vss hvtnfet l=6e-08 w=2.1e-07 $X=26138 $Y=37277 $D=616
M964 b_pxca_n<4> 357 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=26370 $Y=336 $D=616
M965 357 358 vss vss hvtnfet l=6e-08 w=5e-07 $X=26370 $Y=6701 $D=616
M966 358 359 vss vss hvtnfet l=6e-08 w=3e-07 $X=26370 $Y=7831 $D=616
M967 360 359 vss vss hvtnfet l=6e-08 w=3e-07 $X=26370 $Y=43002 $D=616
M968 361 360 vss vss hvtnfet l=6e-08 w=5e-07 $X=26370 $Y=43932 $D=616
M969 t_pxca_n<4> 361 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=26370 $Y=49512 $D=616
M970 729 123 733 vss hvtnfet l=6e-08 w=6e-07 $X=26374 $Y=30668 $D=616
M971 1043 323 vss vss hvtnfet l=6e-08 w=8.23e-07 $X=26379 $Y=17143 $D=616
M972 1044 323 vss vss hvtnfet l=6e-08 w=8.23e-07 $X=26379 $Y=18966 $D=616
M973 1045 323 vss vss hvtnfet l=6e-08 w=8.23e-07 $X=26379 $Y=24063 $D=616
M974 1046 323 vss vss hvtnfet l=6e-08 w=8.23e-07 $X=26379 $Y=25886 $D=616
M975 vss 366 727 vss hvtnfet l=6e-08 w=4.8e-07 $X=26393 $Y=11276 $D=616
M976 724 362 vss vss hvtnfet l=6e-08 w=2.1e-07 $X=26398 $Y=37277 $D=616
M977 vss 357 b_pxca_n<4> vss hvtnfet l=6e-08 w=1.285e-06 $X=26630 $Y=336 $D=616
M978 vss 358 357 vss hvtnfet l=6e-08 w=5e-07 $X=26630 $Y=6701 $D=616
M979 vss 359 358 vss hvtnfet l=6e-08 w=3e-07 $X=26630 $Y=7831 $D=616
M980 vss 359 360 vss hvtnfet l=6e-08 w=3e-07 $X=26630 $Y=43002 $D=616
M981 vss 360 361 vss hvtnfet l=6e-08 w=5e-07 $X=26630 $Y=43932 $D=616
M982 vss 361 t_pxca_n<4> vss hvtnfet l=6e-08 w=1.285e-06 $X=26630 $Y=49512 $D=616
M983 733 123 729 vss hvtnfet l=6e-08 w=6e-07 $X=26634 $Y=30668 $D=616
M984 1047 364 1043 vss hvtnfet l=6e-08 w=5.49e-07 $X=26649 $Y=17417 $D=616
M985 1048 364 1044 vss hvtnfet l=6e-08 w=5.49e-07 $X=26649 $Y=18966 $D=616
M986 1049 365 1045 vss hvtnfet l=6e-08 w=5.49e-07 $X=26649 $Y=24337 $D=616
M987 1050 365 1046 vss hvtnfet l=6e-08 w=5.49e-07 $X=26649 $Y=25886 $D=616
M988 727 325 vss vss hvtnfet l=6e-08 w=4.8e-07 $X=26653 $Y=11276 $D=616
M989 356 363 724 vss hvtnfet l=6e-08 w=2.1e-07 $X=26658 $Y=37277 $D=616
M990 vss tm<7> 726 vss hvtnfet l=6e-08 w=2.74e-07 $X=26820 $Y=39358 $D=616
M991 728 123 vss vss hvtnfet l=6e-08 w=3.2e-07 $X=26839 $Y=32578 $D=616
M992 vss 123 733 vss hvtnfet l=6e-08 w=6e-07 $X=26894 $Y=30668 $D=616
M993 1051 369 1047 vss hvtnfet l=6e-08 w=5.49e-07 $X=26909 $Y=17417 $D=616
M994 1052 369 1048 vss hvtnfet l=6e-08 w=5.49e-07 $X=26909 $Y=18966 $D=616
M995 1053 369 1049 vss hvtnfet l=6e-08 w=5.49e-07 $X=26909 $Y=24337 $D=616
M996 1054 369 1050 vss hvtnfet l=6e-08 w=5.49e-07 $X=26909 $Y=25886 $D=616
M997 730 368 356 vss hvtnfet l=6e-08 w=3.2e-07 $X=26918 $Y=37277 $D=616
M998 vss aa<10> 374 vss hvtnfet l=6e-08 w=2.74e-07 $X=26924 $Y=13476 $D=616
M999 379 123 728 vss hvtnfet l=6e-08 w=3.2e-07 $X=27099 $Y=32578 $D=616
M1000 b_pxca_n<3> 370 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=27140 $Y=336 $D=616
M1001 370 371 vss vss hvtnfet l=6e-08 w=5e-07 $X=27140 $Y=6701 $D=616
M1002 371 351 vss vss hvtnfet l=6e-08 w=3e-07 $X=27140 $Y=7831 $D=616
M1003 372 351 vss vss hvtnfet l=6e-08 w=3e-07 $X=27140 $Y=43002 $D=616
M1004 373 372 vss vss hvtnfet l=6e-08 w=5e-07 $X=27140 $Y=43932 $D=616
M1005 t_pxca_n<3> 373 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=27140 $Y=49512 $D=616
M1006 733 123 vss vss hvtnfet l=6e-08 w=6e-07 $X=27154 $Y=30668 $D=616
M1007 vss tm<9> 325 vss hvtnfet l=7e-08 w=3.2e-07 $X=27163 $Y=11276 $D=616
M1008 352 374 1051 vss hvtnfet l=6e-08 w=5.49e-07 $X=27169 $Y=17417 $D=616
M1009 353 375 1052 vss hvtnfet l=6e-08 w=5.49e-07 $X=27169 $Y=18966 $D=616
M1010 354 374 1053 vss hvtnfet l=6e-08 w=5.49e-07 $X=27169 $Y=24337 $D=616
M1011 355 375 1054 vss hvtnfet l=6e-08 w=5.49e-07 $X=27169 $Y=25886 $D=616
M1012 vss 376 730 vss hvtnfet l=6e-08 w=3.2e-07 $X=27178 $Y=37277 $D=616
M1013 375 374 vss vss hvtnfet l=6e-08 w=2.74e-07 $X=27184 $Y=13476 $D=616
M1014 734 377 379 vss hvtnfet l=6e-08 w=2.1e-07 $X=27359 $Y=32688 $D=616
M1015 vss 370 b_pxca_n<3> vss hvtnfet l=6e-08 w=1.285e-06 $X=27400 $Y=336 $D=616
M1016 vss 371 370 vss hvtnfet l=6e-08 w=5e-07 $X=27400 $Y=6701 $D=616
M1017 vss 351 371 vss hvtnfet l=6e-08 w=3e-07 $X=27400 $Y=7831 $D=616
M1018 vss 351 372 vss hvtnfet l=6e-08 w=3e-07 $X=27400 $Y=43002 $D=616
M1019 vss 372 373 vss hvtnfet l=6e-08 w=5e-07 $X=27400 $Y=43932 $D=616
M1020 vss 373 t_pxca_n<3> vss hvtnfet l=6e-08 w=1.285e-06 $X=27400 $Y=49512 $D=616
M1021 366 tm<8> vss vss hvtnfet l=7e-08 w=3.2e-07 $X=27433 $Y=11276 $D=616
M1022 vss 131 734 vss hvtnfet l=6e-08 w=2.1e-07 $X=27619 $Y=32688 $D=616
M1023 vss tm<1> 735 vss hvtnfet l=6e-08 w=2.74e-07 $X=27620 $Y=39358 $D=616
M1024 vss 380 369 vss hvtnfet l=6e-08 w=2.74e-07 $X=27784 $Y=13476 $D=616
M1025 737 362 386 vss hvtnfet l=6e-08 w=4e-07 $X=27858 $Y=37045 $D=616
M1026 377 379 vss vss hvtnfet l=6e-08 w=2.1e-07 $X=27879 $Y=32688 $D=616
M1027 b_pxca_n<2> 381 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=27910 $Y=336 $D=616
M1028 381 382 vss vss hvtnfet l=6e-08 w=5e-07 $X=27910 $Y=6701 $D=616
M1029 382 350 vss vss hvtnfet l=6e-08 w=3e-07 $X=27910 $Y=7831 $D=616
M1030 383 350 vss vss hvtnfet l=6e-08 w=3e-07 $X=27910 $Y=43002 $D=616
M1031 384 383 vss vss hvtnfet l=6e-08 w=5e-07 $X=27910 $Y=43932 $D=616
M1032 t_pxca_n<2> 384 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=27910 $Y=49512 $D=616
M1033 vss 323 317 vss hvtnfet l=6e-08 w=7e-07 $X=27924 $Y=30668 $D=616
M1034 380 aa<11> vss vss hvtnfet l=6e-08 w=2.74e-07 $X=28044 $Y=13476 $D=616
M1035 vss 356 737 vss hvtnfet l=6e-08 w=4e-07 $X=28118 $Y=37045 $D=616
M1036 vss 381 b_pxca_n<2> vss hvtnfet l=6e-08 w=1.285e-06 $X=28170 $Y=336 $D=616
M1037 vss 382 381 vss hvtnfet l=6e-08 w=5e-07 $X=28170 $Y=6701 $D=616
M1038 vss 350 382 vss hvtnfet l=6e-08 w=3e-07 $X=28170 $Y=7831 $D=616
M1039 vss 350 383 vss hvtnfet l=6e-08 w=3e-07 $X=28170 $Y=43002 $D=616
M1040 vss 383 384 vss hvtnfet l=6e-08 w=5e-07 $X=28170 $Y=43932 $D=616
M1041 vss 384 t_pxca_n<2> vss hvtnfet l=6e-08 w=1.285e-06 $X=28170 $Y=49512 $D=616
M1042 317 323 vss vss hvtnfet l=6e-08 w=7e-07 $X=28184 $Y=30668 $D=616
M1043 vss 392 541 vss hvtnfet l=6e-08 w=2e-07 $X=28514 $Y=11276 $D=616
M1044 vss 393 544 vss hvtnfet l=6e-08 w=2e-07 $X=28514 $Y=39657 $D=616
M1045 494 386 vss vss hvtnfet l=6e-08 w=2e-07 $X=28628 $Y=37045 $D=616
M1046 b_pxca_n<1> 387 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=28680 $Y=336 $D=616
M1047 387 388 vss vss hvtnfet l=6e-08 w=5e-07 $X=28680 $Y=6701 $D=616
M1048 388 389 vss vss hvtnfet l=6e-08 w=3e-07 $X=28680 $Y=7831 $D=616
M1049 390 389 vss vss hvtnfet l=6e-08 w=3e-07 $X=28680 $Y=43002 $D=616
M1050 391 390 vss vss hvtnfet l=6e-08 w=5e-07 $X=28680 $Y=43932 $D=616
M1051 t_pxca_n<1> 391 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=28680 $Y=49512 $D=616
M1052 742 123 vss vss hvtnfet l=6e-08 w=6e-07 $X=28704 $Y=30668 $D=616
M1053 vss 387 b_pxca_n<1> vss hvtnfet l=6e-08 w=1.285e-06 $X=28940 $Y=336 $D=616
M1054 vss 388 387 vss hvtnfet l=6e-08 w=5e-07 $X=28940 $Y=6701 $D=616
M1055 vss 389 388 vss hvtnfet l=6e-08 w=3e-07 $X=28940 $Y=7831 $D=616
M1056 vss 389 390 vss hvtnfet l=6e-08 w=3e-07 $X=28940 $Y=43002 $D=616
M1057 vss 390 391 vss hvtnfet l=6e-08 w=5e-07 $X=28940 $Y=43932 $D=616
M1058 vss 391 t_pxca_n<1> vss hvtnfet l=6e-08 w=1.285e-06 $X=28940 $Y=49512 $D=616
M1059 1055 374 407 vss hvtnfet l=6e-08 w=5.49e-07 $X=29009 $Y=17417 $D=616
M1060 1056 375 408 vss hvtnfet l=6e-08 w=5.49e-07 $X=29009 $Y=18966 $D=616
M1061 1057 374 409 vss hvtnfet l=6e-08 w=5.49e-07 $X=29009 $Y=24337 $D=616
M1062 1058 375 410 vss hvtnfet l=6e-08 w=5.49e-07 $X=29009 $Y=25886 $D=616
M1063 1059 308 vss vss hvtnfet l=6e-08 w=4.11e-07 $X=29024 $Y=11276 $D=616
M1064 1060 308 vss vss hvtnfet l=6e-08 w=4.11e-07 $X=29024 $Y=39446 $D=616
M1065 vss aa<12> 365 vss hvtnfet l=6e-08 w=2.74e-07 $X=29054 $Y=13476 $D=616
M1066 1061 380 1055 vss hvtnfet l=6e-08 w=5.49e-07 $X=29269 $Y=17417 $D=616
M1067 1062 380 1056 vss hvtnfet l=6e-08 w=5.49e-07 $X=29269 $Y=18966 $D=616
M1068 1063 380 1057 vss hvtnfet l=6e-08 w=5.49e-07 $X=29269 $Y=24337 $D=616
M1069 1064 380 1058 vss hvtnfet l=6e-08 w=5.49e-07 $X=29269 $Y=25886 $D=616
M1070 392 dwla<1> 1059 vss hvtnfet l=6e-08 w=4.11e-07 $X=29284 $Y=11276 $D=616
M1071 393 dwla<0> 1060 vss hvtnfet l=6e-08 w=4.11e-07 $X=29284 $Y=39446 $D=616
M1072 vss 395 403 vss hvtnfet l=6e-08 w=2e-07 $X=29298 $Y=32533 $D=616
M1073 b_pxca_n<0> 396 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=29450 $Y=336 $D=616
M1074 396 397 vss vss hvtnfet l=6e-08 w=5e-07 $X=29450 $Y=6701 $D=616
M1075 397 398 vss vss hvtnfet l=6e-08 w=3e-07 $X=29450 $Y=7831 $D=616
M1076 399 398 vss vss hvtnfet l=6e-08 w=3e-07 $X=29450 $Y=43002 $D=616
M1077 400 399 vss vss hvtnfet l=6e-08 w=5e-07 $X=29450 $Y=43932 $D=616
M1078 t_pxca_n<0> 400 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=29450 $Y=49512 $D=616
M1079 1065 364 1061 vss hvtnfet l=6e-08 w=5.49e-07 $X=29529 $Y=17417 $D=616
M1080 1066 364 1062 vss hvtnfet l=6e-08 w=5.49e-07 $X=29529 $Y=18966 $D=616
M1081 1067 365 1063 vss hvtnfet l=6e-08 w=5.49e-07 $X=29529 $Y=24337 $D=616
M1082 1068 365 1064 vss hvtnfet l=6e-08 w=5.49e-07 $X=29529 $Y=25886 $D=616
M1083 403 405 vss vss hvtnfet l=6e-08 w=2e-07 $X=29558 $Y=32533 $D=616
M1084 364 365 vss vss hvtnfet l=6e-08 w=2.74e-07 $X=29564 $Y=13476 $D=616
M1085 vss 404 395 vss hvtnfet l=6e-08 w=3.5e-07 $X=29621 $Y=30853 $D=616
M1086 vss 396 b_pxca_n<0> vss hvtnfet l=6e-08 w=1.285e-06 $X=29710 $Y=336 $D=616
M1087 vss 397 396 vss hvtnfet l=6e-08 w=5e-07 $X=29710 $Y=6701 $D=616
M1088 vss 398 397 vss hvtnfet l=6e-08 w=3e-07 $X=29710 $Y=7831 $D=616
M1089 vss 398 399 vss hvtnfet l=6e-08 w=3e-07 $X=29710 $Y=43002 $D=616
M1090 vss 399 400 vss hvtnfet l=6e-08 w=5e-07 $X=29710 $Y=43932 $D=616
M1091 vss 400 t_pxca_n<0> vss hvtnfet l=6e-08 w=1.285e-06 $X=29710 $Y=49512 $D=616
M1092 456 403 vss vss hvtnfet l=6e-08 w=6e-07 $X=29747 $Y=37037 $D=616
M1093 vss 323 1065 vss hvtnfet l=6e-08 w=8.23e-07 $X=29799 $Y=17143 $D=616
M1094 vss 323 1066 vss hvtnfet l=6e-08 w=8.23e-07 $X=29799 $Y=18966 $D=616
M1095 vss 323 1067 vss hvtnfet l=6e-08 w=8.23e-07 $X=29799 $Y=24063 $D=616
M1096 vss 323 1068 vss hvtnfet l=6e-08 w=8.23e-07 $X=29799 $Y=25886 $D=616
M1097 404 406 vss vss hvtnfet l=2.5e-07 w=3.5e-07 $X=29881 $Y=30853 $D=616
M1098 405 tm<7> vss vss hvtnfet l=6e-08 w=2e-07 $X=30068 $Y=32533 $D=616
M1099 dbl_pd_n<3> 131 vss vss hvtnfet l=6e-08 w=2.14e-07 $X=30204 $Y=13361 $D=616
M1100 b_pxba_n<7> 411 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=30220 $Y=336 $D=616
M1101 411 412 vss vss hvtnfet l=6e-08 w=5e-07 $X=30220 $Y=6701 $D=616
M1102 412 413 vss vss hvtnfet l=6e-08 w=3e-07 $X=30220 $Y=7831 $D=616
M1103 414 413 vss vss hvtnfet l=6e-08 w=3e-07 $X=30220 $Y=43002 $D=616
M1104 415 414 vss vss hvtnfet l=6e-08 w=5e-07 $X=30220 $Y=43932 $D=616
M1105 t_pxba_n<7> 415 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=30220 $Y=49512 $D=616
M1106 359 407 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=30294 $Y=17812 $D=616
M1107 347 408 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=30294 $Y=18983 $D=616
M1108 398 409 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=30294 $Y=24732 $D=616
M1109 389 410 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=30294 $Y=25903 $D=616
M1110 1069 317 407 vss hvtnfet l=6e-08 w=1.8e-07 $X=30309 $Y=17143 $D=616
M1111 1070 317 408 vss hvtnfet l=6e-08 w=1.8e-07 $X=30309 $Y=19609 $D=616
M1112 1071 317 409 vss hvtnfet l=6e-08 w=1.8e-07 $X=30309 $Y=24063 $D=616
M1113 1072 317 410 vss hvtnfet l=6e-08 w=1.8e-07 $X=30309 $Y=26529 $D=616
M1114 vss 131 dbl_pd_n<3> vss hvtnfet l=6e-08 w=2.14e-07 $X=30464 $Y=13361 $D=616
M1115 vss 411 b_pxba_n<7> vss hvtnfet l=6e-08 w=1.285e-06 $X=30480 $Y=336 $D=616
M1116 vss 412 411 vss hvtnfet l=6e-08 w=5e-07 $X=30480 $Y=6701 $D=616
M1117 vss 413 412 vss hvtnfet l=6e-08 w=3e-07 $X=30480 $Y=7831 $D=616
M1118 vss 413 414 vss hvtnfet l=6e-08 w=3e-07 $X=30480 $Y=43002 $D=616
M1119 vss 414 415 vss hvtnfet l=6e-08 w=5e-07 $X=30480 $Y=43932 $D=616
M1120 vss 415 t_pxba_n<7> vss hvtnfet l=6e-08 w=1.285e-06 $X=30480 $Y=49512 $D=616
M1121 456 416 vss vss hvtnfet l=6e-08 w=6e-07 $X=30527 $Y=37037 $D=616
M1122 vss 407 359 vss hvtnfet l=6e-08 w=1.37e-07 $X=30554 $Y=17812 $D=616
M1123 vss 408 347 vss hvtnfet l=6e-08 w=1.37e-07 $X=30554 $Y=18983 $D=616
M1124 vss 409 398 vss hvtnfet l=6e-08 w=1.37e-07 $X=30554 $Y=24732 $D=616
M1125 vss 410 389 vss hvtnfet l=6e-08 w=1.37e-07 $X=30554 $Y=25903 $D=616
M1126 vss 359 1069 vss hvtnfet l=6e-08 w=1.8e-07 $X=30569 $Y=17143 $D=616
M1127 vss 347 1070 vss hvtnfet l=6e-08 w=1.8e-07 $X=30569 $Y=19609 $D=616
M1128 vss 398 1071 vss hvtnfet l=6e-08 w=1.8e-07 $X=30569 $Y=24063 $D=616
M1129 vss 389 1072 vss hvtnfet l=6e-08 w=1.8e-07 $X=30569 $Y=26529 $D=616
M1130 1073 dwla<1> 426 vss hvtnfet l=6e-08 w=4.11e-07 $X=30584 $Y=11276 $D=616
M1131 1074 dwla<0> 427 vss hvtnfet l=6e-08 w=4.11e-07 $X=30584 $Y=39446 $D=616
M1132 vss 406 416 vss hvtnfet l=6e-08 w=2e-07 $X=30644 $Y=32533 $D=616
M1133 dbl_pd_n<3> 131 vss vss hvtnfet l=6e-08 w=2.14e-07 $X=30724 $Y=13361 $D=616
M1134 vss 417 406 vss hvtnfet l=6e-08 w=3.5e-07 $X=30741 $Y=30853 $D=616
M1135 vss 309 1073 vss hvtnfet l=6e-08 w=4.11e-07 $X=30844 $Y=11276 $D=616
M1136 vss 309 1074 vss hvtnfet l=6e-08 w=4.11e-07 $X=30844 $Y=39446 $D=616
M1137 416 423 vss vss hvtnfet l=6e-08 w=2e-07 $X=30904 $Y=32533 $D=616
M1138 b_pxba_n<6> 418 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=30990 $Y=336 $D=616
M1139 418 419 vss vss hvtnfet l=6e-08 w=5e-07 $X=30990 $Y=6701 $D=616
M1140 419 420 vss vss hvtnfet l=6e-08 w=3e-07 $X=30990 $Y=7831 $D=616
M1141 421 420 vss vss hvtnfet l=6e-08 w=3e-07 $X=30990 $Y=43002 $D=616
M1142 422 421 vss vss hvtnfet l=6e-08 w=5e-07 $X=30990 $Y=43932 $D=616
M1143 t_pxba_n<6> 422 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=30990 $Y=49512 $D=616
M1144 417 368 vss vss hvtnfet l=2.5e-07 w=3.5e-07 $X=31001 $Y=30853 $D=616
M1145 1075 420 vss vss hvtnfet l=6e-08 w=1.8e-07 $X=31079 $Y=17143 $D=616
M1146 1076 413 vss vss hvtnfet l=6e-08 w=1.8e-07 $X=31079 $Y=19609 $D=616
M1147 1077 424 vss vss hvtnfet l=6e-08 w=1.8e-07 $X=31079 $Y=24063 $D=616
M1148 1078 425 vss vss hvtnfet l=6e-08 w=1.8e-07 $X=31079 $Y=26529 $D=616
M1149 420 428 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=31094 $Y=17812 $D=616
M1150 413 429 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=31094 $Y=18983 $D=616
M1151 424 430 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=31094 $Y=24732 $D=616
M1152 425 431 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=31094 $Y=25903 $D=616
M1153 dbl_pd_n<1> tm<1> vss vss hvtnfet l=6e-08 w=2.14e-07 $X=31234 $Y=13361 $D=616
M1154 vss 418 b_pxba_n<6> vss hvtnfet l=6e-08 w=1.285e-06 $X=31250 $Y=336 $D=616
M1155 vss 419 418 vss hvtnfet l=6e-08 w=5e-07 $X=31250 $Y=6701 $D=616
M1156 vss 420 419 vss hvtnfet l=6e-08 w=3e-07 $X=31250 $Y=7831 $D=616
M1157 vss 420 421 vss hvtnfet l=6e-08 w=3e-07 $X=31250 $Y=43002 $D=616
M1158 vss 421 422 vss hvtnfet l=6e-08 w=5e-07 $X=31250 $Y=43932 $D=616
M1159 vss 422 t_pxba_n<6> vss hvtnfet l=6e-08 w=1.285e-06 $X=31250 $Y=49512 $D=616
M1160 456 362 vss vss hvtnfet l=6e-08 w=6e-07 $X=31307 $Y=37037 $D=616
M1161 428 317 1075 vss hvtnfet l=6e-08 w=1.8e-07 $X=31339 $Y=17143 $D=616
M1162 429 317 1076 vss hvtnfet l=6e-08 w=1.8e-07 $X=31339 $Y=19609 $D=616
M1163 430 317 1077 vss hvtnfet l=6e-08 w=1.8e-07 $X=31339 $Y=24063 $D=616
M1164 431 317 1078 vss hvtnfet l=6e-08 w=1.8e-07 $X=31339 $Y=26529 $D=616
M1165 556 426 vss vss hvtnfet l=6e-08 w=2e-07 $X=31354 $Y=11276 $D=616
M1166 vss 428 420 vss hvtnfet l=6e-08 w=1.37e-07 $X=31354 $Y=17812 $D=616
M1167 vss 429 413 vss hvtnfet l=6e-08 w=1.37e-07 $X=31354 $Y=18983 $D=616
M1168 vss 430 424 vss hvtnfet l=6e-08 w=1.37e-07 $X=31354 $Y=24732 $D=616
M1169 vss 431 425 vss hvtnfet l=6e-08 w=1.37e-07 $X=31354 $Y=25903 $D=616
M1170 558 427 vss vss hvtnfet l=6e-08 w=2e-07 $X=31354 $Y=39657 $D=616
M1171 vss 173 423 vss hvtnfet l=6e-08 w=2e-07 $X=31414 $Y=32533 $D=616
M1172 vss tm<1> dbl_pd_n<1> vss hvtnfet l=6e-08 w=2.14e-07 $X=31494 $Y=13361 $D=616
M1173 dbl_pd_n<1> tm<1> vss vss hvtnfet l=6e-08 w=2.14e-07 $X=31754 $Y=13361 $D=616
M1174 b_pxba_n<5> 432 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=31760 $Y=336 $D=616
M1175 432 433 vss vss hvtnfet l=6e-08 w=5e-07 $X=31760 $Y=6701 $D=616
M1176 433 434 vss vss hvtnfet l=6e-08 w=3e-07 $X=31760 $Y=7831 $D=616
M1177 435 434 vss vss hvtnfet l=6e-08 w=3e-07 $X=31760 $Y=43002 $D=616
M1178 436 435 vss vss hvtnfet l=6e-08 w=5e-07 $X=31760 $Y=43932 $D=616
M1179 t_pxba_n<5> 436 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=31760 $Y=49512 $D=616
M1180 vss 368 362 vss hvtnfet l=6e-08 w=2e-07 $X=31761 $Y=31098 $D=616
M1181 1079 323 vss vss hvtnfet l=6e-08 w=8.23e-07 $X=31849 $Y=17143 $D=616
M1182 1080 323 vss vss hvtnfet l=6e-08 w=8.23e-07 $X=31849 $Y=18966 $D=616
M1183 1081 323 vss vss hvtnfet l=6e-08 w=8.23e-07 $X=31849 $Y=24063 $D=616
M1184 1082 323 vss vss hvtnfet l=6e-08 w=8.23e-07 $X=31849 $Y=25886 $D=616
M1185 vss 437 540 vss hvtnfet l=6e-08 w=2e-07 $X=31864 $Y=11276 $D=616
M1186 vss 438 545 vss hvtnfet l=6e-08 w=2e-07 $X=31864 $Y=39657 $D=616
M1187 vss 432 b_pxba_n<5> vss hvtnfet l=6e-08 w=1.285e-06 $X=32020 $Y=336 $D=616
M1188 vss 433 432 vss hvtnfet l=6e-08 w=5e-07 $X=32020 $Y=6701 $D=616
M1189 vss 434 433 vss hvtnfet l=6e-08 w=3e-07 $X=32020 $Y=7831 $D=616
M1190 vss 434 435 vss hvtnfet l=6e-08 w=3e-07 $X=32020 $Y=43002 $D=616
M1191 vss 435 436 vss hvtnfet l=6e-08 w=5e-07 $X=32020 $Y=43932 $D=616
M1192 vss 436 t_pxba_n<5> vss hvtnfet l=6e-08 w=1.285e-06 $X=32020 $Y=49512 $D=616
M1193 1083 439 1079 vss hvtnfet l=6e-08 w=5.49e-07 $X=32119 $Y=17417 $D=616
M1194 1084 439 1080 vss hvtnfet l=6e-08 w=5.49e-07 $X=32119 $Y=18966 $D=616
M1195 1085 440 1081 vss hvtnfet l=6e-08 w=5.49e-07 $X=32119 $Y=24337 $D=616
M1196 1086 440 1082 vss hvtnfet l=6e-08 w=5.49e-07 $X=32119 $Y=25886 $D=616
M1197 dwla<1> 442 vss vss hvtnfet l=6e-08 w=3e-07 $X=32271 $Y=31098 $D=616
M1198 497 442 vss vss hvtnfet l=6e-08 w=3e-07 $X=32271 $Y=37457 $D=616
M1199 1087 310 vss vss hvtnfet l=6e-08 w=4.11e-07 $X=32374 $Y=11276 $D=616
M1200 1088 310 vss vss hvtnfet l=6e-08 w=4.11e-07 $X=32374 $Y=39446 $D=616
M1201 1089 443 1083 vss hvtnfet l=6e-08 w=5.49e-07 $X=32379 $Y=17417 $D=616
M1202 1090 443 1084 vss hvtnfet l=6e-08 w=5.49e-07 $X=32379 $Y=18966 $D=616
M1203 1091 443 1085 vss hvtnfet l=6e-08 w=5.49e-07 $X=32379 $Y=24337 $D=616
M1204 1092 443 1086 vss hvtnfet l=6e-08 w=5.49e-07 $X=32379 $Y=25886 $D=616
M1205 vss aa<7> 449 vss hvtnfet l=6e-08 w=2.74e-07 $X=32394 $Y=13476 $D=616
M1206 vss 324 442 vss hvtnfet l=6e-08 w=5e-07 $X=32394 $Y=32443 $D=616
M1207 b_pxba_n<4> 444 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=32530 $Y=336 $D=616
M1208 444 445 vss vss hvtnfet l=6e-08 w=5e-07 $X=32530 $Y=6701 $D=616
M1209 445 446 vss vss hvtnfet l=6e-08 w=3e-07 $X=32530 $Y=7831 $D=616
M1210 447 446 vss vss hvtnfet l=6e-08 w=3e-07 $X=32530 $Y=43002 $D=616
M1211 448 447 vss vss hvtnfet l=6e-08 w=5e-07 $X=32530 $Y=43932 $D=616
M1212 t_pxba_n<4> 448 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=32530 $Y=49512 $D=616
M1213 vss 442 dwla<1> vss hvtnfet l=6e-08 w=3e-07 $X=32531 $Y=31098 $D=616
M1214 vss 442 497 vss hvtnfet l=6e-08 w=3e-07 $X=32531 $Y=37457 $D=616
M1215 437 dwla<1> 1087 vss hvtnfet l=6e-08 w=4.11e-07 $X=32634 $Y=11276 $D=616
M1216 438 dwla<0> 1088 vss hvtnfet l=6e-08 w=4.11e-07 $X=32634 $Y=39446 $D=616
M1217 428 449 1089 vss hvtnfet l=6e-08 w=5.49e-07 $X=32639 $Y=17417 $D=616
M1218 429 450 1090 vss hvtnfet l=6e-08 w=5.49e-07 $X=32639 $Y=18966 $D=616
M1219 430 449 1091 vss hvtnfet l=6e-08 w=5.49e-07 $X=32639 $Y=24337 $D=616
M1220 431 450 1092 vss hvtnfet l=6e-08 w=5.49e-07 $X=32639 $Y=25886 $D=616
M1221 450 449 vss vss hvtnfet l=6e-08 w=2.74e-07 $X=32654 $Y=13476 $D=616
M1222 vss 444 b_pxba_n<4> vss hvtnfet l=6e-08 w=1.285e-06 $X=32790 $Y=336 $D=616
M1223 vss 445 444 vss hvtnfet l=6e-08 w=5e-07 $X=32790 $Y=6701 $D=616
M1224 vss 446 445 vss hvtnfet l=6e-08 w=3e-07 $X=32790 $Y=7831 $D=616
M1225 vss 446 447 vss hvtnfet l=6e-08 w=3e-07 $X=32790 $Y=43002 $D=616
M1226 vss 447 448 vss hvtnfet l=6e-08 w=5e-07 $X=32790 $Y=43932 $D=616
M1227 vss 448 t_pxba_n<4> vss hvtnfet l=6e-08 w=1.285e-06 $X=32790 $Y=49512 $D=616
M1228 dwla<1> 368 vss vss hvtnfet l=6e-08 w=3e-07 $X=33041 $Y=31098 $D=616
M1229 497 456 vss vss hvtnfet l=6e-08 w=3e-07 $X=33041 $Y=37457 $D=616
M1230 465 442 vss vss hvtnfet l=6e-08 w=4e-07 $X=33094 $Y=32543 $D=616
M1231 1093 dwla<1> 458 vss hvtnfet l=6e-08 w=4.11e-07 $X=33144 $Y=11276 $D=616
M1232 1094 dwla<0> 459 vss hvtnfet l=6e-08 w=4.11e-07 $X=33144 $Y=39446 $D=616
M1233 vss 455 443 vss hvtnfet l=6e-08 w=2.74e-07 $X=33254 $Y=13476 $D=616
M1234 b_pxba_n<3> 451 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=33300 $Y=336 $D=616
M1235 451 452 vss vss hvtnfet l=6e-08 w=5e-07 $X=33300 $Y=6701 $D=616
M1236 452 425 vss vss hvtnfet l=6e-08 w=3e-07 $X=33300 $Y=7831 $D=616
M1237 453 425 vss vss hvtnfet l=6e-08 w=3e-07 $X=33300 $Y=43002 $D=616
M1238 454 453 vss vss hvtnfet l=6e-08 w=5e-07 $X=33300 $Y=43932 $D=616
M1239 t_pxba_n<3> 454 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=33300 $Y=49512 $D=616
M1240 vss 368 dwla<1> vss hvtnfet l=6e-08 w=3e-07 $X=33301 $Y=31098 $D=616
M1241 vss 456 497 vss hvtnfet l=6e-08 w=3e-07 $X=33301 $Y=37457 $D=616
M1242 vss 311 1093 vss hvtnfet l=6e-08 w=4.11e-07 $X=33404 $Y=11276 $D=616
M1243 vss 311 1094 vss hvtnfet l=6e-08 w=4.11e-07 $X=33404 $Y=39446 $D=616
M1244 455 aa<8> vss vss hvtnfet l=6e-08 w=2.74e-07 $X=33514 $Y=13476 $D=616
M1245 vss 451 b_pxba_n<3> vss hvtnfet l=6e-08 w=1.285e-06 $X=33560 $Y=336 $D=616
M1246 vss 452 451 vss hvtnfet l=6e-08 w=5e-07 $X=33560 $Y=6701 $D=616
M1247 vss 425 452 vss hvtnfet l=6e-08 w=3e-07 $X=33560 $Y=7831 $D=616
M1248 vss 425 453 vss hvtnfet l=6e-08 w=3e-07 $X=33560 $Y=43002 $D=616
M1249 vss 453 454 vss hvtnfet l=6e-08 w=5e-07 $X=33560 $Y=43932 $D=616
M1250 vss 454 t_pxba_n<3> vss hvtnfet l=6e-08 w=1.285e-06 $X=33560 $Y=49512 $D=616
M1251 dwla<0> 368 vss vss hvtnfet l=6e-08 w=3e-07 $X=33811 $Y=31098 $D=616
M1252 498 456 vss vss hvtnfet l=6e-08 w=3e-07 $X=33811 $Y=37457 $D=616
M1253 555 458 vss vss hvtnfet l=6e-08 w=2e-07 $X=33914 $Y=11276 $D=616
M1254 559 459 vss vss hvtnfet l=6e-08 w=2e-07 $X=33914 $Y=39657 $D=616
M1255 b_pxba_n<2> 460 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=34070 $Y=336 $D=616
M1256 460 461 vss vss hvtnfet l=6e-08 w=5e-07 $X=34070 $Y=6701 $D=616
M1257 461 424 vss vss hvtnfet l=6e-08 w=3e-07 $X=34070 $Y=7831 $D=616
M1258 462 424 vss vss hvtnfet l=6e-08 w=3e-07 $X=34070 $Y=43002 $D=616
M1259 463 462 vss vss hvtnfet l=6e-08 w=5e-07 $X=34070 $Y=43932 $D=616
M1260 t_pxba_n<2> 463 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=34070 $Y=49512 $D=616
M1261 vss 368 dwla<0> vss hvtnfet l=6e-08 w=3e-07 $X=34071 $Y=31098 $D=616
M1262 vss 456 498 vss hvtnfet l=6e-08 w=3e-07 $X=34071 $Y=37457 $D=616
M1263 vss 460 b_pxba_n<2> vss hvtnfet l=6e-08 w=1.285e-06 $X=34330 $Y=336 $D=616
M1264 vss 461 460 vss hvtnfet l=6e-08 w=5e-07 $X=34330 $Y=6701 $D=616
M1265 vss 424 461 vss hvtnfet l=6e-08 w=3e-07 $X=34330 $Y=7831 $D=616
M1266 vss 424 462 vss hvtnfet l=6e-08 w=3e-07 $X=34330 $Y=43002 $D=616
M1267 vss 462 463 vss hvtnfet l=6e-08 w=5e-07 $X=34330 $Y=43932 $D=616
M1268 vss 463 t_pxba_n<2> vss hvtnfet l=6e-08 w=1.285e-06 $X=34330 $Y=49512 $D=616
M1269 1095 449 479 vss hvtnfet l=6e-08 w=5.49e-07 $X=34479 $Y=17417 $D=616
M1270 1096 450 480 vss hvtnfet l=6e-08 w=5.49e-07 $X=34479 $Y=18966 $D=616
M1271 1097 449 481 vss hvtnfet l=6e-08 w=5.49e-07 $X=34479 $Y=24337 $D=616
M1272 1098 450 482 vss hvtnfet l=6e-08 w=5.49e-07 $X=34479 $Y=25886 $D=616
M1273 vss aa<9> 440 vss hvtnfet l=6e-08 w=2.74e-07 $X=34524 $Y=13476 $D=616
M1274 dwla<0> 465 vss vss hvtnfet l=6e-08 w=3e-07 $X=34581 $Y=31098 $D=616
M1275 498 465 vss vss hvtnfet l=6e-08 w=3e-07 $X=34581 $Y=37457 $D=616
M1276 1099 vdd vss vss hvtnfet l=6e-08 w=6.4e-07 $X=34621 $Y=32508 $D=616
M1277 123 131 vss vss hvtnfet l=6e-08 w=2e-07 $X=34646 $Y=11546 $D=616
M1278 1100 455 1095 vss hvtnfet l=6e-08 w=5.49e-07 $X=34739 $Y=17417 $D=616
M1279 1101 455 1096 vss hvtnfet l=6e-08 w=5.49e-07 $X=34739 $Y=18966 $D=616
M1280 1102 455 1097 vss hvtnfet l=6e-08 w=5.49e-07 $X=34739 $Y=24337 $D=616
M1281 1103 455 1098 vss hvtnfet l=6e-08 w=5.49e-07 $X=34739 $Y=25886 $D=616
M1282 b_pxba_n<1> 466 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=34840 $Y=336 $D=616
M1283 466 467 vss vss hvtnfet l=6e-08 w=5e-07 $X=34840 $Y=6701 $D=616
M1284 467 468 vss vss hvtnfet l=6e-08 w=3e-07 $X=34840 $Y=7831 $D=616
M1285 469 468 vss vss hvtnfet l=6e-08 w=3e-07 $X=34840 $Y=43002 $D=616
M1286 470 469 vss vss hvtnfet l=6e-08 w=5e-07 $X=34840 $Y=43932 $D=616
M1287 t_pxba_n<1> 470 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=34840 $Y=49512 $D=616
M1288 vss 465 dwla<0> vss hvtnfet l=6e-08 w=3e-07 $X=34841 $Y=31098 $D=616
M1289 vss 465 498 vss hvtnfet l=6e-08 w=3e-07 $X=34841 $Y=37457 $D=616
M1290 535 471 1099 vss hvtnfet l=6e-08 w=6.4e-07 $X=34881 $Y=32508 $D=616
M1291 vss 123 123 vss hvtnfet l=6e-08 w=2e-07 $X=34906 $Y=11546 $D=616
M1292 1104 439 1100 vss hvtnfet l=6e-08 w=5.49e-07 $X=34999 $Y=17417 $D=616
M1293 1105 439 1101 vss hvtnfet l=6e-08 w=5.49e-07 $X=34999 $Y=18966 $D=616
M1294 1106 440 1102 vss hvtnfet l=6e-08 w=5.49e-07 $X=34999 $Y=24337 $D=616
M1295 1107 440 1103 vss hvtnfet l=6e-08 w=5.49e-07 $X=34999 $Y=25886 $D=616
M1296 439 440 vss vss hvtnfet l=6e-08 w=2.74e-07 $X=35034 $Y=13476 $D=616
M1297 vss 466 b_pxba_n<1> vss hvtnfet l=6e-08 w=1.285e-06 $X=35100 $Y=336 $D=616
M1298 vss 467 466 vss hvtnfet l=6e-08 w=5e-07 $X=35100 $Y=6701 $D=616
M1299 vss 468 467 vss hvtnfet l=6e-08 w=3e-07 $X=35100 $Y=7831 $D=616
M1300 vss 468 469 vss hvtnfet l=6e-08 w=3e-07 $X=35100 $Y=43002 $D=616
M1301 vss 469 470 vss hvtnfet l=6e-08 w=5e-07 $X=35100 $Y=43932 $D=616
M1302 vss 470 t_pxba_n<1> vss hvtnfet l=6e-08 w=1.285e-06 $X=35100 $Y=49512 $D=616
M1303 vss 323 1104 vss hvtnfet l=6e-08 w=8.23e-07 $X=35269 $Y=17143 $D=616
M1304 vss 323 1105 vss hvtnfet l=6e-08 w=8.23e-07 $X=35269 $Y=18966 $D=616
M1305 vss 323 1106 vss hvtnfet l=6e-08 w=8.23e-07 $X=35269 $Y=24063 $D=616
M1306 vss 323 1107 vss hvtnfet l=6e-08 w=8.23e-07 $X=35269 $Y=25886 $D=616
M1307 vss 473 484 vss hvtnfet l=6e-08 w=3e-07 $X=35351 $Y=37257 $D=616
M1308 vss 472 471 vss hvtnfet l=6e-08 w=3.5e-07 $X=35446 $Y=32613 $D=616
M1309 b_pxba_n<0> 474 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=35610 $Y=336 $D=616
M1310 474 475 vss vss hvtnfet l=6e-08 w=5e-07 $X=35610 $Y=6701 $D=616
M1311 475 476 vss vss hvtnfet l=6e-08 w=3e-07 $X=35610 $Y=7831 $D=616
M1312 477 476 vss vss hvtnfet l=6e-08 w=3e-07 $X=35610 $Y=43002 $D=616
M1313 478 477 vss vss hvtnfet l=6e-08 w=5e-07 $X=35610 $Y=43932 $D=616
M1314 t_pxba_n<0> 478 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=35610 $Y=49512 $D=616
M1315 472 483 vss vss hvtnfet l=2.5e-07 w=3.5e-07 $X=35706 $Y=32613 $D=616
M1316 446 479 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=35764 $Y=17812 $D=616
M1317 434 480 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=35764 $Y=18983 $D=616
M1318 476 481 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=35764 $Y=24732 $D=616
M1319 468 482 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=35764 $Y=25903 $D=616
M1320 1108 317 479 vss hvtnfet l=6e-08 w=1.8e-07 $X=35779 $Y=17143 $D=616
M1321 1109 317 480 vss hvtnfet l=6e-08 w=1.8e-07 $X=35779 $Y=19609 $D=616
M1322 1110 317 481 vss hvtnfet l=6e-08 w=1.8e-07 $X=35779 $Y=24063 $D=616
M1323 1111 317 482 vss hvtnfet l=6e-08 w=1.8e-07 $X=35779 $Y=26529 $D=616
M1324 473 484 vss vss hvtnfet l=1.2e-07 w=1.5e-07 $X=35861 $Y=37297 $D=616
M1325 vss 474 b_pxba_n<0> vss hvtnfet l=6e-08 w=1.285e-06 $X=35870 $Y=336 $D=616
M1326 vss 475 474 vss hvtnfet l=6e-08 w=5e-07 $X=35870 $Y=6701 $D=616
M1327 vss 476 475 vss hvtnfet l=6e-08 w=3e-07 $X=35870 $Y=7831 $D=616
M1328 vss 476 477 vss hvtnfet l=6e-08 w=3e-07 $X=35870 $Y=43002 $D=616
M1329 vss 477 478 vss hvtnfet l=6e-08 w=5e-07 $X=35870 $Y=43932 $D=616
M1330 vss 478 t_pxba_n<0> vss hvtnfet l=6e-08 w=1.285e-06 $X=35870 $Y=49512 $D=616
M1331 773 495 vss vss hvtnfet l=6e-08 w=8e-07 $X=35945 $Y=30668 $D=616
M1332 vss 479 446 vss hvtnfet l=6e-08 w=1.37e-07 $X=36024 $Y=17812 $D=616
M1333 vss 480 434 vss hvtnfet l=6e-08 w=1.37e-07 $X=36024 $Y=18983 $D=616
M1334 vss 481 476 vss hvtnfet l=6e-08 w=1.37e-07 $X=36024 $Y=24732 $D=616
M1335 vss 482 468 vss hvtnfet l=6e-08 w=1.37e-07 $X=36024 $Y=25903 $D=616
M1336 vss 446 1108 vss hvtnfet l=6e-08 w=1.8e-07 $X=36039 $Y=17143 $D=616
M1337 vss 434 1109 vss hvtnfet l=6e-08 w=1.8e-07 $X=36039 $Y=19609 $D=616
M1338 vss 476 1110 vss hvtnfet l=6e-08 w=1.8e-07 $X=36039 $Y=24063 $D=616
M1339 vss 468 1111 vss hvtnfet l=6e-08 w=1.8e-07 $X=36039 $Y=26529 $D=616
M1340 vss 495 773 vss hvtnfet l=6e-08 w=8e-07 $X=36205 $Y=30668 $D=616
M1341 vss 491 509 vss hvtnfet l=6e-08 w=2.74e-07 $X=36254 $Y=13476 $D=616
M1342 b_pxaa<3> 485 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=36380 $Y=336 $D=616
M1343 485 486 vss vss hvtnfet l=6e-08 w=5e-07 $X=36380 $Y=6701 $D=616
M1344 486 487 vss vss hvtnfet l=6e-08 w=3e-07 $X=36380 $Y=7831 $D=616
M1345 1112 492 vss vss hvtnfet l=6e-08 w=4.11e-07 $X=36380 $Y=11276 $D=616
M1346 1113 492 vss vss hvtnfet l=6e-08 w=4.11e-07 $X=36380 $Y=39446 $D=616
M1347 489 488 vss vss hvtnfet l=6e-08 w=3e-07 $X=36380 $Y=43002 $D=616
M1348 490 489 vss vss hvtnfet l=6e-08 w=5e-07 $X=36380 $Y=43932 $D=616
M1349 t_pxaa<3> 490 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=36380 $Y=49512 $D=616
M1350 vss 494 473 vss hvtnfet l=6e-08 w=3.2e-07 $X=36431 $Y=37292 $D=616
M1351 vss 496 483 vss hvtnfet l=6e-08 w=3.2e-07 $X=36466 $Y=32828 $D=616
M1352 vss 485 b_pxaa<3> vss hvtnfet l=6e-08 w=1.285e-06 $X=36640 $Y=336 $D=616
M1353 vss 486 485 vss hvtnfet l=6e-08 w=5e-07 $X=36640 $Y=6701 $D=616
M1354 vss 487 486 vss hvtnfet l=6e-08 w=3e-07 $X=36640 $Y=7831 $D=616
M1355 487 497 1112 vss hvtnfet l=6e-08 w=4.11e-07 $X=36640 $Y=11276 $D=616
M1356 488 498 1113 vss hvtnfet l=6e-08 w=4.11e-07 $X=36640 $Y=39446 $D=616
M1357 vss 488 489 vss hvtnfet l=6e-08 w=3e-07 $X=36640 $Y=43002 $D=616
M1358 vss 489 490 vss hvtnfet l=6e-08 w=5e-07 $X=36640 $Y=43932 $D=616
M1359 vss 490 t_pxaa<3> vss hvtnfet l=6e-08 w=1.285e-06 $X=36640 $Y=49512 $D=616
M1360 368 clka 773 vss hvtnfet l=6e-08 w=8e-07 $X=36715 $Y=30668 $D=616
M1361 491 aa<6> vss vss hvtnfet l=6e-08 w=2.74e-07 $X=36764 $Y=13476 $D=616
M1362 773 clka 368 vss hvtnfet l=6e-08 w=8e-07 $X=36975 $Y=30668 $D=616
M1363 vss 473 496 vss hvtnfet l=6e-08 w=3.2e-07 $X=36976 $Y=32828 $D=616
M1364 1114 501 519 vss hvtnfet l=6e-08 w=5.49e-07 $X=37059 $Y=17143 $D=616
M1365 1115 502 520 vss hvtnfet l=6e-08 w=5.49e-07 $X=37059 $Y=19240 $D=616
M1366 1116 501 521 vss hvtnfet l=6e-08 w=5.49e-07 $X=37059 $Y=24063 $D=616
M1367 1117 502 522 vss hvtnfet l=6e-08 w=5.49e-07 $X=37059 $Y=26160 $D=616
M1368 b_pxaa<2> 503 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=37150 $Y=336 $D=616
M1369 503 504 vss vss hvtnfet l=6e-08 w=5e-07 $X=37150 $Y=6701 $D=616
M1370 504 505 vss vss hvtnfet l=6e-08 w=3e-07 $X=37150 $Y=7831 $D=616
M1371 1118 497 505 vss hvtnfet l=6e-08 w=4.11e-07 $X=37150 $Y=11276 $D=616
M1372 1119 498 506 vss hvtnfet l=6e-08 w=4.11e-07 $X=37150 $Y=39446 $D=616
M1373 507 506 vss vss hvtnfet l=6e-08 w=3e-07 $X=37150 $Y=43002 $D=616
M1374 508 507 vss vss hvtnfet l=6e-08 w=5e-07 $X=37150 $Y=43932 $D=616
M1375 t_pxaa<2> 508 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=37150 $Y=49512 $D=616
M1376 vss ddqa_n 493 vss hvtnfet l=6e-08 w=2.4e-07 $X=37161 $Y=37292 $D=616
M1377 vss 502 501 vss hvtnfet l=6e-08 w=2.74e-07 $X=37274 $Y=13476 $D=616
M1378 1120 509 1114 vss hvtnfet l=6e-08 w=5.49e-07 $X=37319 $Y=17143 $D=616
M1379 1121 509 1115 vss hvtnfet l=6e-08 w=5.49e-07 $X=37319 $Y=19240 $D=616
M1380 1122 491 1116 vss hvtnfet l=6e-08 w=5.49e-07 $X=37319 $Y=24063 $D=616
M1381 1123 491 1117 vss hvtnfet l=6e-08 w=5.49e-07 $X=37319 $Y=26160 $D=616
M1382 vss 503 b_pxaa<2> vss hvtnfet l=6e-08 w=1.285e-06 $X=37410 $Y=336 $D=616
M1383 vss 504 503 vss hvtnfet l=6e-08 w=5e-07 $X=37410 $Y=6701 $D=616
M1384 vss 505 504 vss hvtnfet l=6e-08 w=3e-07 $X=37410 $Y=7831 $D=616
M1385 vss 510 1118 vss hvtnfet l=6e-08 w=4.11e-07 $X=37410 $Y=11276 $D=616
M1386 vss 510 1119 vss hvtnfet l=6e-08 w=4.11e-07 $X=37410 $Y=39446 $D=616
M1387 vss 506 507 vss hvtnfet l=6e-08 w=3e-07 $X=37410 $Y=43002 $D=616
M1388 vss 507 508 vss hvtnfet l=6e-08 w=5e-07 $X=37410 $Y=43932 $D=616
M1389 vss 508 t_pxaa<2> vss hvtnfet l=6e-08 w=1.285e-06 $X=37410 $Y=49512 $D=616
M1390 493 ddqa vss vss hvtnfet l=6e-08 w=2.4e-07 $X=37421 $Y=37292 $D=616
M1391 vss clka 524 vss hvtnfet l=6e-08 w=6e-07 $X=37485 $Y=30668 $D=616
M1392 vss 323 1120 vss hvtnfet l=6e-08 w=8.23e-07 $X=37589 $Y=17143 $D=616
M1393 vss 323 1121 vss hvtnfet l=6e-08 w=8.23e-07 $X=37589 $Y=18966 $D=616
M1394 vss 323 1122 vss hvtnfet l=6e-08 w=8.23e-07 $X=37589 $Y=24063 $D=616
M1395 vss 323 1123 vss hvtnfet l=6e-08 w=8.23e-07 $X=37589 $Y=25886 $D=616
M1396 1124 496 557 vss hvtnfet l=6e-08 w=6.4e-07 $X=37661 $Y=32508 $D=616
M1397 502 aa<5> vss vss hvtnfet l=6e-08 w=2.74e-07 $X=37784 $Y=13476 $D=616
M1398 b_pxaa<1> 512 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=37920 $Y=336 $D=616
M1399 512 513 vss vss hvtnfet l=6e-08 w=5e-07 $X=37920 $Y=6701 $D=616
M1400 513 514 vss vss hvtnfet l=6e-08 w=3e-07 $X=37920 $Y=7831 $D=616
M1401 1125 523 vss vss hvtnfet l=6e-08 w=4.11e-07 $X=37920 $Y=11276 $D=616
M1402 1126 523 vss vss hvtnfet l=6e-08 w=4.11e-07 $X=37920 $Y=39446 $D=616
M1403 516 515 vss vss hvtnfet l=6e-08 w=3e-07 $X=37920 $Y=43002 $D=616
M1404 517 516 vss vss hvtnfet l=6e-08 w=5e-07 $X=37920 $Y=43932 $D=616
M1405 t_pxaa<1> 517 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=37920 $Y=49512 $D=616
M1406 vss 386 1124 vss hvtnfet l=6e-08 w=6.4e-07 $X=37921 $Y=32508 $D=616
M1407 1127 317 519 vss hvtnfet l=6e-08 w=1.8e-07 $X=38099 $Y=17143 $D=616
M1408 492 519 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=38099 $Y=17812 $D=616
M1409 510 520 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=38099 $Y=18983 $D=616
M1410 1128 317 520 vss hvtnfet l=6e-08 w=1.8e-07 $X=38099 $Y=19609 $D=616
M1411 1129 317 521 vss hvtnfet l=6e-08 w=1.8e-07 $X=38099 $Y=24063 $D=616
M1412 523 521 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=38099 $Y=24732 $D=616
M1413 525 522 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=38099 $Y=25903 $D=616
M1414 1130 317 522 vss hvtnfet l=6e-08 w=1.8e-07 $X=38099 $Y=26529 $D=616
M1415 vss 493 526 vss hvtnfet l=1.4e-07 w=3.2e-07 $X=38141 $Y=37127 $D=616
M1416 vss 512 b_pxaa<1> vss hvtnfet l=6e-08 w=1.285e-06 $X=38180 $Y=336 $D=616
M1417 vss 513 512 vss hvtnfet l=6e-08 w=5e-07 $X=38180 $Y=6701 $D=616
M1418 vss 514 513 vss hvtnfet l=6e-08 w=3e-07 $X=38180 $Y=7831 $D=616
M1419 514 497 1125 vss hvtnfet l=6e-08 w=4.11e-07 $X=38180 $Y=11276 $D=616
M1420 515 498 1126 vss hvtnfet l=6e-08 w=4.11e-07 $X=38180 $Y=39446 $D=616
M1421 vss 515 516 vss hvtnfet l=6e-08 w=3e-07 $X=38180 $Y=43002 $D=616
M1422 vss 516 517 vss hvtnfet l=6e-08 w=5e-07 $X=38180 $Y=43932 $D=616
M1423 vss 517 t_pxaa<1> vss hvtnfet l=6e-08 w=1.285e-06 $X=38180 $Y=49512 $D=616
M1424 vss 524 534 vss hvtnfet l=6e-08 w=5.49e-07 $X=38255 $Y=30668 $D=616
M1425 vss 492 1127 vss hvtnfet l=6e-08 w=1.8e-07 $X=38359 $Y=17143 $D=616
M1426 vss 519 492 vss hvtnfet l=6e-08 w=1.37e-07 $X=38359 $Y=17812 $D=616
M1427 vss 520 510 vss hvtnfet l=6e-08 w=1.37e-07 $X=38359 $Y=18983 $D=616
M1428 vss 510 1128 vss hvtnfet l=6e-08 w=1.8e-07 $X=38359 $Y=19609 $D=616
M1429 vss 523 1129 vss hvtnfet l=6e-08 w=1.8e-07 $X=38359 $Y=24063 $D=616
M1430 vss 521 523 vss hvtnfet l=6e-08 w=1.37e-07 $X=38359 $Y=24732 $D=616
M1431 vss 522 525 vss hvtnfet l=6e-08 w=1.37e-07 $X=38359 $Y=25903 $D=616
M1432 vss 525 1130 vss hvtnfet l=6e-08 w=1.8e-07 $X=38359 $Y=26529 $D=616
M1433 779 494 vss vss hvtnfet l=6e-08 w=3.2e-07 $X=38431 $Y=32828 $D=616
M1434 780 526 vss vss hvtnfet l=1.4e-07 w=3.2e-07 $X=38481 $Y=37127 $D=616
M1435 534 495 vss vss hvtnfet l=6e-08 w=5.49e-07 $X=38515 $Y=30668 $D=616
M1436 vss 533 546 vss hvtnfet l=6e-08 w=2.74e-07 $X=38574 $Y=13476 $D=616
M1437 b_pxaa<0> 527 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=38690 $Y=336 $D=616
M1438 527 528 vss vss hvtnfet l=6e-08 w=5e-07 $X=38690 $Y=6701 $D=616
M1439 528 529 vss vss hvtnfet l=6e-08 w=3e-07 $X=38690 $Y=7831 $D=616
M1440 1131 497 529 vss hvtnfet l=6e-08 w=4.11e-07 $X=38690 $Y=11276 $D=616
M1441 1132 498 530 vss hvtnfet l=6e-08 w=4.11e-07 $X=38690 $Y=39446 $D=616
M1442 531 530 vss vss hvtnfet l=6e-08 w=3e-07 $X=38690 $Y=43002 $D=616
M1443 532 531 vss vss hvtnfet l=6e-08 w=5e-07 $X=38690 $Y=43932 $D=616
M1444 t_pxaa<0> 532 vss vss hvtnfet l=6e-08 w=1.285e-06 $X=38690 $Y=49512 $D=616
M1445 vss 527 b_pxaa<0> vss hvtnfet l=6e-08 w=1.285e-06 $X=38950 $Y=336 $D=616
M1446 vss 528 527 vss hvtnfet l=6e-08 w=5e-07 $X=38950 $Y=6701 $D=616
M1447 vss 529 528 vss hvtnfet l=6e-08 w=3e-07 $X=38950 $Y=7831 $D=616
M1448 vss 525 1131 vss hvtnfet l=6e-08 w=4.11e-07 $X=38950 $Y=11276 $D=616
M1449 vss 525 1132 vss hvtnfet l=6e-08 w=4.11e-07 $X=38950 $Y=39446 $D=616
M1450 vss 530 531 vss hvtnfet l=6e-08 w=3e-07 $X=38950 $Y=43002 $D=616
M1451 vss 531 532 vss hvtnfet l=6e-08 w=5e-07 $X=38950 $Y=43932 $D=616
M1452 vss 532 t_pxaa<0> vss hvtnfet l=6e-08 w=1.285e-06 $X=38950 $Y=49512 $D=616
M1453 vss 534 495 vss hvtnfet l=6e-08 w=5.49e-07 $X=39025 $Y=30668 $D=616
M1454 533 aa<3> vss vss hvtnfet l=6e-08 w=2.74e-07 $X=39084 $Y=13476 $D=616
M1455 vss clka 323 vss hvtnfet l=6e-08 w=6e-07 $X=39174 $Y=32403 $D=616
M1456 293 535 vss vss hvtnfet l=6e-08 w=6e-07 $X=39185 $Y=37277 $D=616
M1457 495 539 vss vss hvtnfet l=6e-08 w=5.49e-07 $X=39285 $Y=30668 $D=616
M1458 1133 537 549 vss hvtnfet l=6e-08 w=5.49e-07 $X=39379 $Y=17143 $D=616
M1459 1134 538 550 vss hvtnfet l=6e-08 w=5.49e-07 $X=39379 $Y=19240 $D=616
M1460 1135 537 551 vss hvtnfet l=6e-08 w=5.49e-07 $X=39379 $Y=24063 $D=616
M1461 1136 538 552 vss hvtnfet l=6e-08 w=5.49e-07 $X=39379 $Y=26160 $D=616
M1462 323 clka vss vss hvtnfet l=6e-08 w=6e-07 $X=39434 $Y=32403 $D=616
M1463 vss 538 537 vss hvtnfet l=6e-08 w=2.74e-07 $X=39594 $Y=13476 $D=616
M1464 1137 546 1133 vss hvtnfet l=6e-08 w=5.49e-07 $X=39639 $Y=17143 $D=616
M1465 1138 546 1134 vss hvtnfet l=6e-08 w=5.49e-07 $X=39639 $Y=19240 $D=616
M1466 1139 533 1135 vss hvtnfet l=6e-08 w=5.49e-07 $X=39639 $Y=24063 $D=616
M1467 1140 533 1136 vss hvtnfet l=6e-08 w=5.49e-07 $X=39639 $Y=26160 $D=616
M1468 r_sa_prea_n 293 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=39695 $Y=37027 $D=616
M1469 289 540 vss vss hvtnfet l=6e-08 w=6e-07 $X=39705 $Y=336 $D=616
M1470 290 541 vss vss hvtnfet l=6e-08 w=6e-07 $X=39705 $Y=5566 $D=616
M1471 291 542 vss vss hvtnfet l=6e-08 w=6e-07 $X=39705 $Y=6796 $D=616
M1472 292 543 vss vss hvtnfet l=6e-08 w=6e-07 $X=39705 $Y=12026 $D=616
M1473 294 543 vss vss hvtnfet l=6e-08 w=6e-07 $X=39705 $Y=38507 $D=616
M1474 295 542 vss vss hvtnfet l=6e-08 w=6e-07 $X=39705 $Y=43737 $D=616
M1475 296 544 vss vss hvtnfet l=6e-08 w=6e-07 $X=39705 $Y=44967 $D=616
M1476 297 545 vss vss hvtnfet l=6e-08 w=6e-07 $X=39705 $Y=50197 $D=616
M1477 vss stclka 539 vss hvtnfet l=6e-08 w=2.74e-07 $X=39795 $Y=30668 $D=616
M1478 vss 323 1137 vss hvtnfet l=6e-08 w=8.23e-07 $X=39909 $Y=17143 $D=616
M1479 vss 323 1138 vss hvtnfet l=6e-08 w=8.23e-07 $X=39909 $Y=18966 $D=616
M1480 vss 323 1139 vss hvtnfet l=6e-08 w=8.23e-07 $X=39909 $Y=24063 $D=616
M1481 vss 323 1140 vss hvtnfet l=6e-08 w=8.23e-07 $X=39909 $Y=25886 $D=616
M1482 vss 293 r_sa_prea_n vss hvtnfet l=6e-08 w=8.58e-07 $X=39955 $Y=37027 $D=616
M1483 538 aa<2> vss vss hvtnfet l=6e-08 w=2.74e-07 $X=40104 $Y=13476 $D=616
M1484 rb_ca<1> 289 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=40215 $Y=328 $D=616
M1485 rb_ca<3> 290 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=40215 $Y=5316 $D=616
M1486 rb_ma<1> 291 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=40215 $Y=6788 $D=616
M1487 rb_ma<3> 292 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=40215 $Y=11776 $D=616
M1488 r_sa_prea_n 293 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=40215 $Y=37027 $D=616
M1489 rt_ma<3> 294 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=40215 $Y=38499 $D=616
M1490 rt_ma<1> 295 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=40215 $Y=43487 $D=616
M1491 rt_ca<3> 296 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=40215 $Y=44959 $D=616
M1492 rt_ca<1> 297 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=40215 $Y=49947 $D=616
M1493 1141 317 549 vss hvtnfet l=6e-08 w=1.8e-07 $X=40419 $Y=17143 $D=616
M1494 543 549 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=40419 $Y=17812 $D=616
M1495 553 550 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=40419 $Y=18983 $D=616
M1496 1142 317 550 vss hvtnfet l=6e-08 w=1.8e-07 $X=40419 $Y=19609 $D=616
M1497 1143 317 551 vss hvtnfet l=6e-08 w=1.8e-07 $X=40419 $Y=24063 $D=616
M1498 542 551 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=40419 $Y=24732 $D=616
M1499 554 552 vss vss hvtnfet l=6e-08 w=1.37e-07 $X=40419 $Y=25903 $D=616
M1500 1144 317 552 vss hvtnfet l=6e-08 w=1.8e-07 $X=40419 $Y=26529 $D=616
M1501 vss 289 rb_ca<1> vss hvtnfet l=6e-08 w=8.58e-07 $X=40475 $Y=328 $D=616
M1502 vss 290 rb_ca<3> vss hvtnfet l=6e-08 w=8.58e-07 $X=40475 $Y=5316 $D=616
M1503 vss 291 rb_ma<1> vss hvtnfet l=6e-08 w=8.58e-07 $X=40475 $Y=6788 $D=616
M1504 vss 292 rb_ma<3> vss hvtnfet l=6e-08 w=8.58e-07 $X=40475 $Y=11776 $D=616
M1505 vss 294 rt_ma<3> vss hvtnfet l=6e-08 w=8.58e-07 $X=40475 $Y=38499 $D=616
M1506 vss 295 rt_ma<1> vss hvtnfet l=6e-08 w=8.58e-07 $X=40475 $Y=43487 $D=616
M1507 vss 296 rt_ca<3> vss hvtnfet l=6e-08 w=8.58e-07 $X=40475 $Y=44959 $D=616
M1508 vss 297 rt_ca<1> vss hvtnfet l=6e-08 w=8.58e-07 $X=40475 $Y=49947 $D=616
M1509 vss 543 1141 vss hvtnfet l=6e-08 w=1.8e-07 $X=40679 $Y=17143 $D=616
M1510 vss 549 543 vss hvtnfet l=6e-08 w=1.37e-07 $X=40679 $Y=17812 $D=616
M1511 vss 550 553 vss hvtnfet l=6e-08 w=1.37e-07 $X=40679 $Y=18983 $D=616
M1512 vss 553 1142 vss hvtnfet l=6e-08 w=1.8e-07 $X=40679 $Y=19609 $D=616
M1513 vss 542 1143 vss hvtnfet l=6e-08 w=1.8e-07 $X=40679 $Y=24063 $D=616
M1514 vss 551 542 vss hvtnfet l=6e-08 w=1.37e-07 $X=40679 $Y=24732 $D=616
M1515 vss 552 554 vss hvtnfet l=6e-08 w=1.37e-07 $X=40679 $Y=25903 $D=616
M1516 vss 554 1144 vss hvtnfet l=6e-08 w=1.8e-07 $X=40679 $Y=26529 $D=616
M1517 vss 303 r_saea_n vss hvtnfet l=6e-08 w=8.58e-07 $X=40725 $Y=37027 $D=616
M1518 rb_ca<1> 289 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=40735 $Y=328 $D=616
M1519 rb_ca<3> 290 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=40735 $Y=5316 $D=616
M1520 rb_ma<1> 291 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=40735 $Y=6788 $D=616
M1521 rb_ma<3> 292 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=40735 $Y=11776 $D=616
M1522 rt_ma<3> 294 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=40735 $Y=38499 $D=616
M1523 rt_ma<1> 295 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=40735 $Y=43487 $D=616
M1524 rt_ca<3> 296 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=40735 $Y=44959 $D=616
M1525 rt_ca<1> 297 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=40735 $Y=49947 $D=616
M1526 r_saea_n 303 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=40985 $Y=37027 $D=616
M1527 vss 299 rb_ca<0> vss hvtnfet l=6e-08 w=8.58e-07 $X=41245 $Y=328 $D=616
M1528 vss 300 rb_ca<2> vss hvtnfet l=6e-08 w=8.58e-07 $X=41245 $Y=5316 $D=616
M1529 vss 301 rb_ma<0> vss hvtnfet l=6e-08 w=8.58e-07 $X=41245 $Y=6788 $D=616
M1530 vss 302 rb_ma<2> vss hvtnfet l=6e-08 w=8.58e-07 $X=41245 $Y=11776 $D=616
M1531 vss 303 r_saea_n vss hvtnfet l=6e-08 w=8.58e-07 $X=41245 $Y=37027 $D=616
M1532 vss 304 rt_ma<2> vss hvtnfet l=6e-08 w=8.58e-07 $X=41245 $Y=38499 $D=616
M1533 vss 305 rt_ma<0> vss hvtnfet l=6e-08 w=8.58e-07 $X=41245 $Y=43487 $D=616
M1534 vss 306 rt_ca<2> vss hvtnfet l=6e-08 w=8.58e-07 $X=41245 $Y=44959 $D=616
M1535 vss 307 rt_ca<0> vss hvtnfet l=6e-08 w=8.58e-07 $X=41245 $Y=49947 $D=616
M1536 vss clka 287 vss hvtnfet l=6e-08 w=1.05e-06 $X=41495 $Y=22251 $D=616
M1537 vss 340 288 vss hvtnfet l=6e-08 w=1.05e-06 $X=41495 $Y=29007 $D=616
M1538 rb_ca<0> 299 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=41505 $Y=328 $D=616
M1539 rb_ca<2> 300 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=41505 $Y=5316 $D=616
M1540 rb_ma<0> 301 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=41505 $Y=6788 $D=616
M1541 rb_ma<2> 302 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=41505 $Y=11776 $D=616
M1542 285 497 vss vss hvtnfet l=6e-08 w=6e-07 $X=41505 $Y=13282 $D=616
M1543 286 498 vss vss hvtnfet l=6e-08 w=6e-07 $X=41505 $Y=20809 $D=616
M1544 r_saea_n 303 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=41505 $Y=37027 $D=616
M1545 rt_ma<2> 304 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=41505 $Y=38499 $D=616
M1546 rt_ma<0> 305 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=41505 $Y=43487 $D=616
M1547 rt_ca<2> 306 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=41505 $Y=44959 $D=616
M1548 rt_ca<0> 307 vss vss hvtnfet l=6e-08 w=8.58e-07 $X=41505 $Y=49947 $D=616
M1549 r_clk_dqa 287 vss vss hvtnfet l=6e-08 w=1.26e-06 $X=41755 $Y=22041 $D=616
M1550 r_clk_dqa_n 288 vss vss hvtnfet l=6e-08 w=1.26e-06 $X=41755 $Y=29007 $D=616
M1551 vss 299 rb_ca<0> vss hvtnfet l=6e-08 w=8.58e-07 $X=41765 $Y=328 $D=616
M1552 vss 300 rb_ca<2> vss hvtnfet l=6e-08 w=8.58e-07 $X=41765 $Y=5316 $D=616
M1553 vss 301 rb_ma<0> vss hvtnfet l=6e-08 w=8.58e-07 $X=41765 $Y=6788 $D=616
M1554 vss 302 rb_ma<2> vss hvtnfet l=6e-08 w=8.58e-07 $X=41765 $Y=11776 $D=616
M1555 vss 303 r_saea_n vss hvtnfet l=6e-08 w=8.58e-07 $X=41765 $Y=37027 $D=616
M1556 vss 304 rt_ma<2> vss hvtnfet l=6e-08 w=8.58e-07 $X=41765 $Y=38499 $D=616
M1557 vss 305 rt_ma<0> vss hvtnfet l=6e-08 w=8.58e-07 $X=41765 $Y=43487 $D=616
M1558 vss 306 rt_ca<2> vss hvtnfet l=6e-08 w=8.58e-07 $X=41765 $Y=44959 $D=616
M1559 vss 307 rt_ca<0> vss hvtnfet l=6e-08 w=8.58e-07 $X=41765 $Y=49947 $D=616
M1560 rb_tm_prea_n 285 vss vss hvtnfet l=6e-08 w=1.287e-06 $X=42015 $Y=13280 $D=616
M1561 rt_tm_prea_n 286 vss vss hvtnfet l=6e-08 w=1.287e-06 $X=42015 $Y=20124 $D=616
M1562 vss 287 r_clk_dqa vss hvtnfet l=6e-08 w=1.26e-06 $X=42015 $Y=22041 $D=616
M1563 vss 288 r_clk_dqa_n vss hvtnfet l=6e-08 w=1.26e-06 $X=42015 $Y=29007 $D=616
M1564 r_lwea 284 vss vss hvtnfet l=6e-08 w=1.287e-06 $X=42015 $Y=30897 $D=616
M1565 vss 555 299 vss hvtnfet l=6e-08 w=6e-07 $X=42275 $Y=336 $D=616
M1566 vss 556 300 vss hvtnfet l=6e-08 w=6e-07 $X=42275 $Y=5566 $D=616
M1567 vss 554 301 vss hvtnfet l=6e-08 w=6e-07 $X=42275 $Y=6796 $D=616
M1568 vss 553 302 vss hvtnfet l=6e-08 w=6e-07 $X=42275 $Y=12026 $D=616
M1569 vss 285 rb_tm_prea_n vss hvtnfet l=6e-08 w=1.287e-06 $X=42275 $Y=13280 $D=616
M1570 vss 286 rt_tm_prea_n vss hvtnfet l=6e-08 w=1.287e-06 $X=42275 $Y=20124 $D=616
M1571 r_clk_dqa 287 vss vss hvtnfet l=6e-08 w=1.26e-06 $X=42275 $Y=22041 $D=616
M1572 r_clk_dqa_n 288 vss vss hvtnfet l=6e-08 w=1.26e-06 $X=42275 $Y=29007 $D=616
M1573 vss 284 r_lwea vss hvtnfet l=6e-08 w=1.287e-06 $X=42275 $Y=30897 $D=616
M1574 vss 557 303 vss hvtnfet l=6e-08 w=6e-07 $X=42275 $Y=37277 $D=616
M1575 vss 553 304 vss hvtnfet l=6e-08 w=6e-07 $X=42275 $Y=38507 $D=616
M1576 vss 554 305 vss hvtnfet l=6e-08 w=6e-07 $X=42275 $Y=43737 $D=616
M1577 vss 558 306 vss hvtnfet l=6e-08 w=6e-07 $X=42275 $Y=44967 $D=616
M1578 vss 559 307 vss hvtnfet l=6e-08 w=6e-07 $X=42275 $Y=50197 $D=616
M1579 303 557 vss vss hvtnfet l=6e-08 w=6e-07 $X=42535 $Y=37277 $D=616
M1580 vdd 5 15 vdd hvtpfet l=6e-08 w=1.2e-06 $X=965 $Y=35277 $D=636
M1581 11 1 vdd vdd hvtpfet l=6e-08 w=1.2e-06 $X=1225 $Y=1736 $D=636
M1582 12 2 vdd vdd hvtpfet l=6e-08 w=1.2e-06 $X=1225 $Y=3566 $D=636
M1583 13 3 vdd vdd hvtpfet l=6e-08 w=1.2e-06 $X=1225 $Y=8196 $D=636
M1584 14 4 vdd vdd hvtpfet l=6e-08 w=1.2e-06 $X=1225 $Y=10026 $D=636
M1585 lb_tm_preb_n 20 vdd vdd hvtpfet l=6e-08 w=2.145e-06 $X=1225 $Y=14887 $D=636
M1586 lt_tm_preb_n 21 vdd vdd hvtpfet l=6e-08 w=2.145e-06 $X=1225 $Y=17659 $D=636
M1587 vdd 8 l_clk_dqb vdd hvtpfet l=6e-08 w=2.1e-06 $X=1225 $Y=23621 $D=636
M1588 vdd 9 l_clk_dqb_n vdd hvtpfet l=6e-08 w=2.1e-06 $X=1225 $Y=26587 $D=636
M1589 l_lweb 10 vdd vdd hvtpfet l=6e-08 w=2.145e-06 $X=1225 $Y=32504 $D=636
M1590 15 5 vdd vdd hvtpfet l=6e-08 w=1.2e-06 $X=1225 $Y=35277 $D=636
M1591 16 4 vdd vdd hvtpfet l=6e-08 w=1.2e-06 $X=1225 $Y=39907 $D=636
M1592 17 3 vdd vdd hvtpfet l=6e-08 w=1.2e-06 $X=1225 $Y=41737 $D=636
M1593 18 6 vdd vdd hvtpfet l=6e-08 w=1.2e-06 $X=1225 $Y=46367 $D=636
M1594 19 7 vdd vdd hvtpfet l=6e-08 w=1.2e-06 $X=1225 $Y=48197 $D=636
M1595 vdd 20 lb_tm_preb_n vdd hvtpfet l=6e-08 w=2.145e-06 $X=1485 $Y=14887 $D=636
M1596 vdd 21 lt_tm_preb_n vdd hvtpfet l=6e-08 w=2.145e-06 $X=1485 $Y=17659 $D=636
M1597 l_clk_dqb 8 vdd vdd hvtpfet l=6e-08 w=2.1e-06 $X=1485 $Y=23621 $D=636
M1598 l_clk_dqb_n 9 vdd vdd hvtpfet l=6e-08 w=2.1e-06 $X=1485 $Y=26587 $D=636
M1599 vdd 10 l_lweb vdd hvtpfet l=6e-08 w=2.145e-06 $X=1485 $Y=32504 $D=636
M1600 lb_cb<0> 11 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=1735 $Y=1506 $D=636
M1601 lb_cb<2> 12 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=1735 $Y=3566 $D=636
M1602 lb_mb<0> 13 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=1735 $Y=7966 $D=636
M1603 lb_mb<2> 14 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=1735 $Y=10026 $D=636
M1604 l_saeb_n 15 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=1735 $Y=35277 $D=636
M1605 lt_mb<2> 16 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=1735 $Y=39677 $D=636
M1606 lt_mb<0> 17 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=1735 $Y=41737 $D=636
M1607 lt_cb<2> 18 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=1735 $Y=46137 $D=636
M1608 lt_cb<0> 19 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=1735 $Y=48197 $D=636
M1609 vdd 8 l_clk_dqb vdd hvtpfet l=6e-08 w=2.1e-06 $X=1745 $Y=23621 $D=636
M1610 vdd 9 l_clk_dqb_n vdd hvtpfet l=6e-08 w=2.1e-06 $X=1745 $Y=26587 $D=636
M1611 vdd 11 lb_cb<0> vdd hvtpfet l=6e-08 w=1.43e-06 $X=1995 $Y=1506 $D=636
M1612 vdd 12 lb_cb<2> vdd hvtpfet l=6e-08 w=1.43e-06 $X=1995 $Y=3566 $D=636
M1613 vdd 13 lb_mb<0> vdd hvtpfet l=6e-08 w=1.43e-06 $X=1995 $Y=7966 $D=636
M1614 vdd 14 lb_mb<2> vdd hvtpfet l=6e-08 w=1.43e-06 $X=1995 $Y=10026 $D=636
M1615 vdd 24 20 vdd hvtpfet l=6e-08 w=1.2e-06 $X=1995 $Y=15067 $D=636
M1616 vdd 25 21 vdd hvtpfet l=6e-08 w=1.2e-06 $X=1995 $Y=18424 $D=636
M1617 vdd 15 l_saeb_n vdd hvtpfet l=6e-08 w=1.43e-06 $X=1995 $Y=35277 $D=636
M1618 vdd 16 lt_mb<2> vdd hvtpfet l=6e-08 w=1.43e-06 $X=1995 $Y=39677 $D=636
M1619 vdd 17 lt_mb<0> vdd hvtpfet l=6e-08 w=1.43e-06 $X=1995 $Y=41737 $D=636
M1620 vdd 18 lt_cb<2> vdd hvtpfet l=6e-08 w=1.43e-06 $X=1995 $Y=46137 $D=636
M1621 vdd 19 lt_cb<0> vdd hvtpfet l=6e-08 w=1.43e-06 $X=1995 $Y=48197 $D=636
M1622 8 clkb vdd vdd hvtpfet l=6e-08 w=2.1e-06 $X=2005 $Y=23621 $D=636
M1623 9 23 vdd vdd hvtpfet l=6e-08 w=2.1e-06 $X=2005 $Y=26587 $D=636
M1624 lb_cb<0> 11 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=2255 $Y=1506 $D=636
M1625 lb_cb<2> 12 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=2255 $Y=3566 $D=636
M1626 lb_mb<0> 13 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=2255 $Y=7966 $D=636
M1627 lb_mb<2> 14 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=2255 $Y=10026 $D=636
M1628 l_saeb_n 15 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=2255 $Y=35277 $D=636
M1629 lt_mb<2> 16 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=2255 $Y=39677 $D=636
M1630 lt_mb<0> 17 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=2255 $Y=41737 $D=636
M1631 lt_cb<2> 18 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=2255 $Y=46137 $D=636
M1632 lt_cb<0> 19 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=2255 $Y=48197 $D=636
M1633 vdd 15 l_saeb_n vdd hvtpfet l=6e-08 w=1.43e-06 $X=2515 $Y=35277 $D=636
M1634 vdd 34 lb_cb<1> vdd hvtpfet l=6e-08 w=1.43e-06 $X=2765 $Y=1506 $D=636
M1635 vdd 35 lb_cb<3> vdd hvtpfet l=6e-08 w=1.43e-06 $X=2765 $Y=3566 $D=636
M1636 vdd 36 lb_mb<1> vdd hvtpfet l=6e-08 w=1.43e-06 $X=2765 $Y=7966 $D=636
M1637 vdd 37 lb_mb<3> vdd hvtpfet l=6e-08 w=1.43e-06 $X=2765 $Y=10026 $D=636
M1638 vdd 39 lt_mb<3> vdd hvtpfet l=6e-08 w=1.43e-06 $X=2765 $Y=39677 $D=636
M1639 vdd 40 lt_mb<1> vdd hvtpfet l=6e-08 w=1.43e-06 $X=2765 $Y=41737 $D=636
M1640 vdd 41 lt_cb<3> vdd hvtpfet l=6e-08 w=1.43e-06 $X=2765 $Y=46137 $D=636
M1641 vdd 42 lt_cb<1> vdd hvtpfet l=6e-08 w=1.43e-06 $X=2765 $Y=48197 $D=636
M1642 l_saeb_n 15 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=2775 $Y=35277 $D=636
M1643 26 28 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=2821 $Y=15321 $D=636
M1644 1145 26 vdd vdd hvtpfet l=6e-08 w=2.74e-07 $X=2821 $Y=16069 $D=636
M1645 1146 4 vdd vdd hvtpfet l=6e-08 w=2.74e-07 $X=2821 $Y=20589 $D=636
M1646 4 29 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=2821 $Y=21405 $D=636
M1647 27 30 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=2821 $Y=22241 $D=636
M1648 1147 27 vdd vdd hvtpfet l=6e-08 w=2.74e-07 $X=2821 $Y=22989 $D=636
M1649 1148 3 vdd vdd hvtpfet l=6e-08 w=2.74e-07 $X=2821 $Y=27509 $D=636
M1650 3 31 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=2821 $Y=28325 $D=636
M1651 lb_cb<1> 34 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=3025 $Y=1506 $D=636
M1652 lb_cb<3> 35 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=3025 $Y=3566 $D=636
M1653 lb_mb<1> 36 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=3025 $Y=7966 $D=636
M1654 lb_mb<3> 37 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=3025 $Y=10026 $D=636
M1655 lt_mb<3> 39 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=3025 $Y=39677 $D=636
M1656 lt_mb<1> 40 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=3025 $Y=41737 $D=636
M1657 lt_cb<3> 41 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=3025 $Y=46137 $D=636
M1658 lt_cb<1> 42 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=3025 $Y=48197 $D=636
M1659 vdd 28 26 vdd hvtpfet l=6e-08 w=2.06e-07 $X=3081 $Y=15321 $D=636
M1660 28 43 1145 vdd hvtpfet l=6e-08 w=2.74e-07 $X=3081 $Y=16069 $D=636
M1661 29 43 1146 vdd hvtpfet l=6e-08 w=2.74e-07 $X=3081 $Y=20589 $D=636
M1662 vdd 29 4 vdd hvtpfet l=6e-08 w=2.06e-07 $X=3081 $Y=21405 $D=636
M1663 vdd 30 27 vdd hvtpfet l=6e-08 w=2.06e-07 $X=3081 $Y=22241 $D=636
M1664 30 43 1147 vdd hvtpfet l=6e-08 w=2.74e-07 $X=3081 $Y=22989 $D=636
M1665 31 43 1148 vdd hvtpfet l=6e-08 w=2.74e-07 $X=3081 $Y=27509 $D=636
M1666 vdd 31 3 vdd hvtpfet l=6e-08 w=2.06e-07 $X=3081 $Y=28325 $D=636
M1667 vdd 34 lb_cb<1> vdd hvtpfet l=6e-08 w=1.43e-06 $X=3285 $Y=1506 $D=636
M1668 vdd 35 lb_cb<3> vdd hvtpfet l=6e-08 w=1.43e-06 $X=3285 $Y=3566 $D=636
M1669 vdd 36 lb_mb<1> vdd hvtpfet l=6e-08 w=1.43e-06 $X=3285 $Y=7966 $D=636
M1670 vdd 37 lb_mb<3> vdd hvtpfet l=6e-08 w=1.43e-06 $X=3285 $Y=10026 $D=636
M1671 vdd 51 l_sa_preb_n vdd hvtpfet l=6e-08 w=1.43e-06 $X=3285 $Y=35277 $D=636
M1672 vdd 39 lt_mb<3> vdd hvtpfet l=6e-08 w=1.43e-06 $X=3285 $Y=39677 $D=636
M1673 vdd 40 lt_mb<1> vdd hvtpfet l=6e-08 w=1.43e-06 $X=3285 $Y=41737 $D=636
M1674 vdd 41 lt_cb<3> vdd hvtpfet l=6e-08 w=1.43e-06 $X=3285 $Y=46137 $D=636
M1675 vdd 42 lt_cb<1> vdd hvtpfet l=6e-08 w=1.43e-06 $X=3285 $Y=48197 $D=636
M1676 vdd ab<2> 44 vdd hvtpfet l=6e-08 w=4.11e-07 $X=3396 $Y=14280 $D=636
M1677 l_sa_preb_n 51 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=3545 $Y=35277 $D=636
M1678 vdd clkb 43 vdd hvtpfet l=6e-08 w=6e-07 $X=3546 $Y=33747 $D=636
M1679 1149 33 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=3591 $Y=15520 $D=636
M1680 1150 33 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=3591 $Y=20589 $D=636
M1681 1151 33 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=3591 $Y=22440 $D=636
M1682 1152 33 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=3591 $Y=27509 $D=636
M1683 52 stclkb vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=3705 $Y=29937 $D=636
M1684 vdd 47 34 vdd hvtpfet l=6e-08 w=1.2e-06 $X=3795 $Y=1736 $D=636
M1685 vdd 48 35 vdd hvtpfet l=6e-08 w=1.2e-06 $X=3795 $Y=3566 $D=636
M1686 vdd 27 36 vdd hvtpfet l=6e-08 w=1.2e-06 $X=3795 $Y=8196 $D=636
M1687 vdd 26 37 vdd hvtpfet l=6e-08 w=1.2e-06 $X=3795 $Y=10026 $D=636
M1688 vdd 26 39 vdd hvtpfet l=6e-08 w=1.2e-06 $X=3795 $Y=39907 $D=636
M1689 vdd 27 40 vdd hvtpfet l=6e-08 w=1.2e-06 $X=3795 $Y=41737 $D=636
M1690 vdd 49 41 vdd hvtpfet l=6e-08 w=1.2e-06 $X=3795 $Y=46367 $D=636
M1691 vdd 50 42 vdd hvtpfet l=6e-08 w=1.2e-06 $X=3795 $Y=48197 $D=636
M1692 vdd 51 l_sa_preb_n vdd hvtpfet l=6e-08 w=1.43e-06 $X=3805 $Y=35277 $D=636
M1693 43 clkb vdd vdd hvtpfet l=6e-08 w=6e-07 $X=3806 $Y=33747 $D=636
M1694 28 45 1149 vdd hvtpfet l=6e-08 w=4.11e-07 $X=3861 $Y=15932 $D=636
M1695 29 45 1150 vdd hvtpfet l=6e-08 w=4.11e-07 $X=3861 $Y=20589 $D=636
M1696 30 46 1151 vdd hvtpfet l=6e-08 w=4.11e-07 $X=3861 $Y=22852 $D=636
M1697 31 46 1152 vdd hvtpfet l=6e-08 w=4.11e-07 $X=3861 $Y=27509 $D=636
M1698 53 44 vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=3906 $Y=14280 $D=636
M1699 vdd clkb 43 vdd hvtpfet l=6e-08 w=6e-07 $X=4066 $Y=33747 $D=636
M1700 1153 53 28 vdd hvtpfet l=6e-08 w=4.11e-07 $X=4121 $Y=15932 $D=636
M1701 1154 44 29 vdd hvtpfet l=6e-08 w=4.11e-07 $X=4121 $Y=20589 $D=636
M1702 1155 53 30 vdd hvtpfet l=6e-08 w=4.11e-07 $X=4121 $Y=22852 $D=636
M1703 1156 44 31 vdd hvtpfet l=6e-08 w=4.11e-07 $X=4121 $Y=27509 $D=636
M1704 1157 52 59 vdd hvtpfet l=6e-08 w=8.23e-07 $X=4215 $Y=29525 $D=636
M1705 vdd 55 51 vdd hvtpfet l=6e-08 w=1.2e-06 $X=4315 $Y=35277 $D=636
M1706 43 clkb vdd vdd hvtpfet l=6e-08 w=6e-07 $X=4326 $Y=33747 $D=636
M1707 vdd 33 1153 vdd hvtpfet l=6e-08 w=8.23e-07 $X=4391 $Y=15520 $D=636
M1708 vdd 33 1154 vdd hvtpfet l=6e-08 w=8.23e-07 $X=4391 $Y=20589 $D=636
M1709 vdd 33 1155 vdd hvtpfet l=6e-08 w=8.23e-07 $X=4391 $Y=22440 $D=636
M1710 vdd 33 1156 vdd hvtpfet l=6e-08 w=8.23e-07 $X=4391 $Y=27509 $D=636
M1711 vdd ab<3> 46 vdd hvtpfet l=6e-08 w=4.11e-07 $X=4416 $Y=14280 $D=636
M1712 vdd 56 1157 vdd hvtpfet l=6e-08 w=8.23e-07 $X=4475 $Y=29525 $D=636
M1713 b_pxab<0> 60 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=4550 $Y=1941 $D=636
M1714 60 61 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=4550 $Y=5141 $D=636
M1715 61 62 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=4550 $Y=8691 $D=636
M1716 vdd 57 62 vdd hvtpfet l=6e-08 w=4.11e-07 $X=4550 $Y=10156 $D=636
M1717 vdd 57 63 vdd hvtpfet l=6e-08 w=4.11e-07 $X=4550 $Y=40566 $D=636
M1718 64 63 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=4550 $Y=41842 $D=636
M1719 65 64 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=4550 $Y=44992 $D=636
M1720 t_pxab<0> 65 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=4550 $Y=46622 $D=636
M1721 vdd 60 b_pxab<0> vdd hvtpfet l=6e-08 w=2.57e-06 $X=4810 $Y=1941 $D=636
M1722 vdd 61 60 vdd hvtpfet l=6e-08 w=1e-06 $X=4810 $Y=5141 $D=636
M1723 vdd 62 61 vdd hvtpfet l=6e-08 w=6e-07 $X=4810 $Y=8691 $D=636
M1724 62 24 vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=4810 $Y=10156 $D=636
M1725 63 25 vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=4810 $Y=40566 $D=636
M1726 vdd 63 64 vdd hvtpfet l=6e-08 w=6e-07 $X=4810 $Y=41842 $D=636
M1727 vdd 64 65 vdd hvtpfet l=6e-08 w=1e-06 $X=4810 $Y=44992 $D=636
M1728 vdd 65 t_pxab<0> vdd hvtpfet l=6e-08 w=2.57e-06 $X=4810 $Y=46622 $D=636
M1729 45 46 vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=4926 $Y=14280 $D=636
M1730 vdd 66 586 vdd hvtpfet l=1.4e-07 w=6.4e-07 $X=4939 $Y=36067 $D=636
M1731 1158 59 56 vdd hvtpfet l=6e-08 w=8.23e-07 $X=4985 $Y=29525 $D=636
M1732 vdd 58 587 vdd hvtpfet l=6e-08 w=6.4e-07 $X=5069 $Y=33468 $D=636
M1733 67 73 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=5141 $Y=15321 $D=636
M1734 1159 67 vdd vdd hvtpfet l=6e-08 w=2.74e-07 $X=5141 $Y=16069 $D=636
M1735 1160 68 vdd vdd hvtpfet l=6e-08 w=2.74e-07 $X=5141 $Y=20589 $D=636
M1736 68 74 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=5141 $Y=21405 $D=636
M1737 69 75 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=5141 $Y=22241 $D=636
M1738 1161 69 vdd vdd hvtpfet l=6e-08 w=2.74e-07 $X=5141 $Y=22989 $D=636
M1739 1162 57 vdd vdd hvtpfet l=6e-08 w=2.74e-07 $X=5141 $Y=27509 $D=636
M1740 57 76 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=5141 $Y=28325 $D=636
M1741 vdd 70 1158 vdd hvtpfet l=6e-08 w=8.23e-07 $X=5245 $Y=29525 $D=636
M1742 66 71 vdd vdd hvtpfet l=1.4e-07 w=6.4e-07 $X=5279 $Y=36067 $D=636
M1743 b_pxab<1> 78 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=5320 $Y=1941 $D=636
M1744 78 79 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=5320 $Y=5141 $D=636
M1745 79 80 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=5320 $Y=8691 $D=636
M1746 vdd 24 80 vdd hvtpfet l=6e-08 w=4.11e-07 $X=5320 $Y=10156 $D=636
M1747 vdd 25 81 vdd hvtpfet l=6e-08 w=4.11e-07 $X=5320 $Y=40566 $D=636
M1748 82 81 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=5320 $Y=41842 $D=636
M1749 83 82 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=5320 $Y=44992 $D=636
M1750 t_pxab<1> 83 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=5320 $Y=46622 $D=636
M1751 vdd 73 67 vdd hvtpfet l=6e-08 w=2.06e-07 $X=5401 $Y=15321 $D=636
M1752 73 43 1159 vdd hvtpfet l=6e-08 w=2.74e-07 $X=5401 $Y=16069 $D=636
M1753 74 43 1160 vdd hvtpfet l=6e-08 w=2.74e-07 $X=5401 $Y=20589 $D=636
M1754 vdd 74 68 vdd hvtpfet l=6e-08 w=2.06e-07 $X=5401 $Y=21405 $D=636
M1755 vdd 75 69 vdd hvtpfet l=6e-08 w=2.06e-07 $X=5401 $Y=22241 $D=636
M1756 75 43 1161 vdd hvtpfet l=6e-08 w=2.74e-07 $X=5401 $Y=22989 $D=636
M1757 76 43 1162 vdd hvtpfet l=6e-08 w=2.74e-07 $X=5401 $Y=27509 $D=636
M1758 vdd 76 57 vdd hvtpfet l=6e-08 w=2.06e-07 $X=5401 $Y=28325 $D=636
M1759 vdd 72 5 vdd hvtpfet l=6e-08 w=6.4e-07 $X=5579 $Y=33693 $D=636
M1760 vdd 78 b_pxab<1> vdd hvtpfet l=6e-08 w=2.57e-06 $X=5580 $Y=1941 $D=636
M1761 vdd 79 78 vdd hvtpfet l=6e-08 w=1e-06 $X=5580 $Y=5141 $D=636
M1762 vdd 80 79 vdd hvtpfet l=6e-08 w=6e-07 $X=5580 $Y=8691 $D=636
M1763 80 69 vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=5580 $Y=10156 $D=636
M1764 81 69 vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=5580 $Y=40566 $D=636
M1765 vdd 81 82 vdd hvtpfet l=6e-08 w=6e-07 $X=5580 $Y=41842 $D=636
M1766 vdd 82 83 vdd hvtpfet l=6e-08 w=1e-06 $X=5580 $Y=44992 $D=636
M1767 vdd 83 t_pxab<1> vdd hvtpfet l=6e-08 w=2.57e-06 $X=5580 $Y=46622 $D=636
M1768 vdd ab<5> 86 vdd hvtpfet l=6e-08 w=4.11e-07 $X=5716 $Y=14280 $D=636
M1769 5 85 vdd vdd hvtpfet l=6e-08 w=6.4e-07 $X=5839 $Y=33693 $D=636
M1770 1163 33 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=5911 $Y=15520 $D=636
M1771 1164 33 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=5911 $Y=20589 $D=636
M1772 1165 33 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=5911 $Y=22440 $D=636
M1773 1166 33 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=5911 $Y=27509 $D=636
M1774 70 clkb vdd vdd hvtpfet l=6e-08 w=1.2e-06 $X=6015 $Y=29148 $D=636
M1775 592 ddqb 71 vdd hvtpfet l=6e-08 w=6.4e-07 $X=6079 $Y=35802 $D=636
M1776 b_pxab<2> 90 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=6090 $Y=1941 $D=636
M1777 90 91 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=6090 $Y=5141 $D=636
M1778 91 92 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=6090 $Y=8691 $D=636
M1779 vdd 68 92 vdd hvtpfet l=6e-08 w=4.11e-07 $X=6090 $Y=10156 $D=636
M1780 vdd 68 93 vdd hvtpfet l=6e-08 w=4.11e-07 $X=6090 $Y=40566 $D=636
M1781 94 93 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=6090 $Y=41842 $D=636
M1782 95 94 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=6090 $Y=44992 $D=636
M1783 t_pxab<2> 95 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=6090 $Y=46622 $D=636
M1784 73 87 1163 vdd hvtpfet l=6e-08 w=4.11e-07 $X=6181 $Y=15932 $D=636
M1785 74 87 1164 vdd hvtpfet l=6e-08 w=4.11e-07 $X=6181 $Y=20589 $D=636
M1786 75 88 1165 vdd hvtpfet l=6e-08 w=4.11e-07 $X=6181 $Y=22852 $D=636
M1787 76 88 1166 vdd hvtpfet l=6e-08 w=4.11e-07 $X=6181 $Y=27509 $D=636
M1788 97 86 vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=6226 $Y=14280 $D=636
M1789 vdd ddqb_n 592 vdd hvtpfet l=6e-08 w=6.4e-07 $X=6339 $Y=35802 $D=636
M1790 vdd 90 b_pxab<2> vdd hvtpfet l=6e-08 w=2.57e-06 $X=6350 $Y=1941 $D=636
M1791 vdd 91 90 vdd hvtpfet l=6e-08 w=1e-06 $X=6350 $Y=5141 $D=636
M1792 vdd 92 91 vdd hvtpfet l=6e-08 w=6e-07 $X=6350 $Y=8691 $D=636
M1793 92 24 vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=6350 $Y=10156 $D=636
M1794 93 25 vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=6350 $Y=40566 $D=636
M1795 vdd 93 94 vdd hvtpfet l=6e-08 w=6e-07 $X=6350 $Y=41842 $D=636
M1796 vdd 94 95 vdd hvtpfet l=6e-08 w=1e-06 $X=6350 $Y=44992 $D=636
M1797 vdd 95 t_pxab<2> vdd hvtpfet l=6e-08 w=2.57e-06 $X=6350 $Y=46622 $D=636
M1798 1167 97 73 vdd hvtpfet l=6e-08 w=4.11e-07 $X=6441 $Y=15932 $D=636
M1799 1168 86 74 vdd hvtpfet l=6e-08 w=4.11e-07 $X=6441 $Y=20589 $D=636
M1800 1169 97 75 vdd hvtpfet l=6e-08 w=4.11e-07 $X=6441 $Y=22852 $D=636
M1801 1170 86 76 vdd hvtpfet l=6e-08 w=4.11e-07 $X=6441 $Y=27509 $D=636
M1802 85 89 vdd vdd hvtpfet l=6e-08 w=6.4e-07 $X=6524 $Y=33693 $D=636
M1803 142 clkb vdd vdd hvtpfet l=6e-08 w=8e-07 $X=6525 $Y=29548 $D=636
M1804 vdd 33 1167 vdd hvtpfet l=6e-08 w=8.23e-07 $X=6711 $Y=15520 $D=636
M1805 vdd 33 1168 vdd hvtpfet l=6e-08 w=8.23e-07 $X=6711 $Y=20589 $D=636
M1806 vdd 33 1169 vdd hvtpfet l=6e-08 w=8.23e-07 $X=6711 $Y=22440 $D=636
M1807 vdd 33 1170 vdd hvtpfet l=6e-08 w=8.23e-07 $X=6711 $Y=27509 $D=636
M1808 vdd ab<6> 88 vdd hvtpfet l=6e-08 w=4.11e-07 $X=6736 $Y=14280 $D=636
M1809 vdd clkb 142 vdd hvtpfet l=6e-08 w=8e-07 $X=6785 $Y=29548 $D=636
M1810 b_pxab<3> 99 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=6860 $Y=1941 $D=636
M1811 99 100 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=6860 $Y=5141 $D=636
M1812 100 101 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=6860 $Y=8691 $D=636
M1813 vdd 24 101 vdd hvtpfet l=6e-08 w=4.11e-07 $X=6860 $Y=10156 $D=636
M1814 vdd 25 102 vdd hvtpfet l=6e-08 w=4.11e-07 $X=6860 $Y=40566 $D=636
M1815 103 102 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=6860 $Y=41842 $D=636
M1816 104 103 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=6860 $Y=44992 $D=636
M1817 t_pxab<3> 104 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=6860 $Y=46622 $D=636
M1818 109 85 vdd vdd hvtpfet l=6e-08 w=6.4e-07 $X=7034 $Y=33468 $D=636
M1819 89 71 vdd vdd hvtpfet l=6e-08 w=6.4e-07 $X=7069 $Y=35802 $D=636
M1820 vdd 99 b_pxab<3> vdd hvtpfet l=6e-08 w=2.57e-06 $X=7120 $Y=1941 $D=636
M1821 vdd 100 99 vdd hvtpfet l=6e-08 w=1e-06 $X=7120 $Y=5141 $D=636
M1822 vdd 101 100 vdd hvtpfet l=6e-08 w=6e-07 $X=7120 $Y=8691 $D=636
M1823 101 67 vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=7120 $Y=10156 $D=636
M1824 102 67 vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=7120 $Y=40566 $D=636
M1825 vdd 102 103 vdd hvtpfet l=6e-08 w=6e-07 $X=7120 $Y=41842 $D=636
M1826 vdd 103 104 vdd hvtpfet l=6e-08 w=1e-06 $X=7120 $Y=44992 $D=636
M1827 vdd 104 t_pxab<3> vdd hvtpfet l=6e-08 w=2.57e-06 $X=7120 $Y=46622 $D=636
M1828 87 88 vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=7246 $Y=14280 $D=636
M1829 142 59 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=7295 $Y=29548 $D=636
M1830 105 111 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=7461 $Y=15321 $D=636
M1831 1171 105 vdd vdd hvtpfet l=6e-08 w=2.74e-07 $X=7461 $Y=16069 $D=636
M1832 1172 106 vdd vdd hvtpfet l=6e-08 w=2.74e-07 $X=7461 $Y=20589 $D=636
M1833 106 112 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=7461 $Y=21405 $D=636
M1834 107 113 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=7461 $Y=22241 $D=636
M1835 1173 107 vdd vdd hvtpfet l=6e-08 w=2.74e-07 $X=7461 $Y=22989 $D=636
M1836 1174 108 vdd vdd hvtpfet l=6e-08 w=2.74e-07 $X=7461 $Y=27509 $D=636
M1837 108 114 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=7461 $Y=28325 $D=636
M1838 vdd 59 142 vdd hvtpfet l=6e-08 w=8e-07 $X=7555 $Y=29548 $D=636
M1839 vdd 110 89 vdd hvtpfet l=1.2e-07 w=3e-07 $X=7579 $Y=36382 $D=636
M1840 b_pxbb_n<0> 115 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=7630 $Y=1941 $D=636
M1841 115 116 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=7630 $Y=5141 $D=636
M1842 116 107 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=7630 $Y=8691 $D=636
M1843 117 107 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=7630 $Y=41842 $D=636
M1844 118 117 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=7630 $Y=44992 $D=636
M1845 t_pxbb_n<0> 118 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=7630 $Y=46622 $D=636
M1846 vdd 109 119 vdd hvtpfet l=6e-08 w=5e-07 $X=7634 $Y=33503 $D=636
M1847 vdd 111 105 vdd hvtpfet l=6e-08 w=2.06e-07 $X=7721 $Y=15321 $D=636
M1848 111 43 1171 vdd hvtpfet l=6e-08 w=2.74e-07 $X=7721 $Y=16069 $D=636
M1849 112 43 1172 vdd hvtpfet l=6e-08 w=2.74e-07 $X=7721 $Y=20589 $D=636
M1850 vdd 112 106 vdd hvtpfet l=6e-08 w=2.06e-07 $X=7721 $Y=21405 $D=636
M1851 vdd 113 107 vdd hvtpfet l=6e-08 w=2.06e-07 $X=7721 $Y=22241 $D=636
M1852 113 43 1173 vdd hvtpfet l=6e-08 w=2.74e-07 $X=7721 $Y=22989 $D=636
M1853 114 43 1174 vdd hvtpfet l=6e-08 w=2.74e-07 $X=7721 $Y=27509 $D=636
M1854 vdd 114 108 vdd hvtpfet l=6e-08 w=2.06e-07 $X=7721 $Y=28325 $D=636
M1855 vdd 115 b_pxbb_n<0> vdd hvtpfet l=6e-08 w=2.57e-06 $X=7890 $Y=1941 $D=636
M1856 vdd 116 115 vdd hvtpfet l=6e-08 w=1e-06 $X=7890 $Y=5141 $D=636
M1857 vdd 107 116 vdd hvtpfet l=6e-08 w=6e-07 $X=7890 $Y=8691 $D=636
M1858 vdd 107 117 vdd hvtpfet l=6e-08 w=6e-07 $X=7890 $Y=41842 $D=636
M1859 vdd 117 118 vdd hvtpfet l=6e-08 w=1e-06 $X=7890 $Y=44992 $D=636
M1860 vdd 118 t_pxbb_n<0> vdd hvtpfet l=6e-08 w=2.57e-06 $X=7890 $Y=46622 $D=636
M1861 120 119 vdd vdd hvtpfet l=2.5e-07 w=5e-07 $X=7894 $Y=33503 $D=636
M1862 110 89 vdd vdd hvtpfet l=6e-08 w=3e-07 $X=8149 $Y=36377 $D=636
M1863 1175 33 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=8231 $Y=15520 $D=636
M1864 1176 33 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=8231 $Y=20589 $D=636
M1865 1177 33 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=8231 $Y=22440 $D=636
M1866 1178 33 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=8231 $Y=27509 $D=636
M1867 b_pxbb_n<1> 125 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=8400 $Y=1941 $D=636
M1868 125 126 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=8400 $Y=5141 $D=636
M1869 126 108 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=8400 $Y=8691 $D=636
M1870 127 108 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=8400 $Y=41842 $D=636
M1871 128 127 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=8400 $Y=44992 $D=636
M1872 t_pxbb_n<1> 128 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=8400 $Y=46622 $D=636
M1873 vdd 122 121 vdd hvtpfet l=6e-08 w=4.11e-07 $X=8466 $Y=14280 $D=636
M1874 111 121 1175 vdd hvtpfet l=6e-08 w=4.11e-07 $X=8501 $Y=15932 $D=636
M1875 112 121 1176 vdd hvtpfet l=6e-08 w=4.11e-07 $X=8501 $Y=20589 $D=636
M1876 113 122 1177 vdd hvtpfet l=6e-08 w=4.11e-07 $X=8501 $Y=22852 $D=636
M1877 114 122 1178 vdd hvtpfet l=6e-08 w=4.11e-07 $X=8501 $Y=27509 $D=636
M1878 131 123 vdd vdd hvtpfet l=6e-08 w=2e-07 $X=8594 $Y=10756 $D=636
M1879 vdd 120 55 vdd hvtpfet l=6e-08 w=6.4e-07 $X=8619 $Y=33468 $D=636
M1880 602 124 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=8659 $Y=29348 $D=636
M1881 603 124 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=8659 $Y=35707 $D=636
M1882 vdd 125 b_pxbb_n<1> vdd hvtpfet l=6e-08 w=2.57e-06 $X=8660 $Y=1941 $D=636
M1883 vdd 126 125 vdd hvtpfet l=6e-08 w=1e-06 $X=8660 $Y=5141 $D=636
M1884 vdd 108 126 vdd hvtpfet l=6e-08 w=6e-07 $X=8660 $Y=8691 $D=636
M1885 vdd 108 127 vdd hvtpfet l=6e-08 w=6e-07 $X=8660 $Y=41842 $D=636
M1886 vdd 127 128 vdd hvtpfet l=6e-08 w=1e-06 $X=8660 $Y=44992 $D=636
M1887 vdd 128 t_pxbb_n<1> vdd hvtpfet l=6e-08 w=2.57e-06 $X=8660 $Y=46622 $D=636
M1888 1179 129 111 vdd hvtpfet l=6e-08 w=4.11e-07 $X=8761 $Y=15932 $D=636
M1889 1180 129 112 vdd hvtpfet l=6e-08 w=4.11e-07 $X=8761 $Y=20589 $D=636
M1890 1181 129 113 vdd hvtpfet l=6e-08 w=4.11e-07 $X=8761 $Y=22852 $D=636
M1891 1182 129 114 vdd hvtpfet l=6e-08 w=4.11e-07 $X=8761 $Y=27509 $D=636
M1892 55 vdd vdd vdd hvtpfet l=6e-08 w=6.4e-07 $X=8879 $Y=33468 $D=636
M1893 vdd 124 602 vdd hvtpfet l=6e-08 w=1e-06 $X=8919 $Y=29348 $D=636
M1894 vdd 124 603 vdd hvtpfet l=6e-08 w=1e-06 $X=8919 $Y=35707 $D=636
M1895 122 ab<9> vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=8976 $Y=14280 $D=636
M1896 vdd 33 1179 vdd hvtpfet l=6e-08 w=8.23e-07 $X=9031 $Y=15520 $D=636
M1897 vdd 33 1180 vdd hvtpfet l=6e-08 w=8.23e-07 $X=9031 $Y=20589 $D=636
M1898 vdd 33 1181 vdd hvtpfet l=6e-08 w=8.23e-07 $X=9031 $Y=22440 $D=636
M1899 vdd 33 1182 vdd hvtpfet l=6e-08 w=8.23e-07 $X=9031 $Y=27509 $D=636
M1900 b_pxbb_n<2> 135 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=9170 $Y=1941 $D=636
M1901 135 136 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=9170 $Y=5141 $D=636
M1902 136 137 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=9170 $Y=8691 $D=636
M1903 138 137 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=9170 $Y=41842 $D=636
M1904 139 138 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=9170 $Y=44992 $D=636
M1905 t_pxbb_n<2> 139 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=9170 $Y=46622 $D=636
M1906 dwlb<0> 142 602 vdd hvtpfet l=6e-08 w=1e-06 $X=9429 $Y=29348 $D=636
M1907 25 143 603 vdd hvtpfet l=6e-08 w=1e-06 $X=9429 $Y=35707 $D=636
M1908 vdd 135 b_pxbb_n<2> vdd hvtpfet l=6e-08 w=2.57e-06 $X=9430 $Y=1941 $D=636
M1909 vdd 136 135 vdd hvtpfet l=6e-08 w=1e-06 $X=9430 $Y=5141 $D=636
M1910 vdd 137 136 vdd hvtpfet l=6e-08 w=6e-07 $X=9430 $Y=8691 $D=636
M1911 vdd 137 138 vdd hvtpfet l=6e-08 w=6e-07 $X=9430 $Y=41842 $D=636
M1912 vdd 138 139 vdd hvtpfet l=6e-08 w=1e-06 $X=9430 $Y=44992 $D=636
M1913 vdd 139 t_pxbb_n<2> vdd hvtpfet l=6e-08 w=2.57e-06 $X=9430 $Y=46622 $D=636
M1914 1183 132 111 vdd hvtpfet l=6e-08 w=4.11e-07 $X=9541 $Y=15932 $D=636
M1915 1184 133 112 vdd hvtpfet l=6e-08 w=4.11e-07 $X=9541 $Y=20589 $D=636
M1916 1185 132 113 vdd hvtpfet l=6e-08 w=4.11e-07 $X=9541 $Y=22852 $D=636
M1917 1186 133 114 vdd hvtpfet l=6e-08 w=4.11e-07 $X=9541 $Y=27509 $D=636
M1918 vdd 140 1 vdd hvtpfet l=6e-08 w=4e-07 $X=9586 $Y=10167 $D=636
M1919 vdd 141 7 vdd hvtpfet l=6e-08 w=4e-07 $X=9586 $Y=40566 $D=636
M1920 602 142 dwlb<0> vdd hvtpfet l=6e-08 w=1e-06 $X=9689 $Y=29348 $D=636
M1921 603 143 25 vdd hvtpfet l=6e-08 w=1e-06 $X=9689 $Y=35707 $D=636
M1922 vdd 33 1183 vdd hvtpfet l=6e-08 w=8.23e-07 $X=9811 $Y=15520 $D=636
M1923 vdd 33 1184 vdd hvtpfet l=6e-08 w=8.23e-07 $X=9811 $Y=20589 $D=636
M1924 vdd 33 1185 vdd hvtpfet l=6e-08 w=8.23e-07 $X=9811 $Y=22440 $D=636
M1925 vdd 33 1186 vdd hvtpfet l=6e-08 w=8.23e-07 $X=9811 $Y=27509 $D=636
M1926 b_pxbb_n<3> 146 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=9940 $Y=1941 $D=636
M1927 146 147 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=9940 $Y=5141 $D=636
M1928 147 148 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=9940 $Y=8691 $D=636
M1929 149 148 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=9940 $Y=41842 $D=636
M1930 150 149 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=9940 $Y=44992 $D=636
M1931 t_pxbb_n<3> 150 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=9940 $Y=46622 $D=636
M1932 vdd ab<8> 129 vdd hvtpfet l=6e-08 w=4.11e-07 $X=9986 $Y=14280 $D=636
M1933 1187 33 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=10071 $Y=15520 $D=636
M1934 1188 33 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=10071 $Y=20589 $D=636
M1935 1189 33 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=10071 $Y=22440 $D=636
M1936 1190 33 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=10071 $Y=27509 $D=636
M1937 vdd 145 140 vdd hvtpfet l=6e-08 w=4.11e-07 $X=10096 $Y=10156 $D=636
M1938 vdd 145 141 vdd hvtpfet l=6e-08 w=4.11e-07 $X=10096 $Y=40566 $D=636
M1939 dwlb<1> 142 608 vdd hvtpfet l=6e-08 w=1e-06 $X=10199 $Y=29348 $D=636
M1940 24 143 609 vdd hvtpfet l=6e-08 w=1e-06 $X=10199 $Y=35707 $D=636
M1941 vdd 146 b_pxbb_n<3> vdd hvtpfet l=6e-08 w=2.57e-06 $X=10200 $Y=1941 $D=636
M1942 vdd 147 146 vdd hvtpfet l=6e-08 w=1e-06 $X=10200 $Y=5141 $D=636
M1943 vdd 148 147 vdd hvtpfet l=6e-08 w=6e-07 $X=10200 $Y=8691 $D=636
M1944 vdd 148 149 vdd hvtpfet l=6e-08 w=6e-07 $X=10200 $Y=41842 $D=636
M1945 vdd 149 150 vdd hvtpfet l=6e-08 w=1e-06 $X=10200 $Y=44992 $D=636
M1946 vdd 150 t_pxbb_n<3> vdd hvtpfet l=6e-08 w=2.57e-06 $X=10200 $Y=46622 $D=636
M1947 160 129 vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=10246 $Y=14280 $D=636
M1948 168 132 1187 vdd hvtpfet l=6e-08 w=4.11e-07 $X=10341 $Y=15932 $D=636
M1949 169 133 1188 vdd hvtpfet l=6e-08 w=4.11e-07 $X=10341 $Y=20589 $D=636
M1950 170 132 1189 vdd hvtpfet l=6e-08 w=4.11e-07 $X=10341 $Y=22852 $D=636
M1951 171 133 1190 vdd hvtpfet l=6e-08 w=4.11e-07 $X=10341 $Y=27509 $D=636
M1952 140 dwlb<1> vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=10356 $Y=10156 $D=636
M1953 141 dwlb<0> vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=10356 $Y=40566 $D=636
M1954 vdd 153 124 vdd hvtpfet l=6e-08 w=8e-07 $X=10406 $Y=33493 $D=636
M1955 608 142 dwlb<1> vdd hvtpfet l=6e-08 w=1e-06 $X=10459 $Y=29348 $D=636
M1956 609 143 24 vdd hvtpfet l=6e-08 w=1e-06 $X=10459 $Y=35707 $D=636
M1957 b_pxbb_n<4> 156 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=10710 $Y=1941 $D=636
M1958 156 157 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=10710 $Y=5141 $D=636
M1959 157 105 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=10710 $Y=8691 $D=636
M1960 158 105 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=10710 $Y=41842 $D=636
M1961 159 158 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=10710 $Y=44992 $D=636
M1962 t_pxbb_n<4> 159 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=10710 $Y=46622 $D=636
M1963 vdd 132 133 vdd hvtpfet l=6e-08 w=4.11e-07 $X=10846 $Y=14280 $D=636
M1964 1191 33 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=10851 $Y=15520 $D=636
M1965 1192 33 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=10851 $Y=20589 $D=636
M1966 1193 33 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=10851 $Y=22440 $D=636
M1967 1194 33 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=10851 $Y=27509 $D=636
M1968 vdd dwlb<1> 162 vdd hvtpfet l=6e-08 w=4.11e-07 $X=10866 $Y=10156 $D=636
M1969 vdd dwlb<0> 163 vdd hvtpfet l=6e-08 w=4.11e-07 $X=10866 $Y=40566 $D=636
M1970 608 153 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=10969 $Y=29348 $D=636
M1971 609 153 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=10969 $Y=35707 $D=636
M1972 vdd 156 b_pxbb_n<4> vdd hvtpfet l=6e-08 w=2.57e-06 $X=10970 $Y=1941 $D=636
M1973 vdd 157 156 vdd hvtpfet l=6e-08 w=1e-06 $X=10970 $Y=5141 $D=636
M1974 vdd 105 157 vdd hvtpfet l=6e-08 w=6e-07 $X=10970 $Y=8691 $D=636
M1975 vdd 105 158 vdd hvtpfet l=6e-08 w=6e-07 $X=10970 $Y=41842 $D=636
M1976 vdd 158 159 vdd hvtpfet l=6e-08 w=1e-06 $X=10970 $Y=44992 $D=636
M1977 vdd 159 t_pxbb_n<4> vdd hvtpfet l=6e-08 w=2.57e-06 $X=10970 $Y=46622 $D=636
M1978 132 ab<7> vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=11106 $Y=14280 $D=636
M1979 153 154 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=11106 $Y=33493 $D=636
M1980 168 160 1191 vdd hvtpfet l=6e-08 w=4.11e-07 $X=11121 $Y=15932 $D=636
M1981 169 160 1192 vdd hvtpfet l=6e-08 w=4.11e-07 $X=11121 $Y=20589 $D=636
M1982 170 160 1193 vdd hvtpfet l=6e-08 w=4.11e-07 $X=11121 $Y=22852 $D=636
M1983 171 160 1194 vdd hvtpfet l=6e-08 w=4.11e-07 $X=11121 $Y=27509 $D=636
M1984 162 155 vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=11126 $Y=10156 $D=636
M1985 163 155 vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=11126 $Y=40566 $D=636
M1986 vdd 153 608 vdd hvtpfet l=6e-08 w=1e-06 $X=11229 $Y=29348 $D=636
M1987 vdd 153 609 vdd hvtpfet l=6e-08 w=1e-06 $X=11229 $Y=35707 $D=636
M1988 1195 121 168 vdd hvtpfet l=6e-08 w=4.11e-07 $X=11381 $Y=15932 $D=636
M1989 1196 121 169 vdd hvtpfet l=6e-08 w=4.11e-07 $X=11381 $Y=20589 $D=636
M1990 1197 122 170 vdd hvtpfet l=6e-08 w=4.11e-07 $X=11381 $Y=22852 $D=636
M1991 1198 122 171 vdd hvtpfet l=6e-08 w=4.11e-07 $X=11381 $Y=27509 $D=636
M1992 b_pxbb_n<5> 164 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=11480 $Y=1941 $D=636
M1993 164 165 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=11480 $Y=5141 $D=636
M1994 165 106 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=11480 $Y=8691 $D=636
M1995 166 106 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=11480 $Y=41842 $D=636
M1996 167 166 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=11480 $Y=44992 $D=636
M1997 t_pxbb_n<5> 167 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=11480 $Y=46622 $D=636
M1998 47 162 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=11636 $Y=10167 $D=636
M1999 50 163 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=11636 $Y=40566 $D=636
M2000 vdd 33 1195 vdd hvtpfet l=6e-08 w=8.23e-07 $X=11651 $Y=15520 $D=636
M2001 vdd 33 1196 vdd hvtpfet l=6e-08 w=8.23e-07 $X=11651 $Y=20589 $D=636
M2002 vdd 33 1197 vdd hvtpfet l=6e-08 w=8.23e-07 $X=11651 $Y=22440 $D=636
M2003 vdd 33 1198 vdd hvtpfet l=6e-08 w=8.23e-07 $X=11651 $Y=27509 $D=636
M2004 172 142 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=11739 $Y=29948 $D=636
M2005 vdd 164 b_pxbb_n<5> vdd hvtpfet l=6e-08 w=2.57e-06 $X=11740 $Y=1941 $D=636
M2006 vdd 165 164 vdd hvtpfet l=6e-08 w=1e-06 $X=11740 $Y=5141 $D=636
M2007 vdd 106 165 vdd hvtpfet l=6e-08 w=6e-07 $X=11740 $Y=8691 $D=636
M2008 vdd 106 166 vdd hvtpfet l=6e-08 w=6e-07 $X=11740 $Y=41842 $D=636
M2009 vdd 166 167 vdd hvtpfet l=6e-08 w=1e-06 $X=11740 $Y=44992 $D=636
M2010 vdd 167 t_pxbb_n<5> vdd hvtpfet l=6e-08 w=2.57e-06 $X=11740 $Y=46622 $D=636
M2011 vdd tm<0> dbl_pd_n<0> vdd hvtpfet l=6e-08 w=4.28e-07 $X=11746 $Y=14263 $D=636
M2012 616 172 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=11933 $Y=35707 $D=636
M2013 dbl_pd_n<0> tm<0> vdd vdd hvtpfet l=6e-08 w=4.28e-07 $X=12006 $Y=14263 $D=636
M2014 179 173 vdd vdd hvtpfet l=6e-08 w=3e-07 $X=12086 $Y=33468 $D=636
M2015 vdd 174 2 vdd hvtpfet l=6e-08 w=4e-07 $X=12146 $Y=10167 $D=636
M2016 vdd 175 6 vdd hvtpfet l=6e-08 w=4e-07 $X=12146 $Y=40566 $D=636
M2017 177 168 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=12161 $Y=15321 $D=636
M2018 1199 43 168 vdd hvtpfet l=6e-08 w=2.74e-07 $X=12161 $Y=16069 $D=636
M2019 1200 43 169 vdd hvtpfet l=6e-08 w=2.74e-07 $X=12161 $Y=20589 $D=636
M2020 178 169 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=12161 $Y=21405 $D=636
M2021 137 170 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=12161 $Y=22241 $D=636
M2022 1201 43 170 vdd hvtpfet l=6e-08 w=2.74e-07 $X=12161 $Y=22989 $D=636
M2023 1202 43 171 vdd hvtpfet l=6e-08 w=2.74e-07 $X=12161 $Y=27509 $D=636
M2024 148 171 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=12161 $Y=28325 $D=636
M2025 vdd 172 616 vdd hvtpfet l=6e-08 w=1e-06 $X=12193 $Y=35707 $D=636
M2026 b_pxbb_n<6> 180 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=12250 $Y=1941 $D=636
M2027 180 181 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=12250 $Y=5141 $D=636
M2028 181 177 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=12250 $Y=8691 $D=636
M2029 182 177 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=12250 $Y=41842 $D=636
M2030 183 182 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=12250 $Y=44992 $D=636
M2031 t_pxbb_n<6> 183 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=12250 $Y=46622 $D=636
M2032 vdd tm<0> dbl_pd_n<0> vdd hvtpfet l=6e-08 w=4.28e-07 $X=12266 $Y=14263 $D=636
M2033 vdd 142 184 vdd hvtpfet l=6e-08 w=5e-07 $X=12339 $Y=29813 $D=636
M2034 vdd 168 177 vdd hvtpfet l=6e-08 w=2.06e-07 $X=12421 $Y=15321 $D=636
M2035 vdd 177 1199 vdd hvtpfet l=6e-08 w=2.74e-07 $X=12421 $Y=16069 $D=636
M2036 vdd 178 1200 vdd hvtpfet l=6e-08 w=2.74e-07 $X=12421 $Y=20589 $D=636
M2037 vdd 169 178 vdd hvtpfet l=6e-08 w=2.06e-07 $X=12421 $Y=21405 $D=636
M2038 vdd 170 137 vdd hvtpfet l=6e-08 w=2.06e-07 $X=12421 $Y=22241 $D=636
M2039 vdd 137 1201 vdd hvtpfet l=6e-08 w=2.74e-07 $X=12421 $Y=22989 $D=636
M2040 vdd 148 1202 vdd hvtpfet l=6e-08 w=2.74e-07 $X=12421 $Y=27509 $D=636
M2041 vdd 171 148 vdd hvtpfet l=6e-08 w=2.06e-07 $X=12421 $Y=28325 $D=636
M2042 616 172 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=12453 $Y=35707 $D=636
M2043 vdd 180 b_pxbb_n<6> vdd hvtpfet l=6e-08 w=2.57e-06 $X=12510 $Y=1941 $D=636
M2044 vdd 181 180 vdd hvtpfet l=6e-08 w=1e-06 $X=12510 $Y=5141 $D=636
M2045 vdd 177 181 vdd hvtpfet l=6e-08 w=6e-07 $X=12510 $Y=8691 $D=636
M2046 vdd 177 182 vdd hvtpfet l=6e-08 w=6e-07 $X=12510 $Y=41842 $D=636
M2047 vdd 182 183 vdd hvtpfet l=6e-08 w=1e-06 $X=12510 $Y=44992 $D=636
M2048 vdd 183 t_pxbb_n<6> vdd hvtpfet l=6e-08 w=2.57e-06 $X=12510 $Y=46622 $D=636
M2049 615 179 186 vdd hvtpfet l=6e-08 w=6e-07 $X=12596 $Y=33468 $D=636
M2050 191 184 vdd vdd hvtpfet l=2.5e-07 w=5e-07 $X=12599 $Y=29813 $D=636
M2051 vdd 185 174 vdd hvtpfet l=6e-08 w=4.11e-07 $X=12656 $Y=10156 $D=636
M2052 vdd 185 175 vdd hvtpfet l=6e-08 w=4.11e-07 $X=12656 $Y=40566 $D=636
M2053 620 186 616 vdd hvtpfet l=6e-08 w=1e-06 $X=12713 $Y=35707 $D=636
M2054 vdd 131 dbl_pd_n<2> vdd hvtpfet l=6e-08 w=4.28e-07 $X=12776 $Y=14263 $D=636
M2055 vdd 191 615 vdd hvtpfet l=6e-08 w=6e-07 $X=12856 $Y=33468 $D=636
M2056 174 dwlb<1> vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=12916 $Y=10156 $D=636
M2057 175 dwlb<0> vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=12916 $Y=40566 $D=636
M2058 187 192 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=12931 $Y=15321 $D=636
M2059 1203 187 vdd vdd hvtpfet l=6e-08 w=2.74e-07 $X=12931 $Y=16069 $D=636
M2060 1204 188 vdd vdd hvtpfet l=6e-08 w=2.74e-07 $X=12931 $Y=20589 $D=636
M2061 188 193 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=12931 $Y=21405 $D=636
M2062 189 194 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=12931 $Y=22241 $D=636
M2063 1205 189 vdd vdd hvtpfet l=6e-08 w=2.74e-07 $X=12931 $Y=22989 $D=636
M2064 1206 190 vdd vdd hvtpfet l=6e-08 w=2.74e-07 $X=12931 $Y=27509 $D=636
M2065 190 195 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=12931 $Y=28325 $D=636
M2066 616 186 620 vdd hvtpfet l=6e-08 w=1e-06 $X=12973 $Y=35707 $D=636
M2067 b_pxbb_n<7> 196 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=13020 $Y=1941 $D=636
M2068 196 197 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=13020 $Y=5141 $D=636
M2069 197 178 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=13020 $Y=8691 $D=636
M2070 198 178 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=13020 $Y=41842 $D=636
M2071 199 198 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=13020 $Y=44992 $D=636
M2072 t_pxbb_n<7> 199 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=13020 $Y=46622 $D=636
M2073 dbl_pd_n<2> 131 vdd vdd hvtpfet l=6e-08 w=4.28e-07 $X=13036 $Y=14263 $D=636
M2074 vdd 192 187 vdd hvtpfet l=6e-08 w=2.06e-07 $X=13191 $Y=15321 $D=636
M2075 192 43 1203 vdd hvtpfet l=6e-08 w=2.74e-07 $X=13191 $Y=16069 $D=636
M2076 193 43 1204 vdd hvtpfet l=6e-08 w=2.74e-07 $X=13191 $Y=20589 $D=636
M2077 vdd 193 188 vdd hvtpfet l=6e-08 w=2.06e-07 $X=13191 $Y=21405 $D=636
M2078 vdd 194 189 vdd hvtpfet l=6e-08 w=2.06e-07 $X=13191 $Y=22241 $D=636
M2079 194 43 1205 vdd hvtpfet l=6e-08 w=2.74e-07 $X=13191 $Y=22989 $D=636
M2080 195 43 1206 vdd hvtpfet l=6e-08 w=2.74e-07 $X=13191 $Y=27509 $D=636
M2081 vdd 195 190 vdd hvtpfet l=6e-08 w=2.06e-07 $X=13191 $Y=28325 $D=636
M2082 620 186 616 vdd hvtpfet l=6e-08 w=1e-06 $X=13233 $Y=35707 $D=636
M2083 vdd 196 b_pxbb_n<7> vdd hvtpfet l=6e-08 w=2.57e-06 $X=13280 $Y=1941 $D=636
M2084 vdd 197 196 vdd hvtpfet l=6e-08 w=1e-06 $X=13280 $Y=5141 $D=636
M2085 vdd 178 197 vdd hvtpfet l=6e-08 w=6e-07 $X=13280 $Y=8691 $D=636
M2086 vdd 178 198 vdd hvtpfet l=6e-08 w=6e-07 $X=13280 $Y=41842 $D=636
M2087 vdd 198 199 vdd hvtpfet l=6e-08 w=1e-06 $X=13280 $Y=44992 $D=636
M2088 vdd 199 t_pxbb_n<7> vdd hvtpfet l=6e-08 w=2.57e-06 $X=13280 $Y=46622 $D=636
M2089 vdd 131 dbl_pd_n<2> vdd hvtpfet l=6e-08 w=4.28e-07 $X=13296 $Y=14263 $D=636
M2090 vdd tm<7> 203 vdd hvtpfet l=6e-08 w=3e-07 $X=13432 $Y=33468 $D=636
M2091 vdd 191 202 vdd hvtpfet l=6e-08 w=5e-07 $X=13459 $Y=29813 $D=636
M2092 143 200 620 vdd hvtpfet l=6e-08 w=1e-06 $X=13493 $Y=35707 $D=636
M2093 1207 33 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=13701 $Y=15520 $D=636
M2094 1208 33 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=13701 $Y=20589 $D=636
M2095 1209 33 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=13701 $Y=22440 $D=636
M2096 1210 33 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=13701 $Y=27509 $D=636
M2097 211 202 vdd vdd hvtpfet l=2.5e-07 w=5e-07 $X=13719 $Y=29813 $D=636
M2098 620 200 143 vdd hvtpfet l=6e-08 w=1e-06 $X=13753 $Y=35707 $D=636
M2099 b_pxcb_n<0> 206 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=13790 $Y=1941 $D=636
M2100 206 207 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=13790 $Y=5141 $D=636
M2101 207 189 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=13790 $Y=8691 $D=636
M2102 208 189 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=13790 $Y=41842 $D=636
M2103 209 208 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=13790 $Y=44992 $D=636
M2104 t_pxcb_n<0> 209 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=13790 $Y=46622 $D=636
M2105 vdd 205 204 vdd hvtpfet l=6e-08 w=4.11e-07 $X=13936 $Y=14280 $D=636
M2106 623 203 200 vdd hvtpfet l=6e-08 w=6e-07 $X=13942 $Y=33468 $D=636
M2107 192 204 1207 vdd hvtpfet l=6e-08 w=4.11e-07 $X=13971 $Y=15932 $D=636
M2108 193 204 1208 vdd hvtpfet l=6e-08 w=4.11e-07 $X=13971 $Y=20589 $D=636
M2109 194 205 1209 vdd hvtpfet l=6e-08 w=4.11e-07 $X=13971 $Y=22852 $D=636
M2110 195 205 1210 vdd hvtpfet l=6e-08 w=4.11e-07 $X=13971 $Y=27509 $D=636
M2111 143 200 620 vdd hvtpfet l=6e-08 w=1e-06 $X=14013 $Y=35707 $D=636
M2112 vdd 206 b_pxcb_n<0> vdd hvtpfet l=6e-08 w=2.57e-06 $X=14050 $Y=1941 $D=636
M2113 vdd 207 206 vdd hvtpfet l=6e-08 w=1e-06 $X=14050 $Y=5141 $D=636
M2114 vdd 189 207 vdd hvtpfet l=6e-08 w=6e-07 $X=14050 $Y=8691 $D=636
M2115 vdd 189 208 vdd hvtpfet l=6e-08 w=6e-07 $X=14050 $Y=41842 $D=636
M2116 vdd 208 209 vdd hvtpfet l=6e-08 w=1e-06 $X=14050 $Y=44992 $D=636
M2117 vdd 209 t_pxcb_n<0> vdd hvtpfet l=6e-08 w=2.57e-06 $X=14050 $Y=46622 $D=636
M2118 vdd 211 623 vdd hvtpfet l=6e-08 w=6e-07 $X=14202 $Y=33468 $D=636
M2119 vdd dwlb<1> 216 vdd hvtpfet l=6e-08 w=4.11e-07 $X=14216 $Y=10156 $D=636
M2120 vdd dwlb<0> 217 vdd hvtpfet l=6e-08 w=4.11e-07 $X=14216 $Y=40566 $D=636
M2121 1211 210 192 vdd hvtpfet l=6e-08 w=4.11e-07 $X=14231 $Y=15932 $D=636
M2122 1212 210 193 vdd hvtpfet l=6e-08 w=4.11e-07 $X=14231 $Y=20589 $D=636
M2123 1213 210 194 vdd hvtpfet l=6e-08 w=4.11e-07 $X=14231 $Y=22852 $D=636
M2124 1214 210 195 vdd hvtpfet l=6e-08 w=4.11e-07 $X=14231 $Y=27509 $D=636
M2125 205 ab<12> vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=14446 $Y=14280 $D=636
M2126 216 212 vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=14476 $Y=10156 $D=636
M2127 217 212 vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=14476 $Y=40566 $D=636
M2128 vdd 33 1211 vdd hvtpfet l=6e-08 w=8.23e-07 $X=14501 $Y=15520 $D=636
M2129 vdd 33 1212 vdd hvtpfet l=6e-08 w=8.23e-07 $X=14501 $Y=20589 $D=636
M2130 vdd 33 1213 vdd hvtpfet l=6e-08 w=8.23e-07 $X=14501 $Y=22440 $D=636
M2131 vdd 33 1214 vdd hvtpfet l=6e-08 w=8.23e-07 $X=14501 $Y=27509 $D=636
M2132 b_pxcb_n<1> 218 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=14560 $Y=1941 $D=636
M2133 218 219 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=14560 $Y=5141 $D=636
M2134 219 190 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=14560 $Y=8691 $D=636
M2135 220 190 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=14560 $Y=41842 $D=636
M2136 221 220 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=14560 $Y=44992 $D=636
M2137 t_pxcb_n<1> 221 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=14560 $Y=46622 $D=636
M2138 vdd 123 624 vdd hvtpfet l=6e-08 w=1.2e-06 $X=14796 $Y=29148 $D=636
M2139 vdd 218 b_pxcb_n<1> vdd hvtpfet l=6e-08 w=2.57e-06 $X=14820 $Y=1941 $D=636
M2140 vdd 219 218 vdd hvtpfet l=6e-08 w=1e-06 $X=14820 $Y=5141 $D=636
M2141 vdd 190 219 vdd hvtpfet l=6e-08 w=6e-07 $X=14820 $Y=8691 $D=636
M2142 vdd 190 220 vdd hvtpfet l=6e-08 w=6e-07 $X=14820 $Y=41842 $D=636
M2143 vdd 220 221 vdd hvtpfet l=6e-08 w=1e-06 $X=14820 $Y=44992 $D=636
M2144 vdd 221 t_pxcb_n<1> vdd hvtpfet l=6e-08 w=2.57e-06 $X=14820 $Y=46622 $D=636
M2145 vdd 72 58 vdd hvtpfet l=6e-08 w=4e-07 $X=14872 $Y=35682 $D=636
M2146 48 216 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=14986 $Y=10167 $D=636
M2147 49 217 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=14986 $Y=40566 $D=636
M2148 1215 213 192 vdd hvtpfet l=6e-08 w=4.11e-07 $X=15011 $Y=15932 $D=636
M2149 1216 214 193 vdd hvtpfet l=6e-08 w=4.11e-07 $X=15011 $Y=20589 $D=636
M2150 1217 213 194 vdd hvtpfet l=6e-08 w=4.11e-07 $X=15011 $Y=22852 $D=636
M2151 1218 214 195 vdd hvtpfet l=6e-08 w=4.11e-07 $X=15011 $Y=27509 $D=636
M2152 33 43 vdd vdd hvtpfet l=6e-08 w=7e-07 $X=15056 $Y=29648 $D=636
M2153 vdd 33 1215 vdd hvtpfet l=6e-08 w=8.23e-07 $X=15281 $Y=15520 $D=636
M2154 vdd 33 1216 vdd hvtpfet l=6e-08 w=8.23e-07 $X=15281 $Y=20589 $D=636
M2155 vdd 33 1217 vdd hvtpfet l=6e-08 w=8.23e-07 $X=15281 $Y=22440 $D=636
M2156 vdd 33 1218 vdd hvtpfet l=6e-08 w=8.23e-07 $X=15281 $Y=27509 $D=636
M2157 vdd 43 33 vdd hvtpfet l=6e-08 w=7e-07 $X=15316 $Y=29648 $D=636
M2158 b_pxcb_n<2> 223 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=15330 $Y=1941 $D=636
M2159 223 224 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=15330 $Y=5141 $D=636
M2160 224 225 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=15330 $Y=8691 $D=636
M2161 226 225 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=15330 $Y=41842 $D=636
M2162 227 226 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=15330 $Y=44992 $D=636
M2163 t_pxcb_n<2> 227 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=15330 $Y=46622 $D=636
M2164 vdd 229 72 vdd hvtpfet l=6e-08 w=4e-07 $X=15382 $Y=35682 $D=636
M2165 vdd ab<11> 210 vdd hvtpfet l=6e-08 w=4.11e-07 $X=15456 $Y=14280 $D=636
M2166 1219 33 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=15541 $Y=15520 $D=636
M2167 1220 33 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=15541 $Y=20589 $D=636
M2168 1221 33 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=15541 $Y=22440 $D=636
M2169 1222 33 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=15541 $Y=27509 $D=636
M2170 33 43 vdd vdd hvtpfet l=6e-08 w=7e-07 $X=15576 $Y=29648 $D=636
M2171 vdd 223 b_pxcb_n<2> vdd hvtpfet l=6e-08 w=2.57e-06 $X=15590 $Y=1941 $D=636
M2172 vdd 224 223 vdd hvtpfet l=6e-08 w=1e-06 $X=15590 $Y=5141 $D=636
M2173 vdd 225 224 vdd hvtpfet l=6e-08 w=6e-07 $X=15590 $Y=8691 $D=636
M2174 vdd 225 226 vdd hvtpfet l=6e-08 w=6e-07 $X=15590 $Y=41842 $D=636
M2175 vdd 226 227 vdd hvtpfet l=6e-08 w=1e-06 $X=15590 $Y=44992 $D=636
M2176 vdd 227 t_pxcb_n<2> vdd hvtpfet l=6e-08 w=2.57e-06 $X=15590 $Y=46622 $D=636
M2177 vdd 228 231 vdd hvtpfet l=6e-08 w=3.2e-07 $X=15621 $Y=33942 $D=636
M2178 72 172 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=15642 $Y=35682 $D=636
M2179 240 210 vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=15716 $Y=14280 $D=636
M2180 249 213 1219 vdd hvtpfet l=6e-08 w=4.11e-07 $X=15811 $Y=15932 $D=636
M2181 250 214 1220 vdd hvtpfet l=6e-08 w=4.11e-07 $X=15811 $Y=20589 $D=636
M2182 251 213 1221 vdd hvtpfet l=6e-08 w=4.11e-07 $X=15811 $Y=22852 $D=636
M2183 252 214 1222 vdd hvtpfet l=6e-08 w=4.11e-07 $X=15811 $Y=27509 $D=636
M2184 vdd 43 33 vdd hvtpfet l=6e-08 w=7e-07 $X=15836 $Y=29648 $D=636
M2185 631 tm<0> vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=15880 $Y=40177 $D=636
M2186 632 123 vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=15881 $Y=33942 $D=636
M2187 vdd tm<3> 242 vdd hvtpfet l=7e-08 w=4.8e-07 $X=16057 $Y=10476 $D=636
M2188 b_pxcb_n<3> 235 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=16100 $Y=1941 $D=636
M2189 235 236 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=16100 $Y=5141 $D=636
M2190 236 237 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=16100 $Y=8691 $D=636
M2191 238 237 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=16100 $Y=41842 $D=636
M2192 239 238 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=16100 $Y=44992 $D=636
M2193 t_pxcb_n<3> 239 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=16100 $Y=46622 $D=636
M2194 228 231 632 vdd hvtpfet l=6e-08 w=3.2e-07 $X=16141 $Y=33942 $D=636
M2195 vdd 213 214 vdd hvtpfet l=6e-08 w=4.11e-07 $X=16316 $Y=14280 $D=636
M2196 1225 33 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=16321 $Y=15520 $D=636
M2197 1226 33 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=16321 $Y=20589 $D=636
M2198 1227 33 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=16321 $Y=22440 $D=636
M2199 1228 33 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=16321 $Y=27509 $D=636
M2200 1223 232 vdd vdd hvtpfet l=6e-08 w=4.8e-07 $X=16322 $Y=35753 $D=636
M2201 243 tm<4> vdd vdd hvtpfet l=7e-08 w=4.8e-07 $X=16327 $Y=10476 $D=636
M2202 642 123 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=16346 $Y=29274 $D=636
M2203 vdd 235 b_pxcb_n<3> vdd hvtpfet l=6e-08 w=2.57e-06 $X=16360 $Y=1941 $D=636
M2204 vdd 236 235 vdd hvtpfet l=6e-08 w=1e-06 $X=16360 $Y=5141 $D=636
M2205 vdd 237 236 vdd hvtpfet l=6e-08 w=6e-07 $X=16360 $Y=8691 $D=636
M2206 vdd 237 238 vdd hvtpfet l=6e-08 w=6e-07 $X=16360 $Y=41842 $D=636
M2207 vdd 238 239 vdd hvtpfet l=6e-08 w=1e-06 $X=16360 $Y=44992 $D=636
M2208 vdd 239 t_pxcb_n<3> vdd hvtpfet l=6e-08 w=2.57e-06 $X=16360 $Y=46622 $D=636
M2209 1224 131 228 vdd hvtpfet l=6e-08 w=4.8e-07 $X=16401 $Y=33942 $D=636
M2210 213 ab<10> vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=16576 $Y=14280 $D=636
M2211 229 172 1223 vdd hvtpfet l=6e-08 w=4.8e-07 $X=16582 $Y=35753 $D=636
M2212 249 240 1225 vdd hvtpfet l=6e-08 w=4.11e-07 $X=16591 $Y=15932 $D=636
M2213 250 240 1226 vdd hvtpfet l=6e-08 w=4.11e-07 $X=16591 $Y=20589 $D=636
M2214 251 240 1227 vdd hvtpfet l=6e-08 w=4.11e-07 $X=16591 $Y=22852 $D=636
M2215 252 240 1228 vdd hvtpfet l=6e-08 w=4.11e-07 $X=16591 $Y=27509 $D=636
M2216 vdd 123 642 vdd hvtpfet l=6e-08 w=6e-07 $X=16606 $Y=29274 $D=636
M2217 vdd 123 1224 vdd hvtpfet l=6e-08 w=4.8e-07 $X=16661 $Y=33942 $D=636
M2218 637 tm<6> vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=16680 $Y=40177 $D=636
M2219 639 244 229 vdd hvtpfet l=6e-08 w=3.2e-07 $X=16842 $Y=35913 $D=636
M2220 1229 243 643 vdd hvtpfet l=6e-08 w=4.8e-07 $X=16847 $Y=10476 $D=636
M2221 1230 204 249 vdd hvtpfet l=6e-08 w=4.11e-07 $X=16851 $Y=15932 $D=636
M2222 1231 204 250 vdd hvtpfet l=6e-08 w=4.11e-07 $X=16851 $Y=20589 $D=636
M2223 1232 205 251 vdd hvtpfet l=6e-08 w=4.11e-07 $X=16851 $Y=22852 $D=636
M2224 1233 205 252 vdd hvtpfet l=6e-08 w=4.11e-07 $X=16851 $Y=27509 $D=636
M2225 642 123 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=16866 $Y=29274 $D=636
M2226 b_pxcb_n<4> 245 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=16870 $Y=1941 $D=636
M2227 245 246 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=16870 $Y=5141 $D=636
M2228 246 187 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=16870 $Y=8691 $D=636
M2229 247 187 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=16870 $Y=41842 $D=636
M2230 248 247 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=16870 $Y=44992 $D=636
M2231 t_pxcb_n<4> 248 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=16870 $Y=46622 $D=636
M2232 vdd 142 639 vdd hvtpfet l=6e-08 w=3.2e-07 $X=17102 $Y=35913 $D=636
M2233 vdd 242 1229 vdd hvtpfet l=6e-08 w=4.8e-07 $X=17107 $Y=10476 $D=636
M2234 vdd 33 1230 vdd hvtpfet l=6e-08 w=8.23e-07 $X=17121 $Y=15520 $D=636
M2235 vdd 33 1231 vdd hvtpfet l=6e-08 w=8.23e-07 $X=17121 $Y=20589 $D=636
M2236 vdd 33 1232 vdd hvtpfet l=6e-08 w=8.23e-07 $X=17121 $Y=22440 $D=636
M2237 vdd 33 1233 vdd hvtpfet l=6e-08 w=8.23e-07 $X=17121 $Y=27509 $D=636
M2238 vdd 123 642 vdd hvtpfet l=6e-08 w=6e-07 $X=17126 $Y=29274 $D=636
M2239 vdd 245 b_pxcb_n<4> vdd hvtpfet l=6e-08 w=2.57e-06 $X=17130 $Y=1941 $D=636
M2240 vdd 246 245 vdd hvtpfet l=6e-08 w=1e-06 $X=17130 $Y=5141 $D=636
M2241 vdd 187 246 vdd hvtpfet l=6e-08 w=6e-07 $X=17130 $Y=8691 $D=636
M2242 vdd 187 247 vdd hvtpfet l=6e-08 w=6e-07 $X=17130 $Y=41842 $D=636
M2243 vdd 247 248 vdd hvtpfet l=6e-08 w=1e-06 $X=17130 $Y=44992 $D=636
M2244 vdd 248 t_pxcb_n<4> vdd hvtpfet l=6e-08 w=2.57e-06 $X=17130 $Y=46622 $D=636
M2245 244 229 vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=17362 $Y=35913 $D=636
M2246 1234 242 vdd vdd hvtpfet l=6e-08 w=4.8e-07 $X=17617 $Y=10476 $D=636
M2247 253 249 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=17631 $Y=15321 $D=636
M2248 1235 43 249 vdd hvtpfet l=6e-08 w=2.74e-07 $X=17631 $Y=16069 $D=636
M2249 1236 43 250 vdd hvtpfet l=6e-08 w=2.74e-07 $X=17631 $Y=20589 $D=636
M2250 254 250 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=17631 $Y=21405 $D=636
M2251 225 251 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=17631 $Y=22241 $D=636
M2252 1237 43 251 vdd hvtpfet l=6e-08 w=2.74e-07 $X=17631 $Y=22989 $D=636
M2253 1238 43 252 vdd hvtpfet l=6e-08 w=2.74e-07 $X=17631 $Y=27509 $D=636
M2254 237 252 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=17631 $Y=28325 $D=636
M2255 b_pxcb_n<5> 255 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=17640 $Y=1941 $D=636
M2256 255 256 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=17640 $Y=5141 $D=636
M2257 256 188 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=17640 $Y=8691 $D=636
M2258 257 188 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=17640 $Y=41842 $D=636
M2259 258 257 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=17640 $Y=44992 $D=636
M2260 t_pxcb_n<5> 258 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=17640 $Y=46622 $D=636
M2261 23 clkb vdd vdd hvtpfet l=6e-08 w=9e-07 $X=17646 $Y=29274 $D=636
M2262 647 tm<4> 1234 vdd hvtpfet l=6e-08 w=4.8e-07 $X=17877 $Y=10476 $D=636
M2263 vdd 249 253 vdd hvtpfet l=6e-08 w=2.06e-07 $X=17891 $Y=15321 $D=636
M2264 vdd 253 1235 vdd hvtpfet l=6e-08 w=2.74e-07 $X=17891 $Y=16069 $D=636
M2265 vdd 254 1236 vdd hvtpfet l=6e-08 w=2.74e-07 $X=17891 $Y=20589 $D=636
M2266 vdd 250 254 vdd hvtpfet l=6e-08 w=2.06e-07 $X=17891 $Y=21405 $D=636
M2267 vdd 251 225 vdd hvtpfet l=6e-08 w=2.06e-07 $X=17891 $Y=22241 $D=636
M2268 vdd 225 1237 vdd hvtpfet l=6e-08 w=2.74e-07 $X=17891 $Y=22989 $D=636
M2269 vdd 237 1238 vdd hvtpfet l=6e-08 w=2.74e-07 $X=17891 $Y=27509 $D=636
M2270 vdd 252 237 vdd hvtpfet l=6e-08 w=2.06e-07 $X=17891 $Y=28325 $D=636
M2271 vdd 255 b_pxcb_n<5> vdd hvtpfet l=6e-08 w=2.57e-06 $X=17900 $Y=1941 $D=636
M2272 vdd 256 255 vdd hvtpfet l=6e-08 w=1e-06 $X=17900 $Y=5141 $D=636
M2273 vdd 188 256 vdd hvtpfet l=6e-08 w=6e-07 $X=17900 $Y=8691 $D=636
M2274 vdd 188 257 vdd hvtpfet l=6e-08 w=6e-07 $X=17900 $Y=41842 $D=636
M2275 vdd 257 258 vdd hvtpfet l=6e-08 w=1e-06 $X=17900 $Y=44992 $D=636
M2276 vdd 258 t_pxcb_n<5> vdd hvtpfet l=6e-08 w=2.57e-06 $X=17900 $Y=46622 $D=636
M2277 vdd 260 273 vdd hvtpfet l=6e-08 w=4.11e-07 $X=18106 $Y=14280 $D=636
M2278 1239 wenb 232 vdd hvtpfet l=6e-08 w=8e-07 $X=18366 $Y=35907 $D=636
M2279 1240 tm<4> 648 vdd hvtpfet l=6e-08 w=4.8e-07 $X=18387 $Y=10476 $D=636
M2280 b_pxcb_n<6> 265 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=18410 $Y=1941 $D=636
M2281 265 266 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=18410 $Y=5141 $D=636
M2282 266 253 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=18410 $Y=8691 $D=636
M2283 267 253 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=18410 $Y=41842 $D=636
M2284 268 267 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=18410 $Y=44992 $D=636
M2285 t_pxcb_n<6> 268 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=18410 $Y=46622 $D=636
M2286 1241 ab<4> vdd vdd hvtpfet l=6e-08 w=4.8e-07 $X=18460 $Y=29394 $D=636
M2287 1242 wenb vdd vdd hvtpfet l=6e-08 w=4.8e-07 $X=18460 $Y=33942 $D=636
M2288 vdd tm<2> 173 vdd hvtpfet l=6e-08 w=4.11e-07 $X=18510 $Y=40177 $D=636
M2289 260 ab<1> vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=18616 $Y=14280 $D=636
M2290 vdd 264 1239 vdd hvtpfet l=6e-08 w=8e-07 $X=18626 $Y=35907 $D=636
M2291 1243 33 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=18641 $Y=15520 $D=636
M2292 1244 33 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=18641 $Y=20589 $D=636
M2293 1245 33 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=18641 $Y=22440 $D=636
M2294 1246 33 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=18641 $Y=27509 $D=636
M2295 vdd tm<3> 1240 vdd hvtpfet l=6e-08 w=4.8e-07 $X=18647 $Y=10476 $D=636
M2296 vdd 265 b_pxcb_n<6> vdd hvtpfet l=6e-08 w=2.57e-06 $X=18670 $Y=1941 $D=636
M2297 vdd 266 265 vdd hvtpfet l=6e-08 w=1e-06 $X=18670 $Y=5141 $D=636
M2298 vdd 253 266 vdd hvtpfet l=6e-08 w=6e-07 $X=18670 $Y=8691 $D=636
M2299 vdd 253 267 vdd hvtpfet l=6e-08 w=6e-07 $X=18670 $Y=41842 $D=636
M2300 vdd 267 268 vdd hvtpfet l=6e-08 w=1e-06 $X=18670 $Y=44992 $D=636
M2301 vdd 268 t_pxcb_n<6> vdd hvtpfet l=6e-08 w=2.57e-06 $X=18670 $Y=46622 $D=636
M2302 154 clkb 1241 vdd hvtpfet l=6e-08 w=4.8e-07 $X=18720 $Y=29394 $D=636
M2303 274 clkb 1242 vdd hvtpfet l=6e-08 w=4.8e-07 $X=18720 $Y=33942 $D=636
M2304 280 269 1243 vdd hvtpfet l=6e-08 w=4.11e-07 $X=18911 $Y=15932 $D=636
M2305 281 270 1244 vdd hvtpfet l=6e-08 w=4.11e-07 $X=18911 $Y=20589 $D=636
M2306 282 269 1245 vdd hvtpfet l=6e-08 w=4.11e-07 $X=18911 $Y=22852 $D=636
M2307 283 270 1246 vdd hvtpfet l=6e-08 w=4.11e-07 $X=18911 $Y=27509 $D=636
M2308 655 271 154 vdd hvtpfet l=6e-08 w=3.2e-07 $X=18980 $Y=29554 $D=636
M2309 656 272 274 vdd hvtpfet l=6e-08 w=3.2e-07 $X=18980 $Y=33942 $D=636
M2310 vdd 270 269 vdd hvtpfet l=6e-08 w=4.11e-07 $X=19126 $Y=14280 $D=636
M2311 1247 tm<3> vdd vdd hvtpfet l=6e-08 w=4.8e-07 $X=19157 $Y=10476 $D=636
M2312 1248 273 280 vdd hvtpfet l=6e-08 w=4.11e-07 $X=19171 $Y=15932 $D=636
M2313 1249 273 281 vdd hvtpfet l=6e-08 w=4.11e-07 $X=19171 $Y=20589 $D=636
M2314 1250 260 282 vdd hvtpfet l=6e-08 w=4.11e-07 $X=19171 $Y=22852 $D=636
M2315 1251 260 283 vdd hvtpfet l=6e-08 w=4.11e-07 $X=19171 $Y=27509 $D=636
M2316 b_pxcb_n<7> 275 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=19180 $Y=1941 $D=636
M2317 275 276 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=19180 $Y=5141 $D=636
M2318 276 254 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=19180 $Y=8691 $D=636
M2319 277 254 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=19180 $Y=41842 $D=636
M2320 278 277 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=19180 $Y=44992 $D=636
M2321 t_pxcb_n<7> 278 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=19180 $Y=46622 $D=636
M2322 vdd 23 655 vdd hvtpfet l=6e-08 w=3.2e-07 $X=19240 $Y=29554 $D=636
M2323 vdd 23 656 vdd hvtpfet l=6e-08 w=3.2e-07 $X=19240 $Y=33942 $D=636
M2324 659 243 1247 vdd hvtpfet l=6e-08 w=4.8e-07 $X=19417 $Y=10476 $D=636
M2325 vdd 275 b_pxcb_n<7> vdd hvtpfet l=6e-08 w=2.57e-06 $X=19440 $Y=1941 $D=636
M2326 vdd 276 275 vdd hvtpfet l=6e-08 w=1e-06 $X=19440 $Y=5141 $D=636
M2327 vdd 254 276 vdd hvtpfet l=6e-08 w=6e-07 $X=19440 $Y=8691 $D=636
M2328 vdd 254 277 vdd hvtpfet l=6e-08 w=6e-07 $X=19440 $Y=41842 $D=636
M2329 vdd 277 278 vdd hvtpfet l=6e-08 w=1e-06 $X=19440 $Y=44992 $D=636
M2330 vdd 278 t_pxcb_n<7> vdd hvtpfet l=6e-08 w=2.57e-06 $X=19440 $Y=46622 $D=636
M2331 vdd 33 1248 vdd hvtpfet l=6e-08 w=8.23e-07 $X=19441 $Y=15520 $D=636
M2332 vdd 33 1249 vdd hvtpfet l=6e-08 w=8.23e-07 $X=19441 $Y=20589 $D=636
M2333 vdd 33 1250 vdd hvtpfet l=6e-08 w=8.23e-07 $X=19441 $Y=22440 $D=636
M2334 vdd 33 1251 vdd hvtpfet l=6e-08 w=8.23e-07 $X=19441 $Y=27509 $D=636
M2335 271 154 vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=19500 $Y=29554 $D=636
M2336 272 274 vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=19500 $Y=33942 $D=636
M2337 270 ab<0> vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=19636 $Y=14280 $D=636
M2338 vdd 15 r_saeb_n vdd hvtpfet l=6e-08 w=1.43e-06 $X=19675 $Y=35277 $D=636
M2339 r_saeb_n 15 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=19935 $Y=35277 $D=636
M2340 212 280 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=19951 $Y=15321 $D=636
M2341 1252 43 280 vdd hvtpfet l=6e-08 w=2.74e-07 $X=19951 $Y=16069 $D=636
M2342 1253 43 281 vdd hvtpfet l=6e-08 w=2.74e-07 $X=19951 $Y=20589 $D=636
M2343 185 281 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=19951 $Y=21405 $D=636
M2344 155 282 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=19951 $Y=22241 $D=636
M2345 1254 43 282 vdd hvtpfet l=6e-08 w=2.74e-07 $X=19951 $Y=22989 $D=636
M2346 1255 43 283 vdd hvtpfet l=6e-08 w=2.74e-07 $X=19951 $Y=27509 $D=636
M2347 145 283 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=19951 $Y=28325 $D=636
M2348 vdd 11 rb_cb<0> vdd hvtpfet l=6e-08 w=1.43e-06 $X=20195 $Y=1506 $D=636
M2349 vdd 12 rb_cb<2> vdd hvtpfet l=6e-08 w=1.43e-06 $X=20195 $Y=3566 $D=636
M2350 vdd 13 rb_mb<0> vdd hvtpfet l=6e-08 w=1.43e-06 $X=20195 $Y=7966 $D=636
M2351 vdd 14 rb_mb<2> vdd hvtpfet l=6e-08 w=1.43e-06 $X=20195 $Y=10026 $D=636
M2352 vdd 15 r_saeb_n vdd hvtpfet l=6e-08 w=1.43e-06 $X=20195 $Y=35277 $D=636
M2353 vdd 16 rt_mb<2> vdd hvtpfet l=6e-08 w=1.43e-06 $X=20195 $Y=39677 $D=636
M2354 vdd 17 rt_mb<0> vdd hvtpfet l=6e-08 w=1.43e-06 $X=20195 $Y=41737 $D=636
M2355 vdd 18 rt_cb<2> vdd hvtpfet l=6e-08 w=1.43e-06 $X=20195 $Y=46137 $D=636
M2356 vdd 19 rt_cb<0> vdd hvtpfet l=6e-08 w=1.43e-06 $X=20195 $Y=48197 $D=636
M2357 vdd 280 212 vdd hvtpfet l=6e-08 w=2.06e-07 $X=20211 $Y=15321 $D=636
M2358 vdd 212 1252 vdd hvtpfet l=6e-08 w=2.74e-07 $X=20211 $Y=16069 $D=636
M2359 vdd 185 1253 vdd hvtpfet l=6e-08 w=2.74e-07 $X=20211 $Y=20589 $D=636
M2360 vdd 281 185 vdd hvtpfet l=6e-08 w=2.06e-07 $X=20211 $Y=21405 $D=636
M2361 vdd 282 155 vdd hvtpfet l=6e-08 w=2.06e-07 $X=20211 $Y=22241 $D=636
M2362 vdd 155 1254 vdd hvtpfet l=6e-08 w=2.74e-07 $X=20211 $Y=22989 $D=636
M2363 vdd 145 1255 vdd hvtpfet l=6e-08 w=2.74e-07 $X=20211 $Y=27509 $D=636
M2364 vdd 283 145 vdd hvtpfet l=6e-08 w=2.06e-07 $X=20211 $Y=28325 $D=636
M2365 rb_cb<0> 11 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=20455 $Y=1506 $D=636
M2366 rb_cb<2> 12 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=20455 $Y=3566 $D=636
M2367 rb_mb<0> 13 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=20455 $Y=7966 $D=636
M2368 rb_mb<2> 14 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=20455 $Y=10026 $D=636
M2369 r_saeb_n 15 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=20455 $Y=35277 $D=636
M2370 rt_mb<2> 16 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=20455 $Y=39677 $D=636
M2371 rt_mb<0> 17 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=20455 $Y=41737 $D=636
M2372 rt_cb<2> 18 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=20455 $Y=46137 $D=636
M2373 rt_cb<0> 19 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=20455 $Y=48197 $D=636
M2374 vdd 11 rb_cb<0> vdd hvtpfet l=6e-08 w=1.43e-06 $X=20715 $Y=1506 $D=636
M2375 vdd 12 rb_cb<2> vdd hvtpfet l=6e-08 w=1.43e-06 $X=20715 $Y=3566 $D=636
M2376 vdd 13 rb_mb<0> vdd hvtpfet l=6e-08 w=1.43e-06 $X=20715 $Y=7966 $D=636
M2377 vdd 14 rb_mb<2> vdd hvtpfet l=6e-08 w=1.43e-06 $X=20715 $Y=10026 $D=636
M2378 vdd 15 r_saeb_n vdd hvtpfet l=6e-08 w=1.43e-06 $X=20715 $Y=35277 $D=636
M2379 vdd 16 rt_mb<2> vdd hvtpfet l=6e-08 w=1.43e-06 $X=20715 $Y=39677 $D=636
M2380 vdd 17 rt_mb<0> vdd hvtpfet l=6e-08 w=1.43e-06 $X=20715 $Y=41737 $D=636
M2381 vdd 18 rt_cb<2> vdd hvtpfet l=6e-08 w=1.43e-06 $X=20715 $Y=46137 $D=636
M2382 vdd 19 rt_cb<0> vdd hvtpfet l=6e-08 w=1.43e-06 $X=20715 $Y=48197 $D=636
M2383 10 274 vdd vdd hvtpfet l=6e-08 w=1.2e-06 $X=20725 $Y=32684 $D=636
M2384 rb_cb<1> 34 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=20975 $Y=1506 $D=636
M2385 rb_cb<3> 35 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=20975 $Y=3566 $D=636
M2386 rb_mb<1> 36 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=20975 $Y=7966 $D=636
M2387 rb_mb<3> 37 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=20975 $Y=10026 $D=636
M2388 r_clk_dqb 8 vdd vdd hvtpfet l=6e-08 w=2.1e-06 $X=20975 $Y=23696 $D=636
M2389 r_clk_dqb_n 9 vdd vdd hvtpfet l=6e-08 w=2.1e-06 $X=20975 $Y=26512 $D=636
M2390 r_sa_preb_n 51 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=20975 $Y=35277 $D=636
M2391 rt_mb<3> 39 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=20975 $Y=39677 $D=636
M2392 rt_mb<1> 40 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=20975 $Y=41737 $D=636
M2393 rt_cb<3> 41 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=20975 $Y=46137 $D=636
M2394 rt_cb<1> 42 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=20975 $Y=48197 $D=636
M2395 vdd 34 rb_cb<1> vdd hvtpfet l=6e-08 w=1.43e-06 $X=21235 $Y=1506 $D=636
M2396 vdd 35 rb_cb<3> vdd hvtpfet l=6e-08 w=1.43e-06 $X=21235 $Y=3566 $D=636
M2397 vdd 36 rb_mb<1> vdd hvtpfet l=6e-08 w=1.43e-06 $X=21235 $Y=7966 $D=636
M2398 vdd 37 rb_mb<3> vdd hvtpfet l=6e-08 w=1.43e-06 $X=21235 $Y=10026 $D=636
M2399 rb_tm_preb_n 20 vdd vdd hvtpfet l=6e-08 w=2.145e-06 $X=21235 $Y=14887 $D=636
M2400 rt_tm_preb_n 21 vdd vdd hvtpfet l=6e-08 w=2.145e-06 $X=21235 $Y=17659 $D=636
M2401 vdd 8 r_clk_dqb vdd hvtpfet l=6e-08 w=2.1e-06 $X=21235 $Y=23696 $D=636
M2402 vdd 9 r_clk_dqb_n vdd hvtpfet l=6e-08 w=2.1e-06 $X=21235 $Y=26512 $D=636
M2403 r_lweb 10 vdd vdd hvtpfet l=6e-08 w=2.145e-06 $X=21235 $Y=32504 $D=636
M2404 vdd 51 r_sa_preb_n vdd hvtpfet l=6e-08 w=1.43e-06 $X=21235 $Y=35277 $D=636
M2405 vdd 39 rt_mb<3> vdd hvtpfet l=6e-08 w=1.43e-06 $X=21235 $Y=39677 $D=636
M2406 vdd 40 rt_mb<1> vdd hvtpfet l=6e-08 w=1.43e-06 $X=21235 $Y=41737 $D=636
M2407 vdd 41 rt_cb<3> vdd hvtpfet l=6e-08 w=1.43e-06 $X=21235 $Y=46137 $D=636
M2408 vdd 42 rt_cb<1> vdd hvtpfet l=6e-08 w=1.43e-06 $X=21235 $Y=48197 $D=636
M2409 rb_cb<1> 34 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=21495 $Y=1506 $D=636
M2410 rb_cb<3> 35 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=21495 $Y=3566 $D=636
M2411 rb_mb<1> 36 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=21495 $Y=7966 $D=636
M2412 rb_mb<3> 37 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=21495 $Y=10026 $D=636
M2413 vdd 20 rb_tm_preb_n vdd hvtpfet l=6e-08 w=2.145e-06 $X=21495 $Y=14887 $D=636
M2414 vdd 21 rt_tm_preb_n vdd hvtpfet l=6e-08 w=2.145e-06 $X=21495 $Y=17659 $D=636
M2415 r_clk_dqb 8 vdd vdd hvtpfet l=6e-08 w=2.1e-06 $X=21495 $Y=23696 $D=636
M2416 r_clk_dqb_n 9 vdd vdd hvtpfet l=6e-08 w=2.1e-06 $X=21495 $Y=26512 $D=636
M2417 vdd 10 r_lweb vdd hvtpfet l=6e-08 w=2.145e-06 $X=21495 $Y=32504 $D=636
M2418 r_sa_preb_n 51 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=21495 $Y=35277 $D=636
M2419 rt_mb<3> 39 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=21495 $Y=39677 $D=636
M2420 rt_mb<1> 40 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=21495 $Y=41737 $D=636
M2421 rt_cb<3> 41 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=21495 $Y=46137 $D=636
M2422 rt_cb<1> 42 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=21495 $Y=48197 $D=636
M2423 vdd 289 lb_ca<1> vdd hvtpfet l=6e-08 w=1.43e-06 $X=22005 $Y=1506 $D=636
M2424 vdd 290 lb_ca<3> vdd hvtpfet l=6e-08 w=1.43e-06 $X=22005 $Y=3566 $D=636
M2425 vdd 291 lb_ma<1> vdd hvtpfet l=6e-08 w=1.43e-06 $X=22005 $Y=7966 $D=636
M2426 vdd 292 lb_ma<3> vdd hvtpfet l=6e-08 w=1.43e-06 $X=22005 $Y=10026 $D=636
M2427 lb_tm_prea_n 285 vdd vdd hvtpfet l=6e-08 w=2.145e-06 $X=22005 $Y=14887 $D=636
M2428 lt_tm_prea_n 286 vdd vdd hvtpfet l=6e-08 w=2.145e-06 $X=22005 $Y=17659 $D=636
M2429 vdd 287 l_clk_dqa vdd hvtpfet l=6e-08 w=2.1e-06 $X=22005 $Y=23696 $D=636
M2430 vdd 288 l_clk_dqa_n vdd hvtpfet l=6e-08 w=2.1e-06 $X=22005 $Y=26512 $D=636
M2431 l_lwea 284 vdd vdd hvtpfet l=6e-08 w=2.145e-06 $X=22005 $Y=32504 $D=636
M2432 vdd 293 l_sa_prea_n vdd hvtpfet l=6e-08 w=1.43e-06 $X=22005 $Y=35277 $D=636
M2433 vdd 294 lt_ma<3> vdd hvtpfet l=6e-08 w=1.43e-06 $X=22005 $Y=39677 $D=636
M2434 vdd 295 lt_ma<1> vdd hvtpfet l=6e-08 w=1.43e-06 $X=22005 $Y=41737 $D=636
M2435 vdd 296 lt_ca<3> vdd hvtpfet l=6e-08 w=1.43e-06 $X=22005 $Y=46137 $D=636
M2436 vdd 297 lt_ca<1> vdd hvtpfet l=6e-08 w=1.43e-06 $X=22005 $Y=48197 $D=636
M2437 lb_ca<1> 289 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=22265 $Y=1506 $D=636
M2438 lb_ca<3> 290 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=22265 $Y=3566 $D=636
M2439 lb_ma<1> 291 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=22265 $Y=7966 $D=636
M2440 lb_ma<3> 292 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=22265 $Y=10026 $D=636
M2441 vdd 285 lb_tm_prea_n vdd hvtpfet l=6e-08 w=2.145e-06 $X=22265 $Y=14887 $D=636
M2442 vdd 286 lt_tm_prea_n vdd hvtpfet l=6e-08 w=2.145e-06 $X=22265 $Y=17659 $D=636
M2443 l_clk_dqa 287 vdd vdd hvtpfet l=6e-08 w=2.1e-06 $X=22265 $Y=23696 $D=636
M2444 l_clk_dqa_n 288 vdd vdd hvtpfet l=6e-08 w=2.1e-06 $X=22265 $Y=26512 $D=636
M2445 vdd 284 l_lwea vdd hvtpfet l=6e-08 w=2.145e-06 $X=22265 $Y=32504 $D=636
M2446 l_sa_prea_n 293 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=22265 $Y=35277 $D=636
M2447 lt_ma<3> 294 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=22265 $Y=39677 $D=636
M2448 lt_ma<1> 295 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=22265 $Y=41737 $D=636
M2449 lt_ca<3> 296 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=22265 $Y=46137 $D=636
M2450 lt_ca<1> 297 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=22265 $Y=48197 $D=636
M2451 vdd 289 lb_ca<1> vdd hvtpfet l=6e-08 w=1.43e-06 $X=22525 $Y=1506 $D=636
M2452 vdd 290 lb_ca<3> vdd hvtpfet l=6e-08 w=1.43e-06 $X=22525 $Y=3566 $D=636
M2453 vdd 291 lb_ma<1> vdd hvtpfet l=6e-08 w=1.43e-06 $X=22525 $Y=7966 $D=636
M2454 vdd 292 lb_ma<3> vdd hvtpfet l=6e-08 w=1.43e-06 $X=22525 $Y=10026 $D=636
M2455 vdd 287 l_clk_dqa vdd hvtpfet l=6e-08 w=2.1e-06 $X=22525 $Y=23696 $D=636
M2456 vdd 288 l_clk_dqa_n vdd hvtpfet l=6e-08 w=2.1e-06 $X=22525 $Y=26512 $D=636
M2457 vdd 293 l_sa_prea_n vdd hvtpfet l=6e-08 w=1.43e-06 $X=22525 $Y=35277 $D=636
M2458 vdd 294 lt_ma<3> vdd hvtpfet l=6e-08 w=1.43e-06 $X=22525 $Y=39677 $D=636
M2459 vdd 295 lt_ma<1> vdd hvtpfet l=6e-08 w=1.43e-06 $X=22525 $Y=41737 $D=636
M2460 vdd 296 lt_ca<3> vdd hvtpfet l=6e-08 w=1.43e-06 $X=22525 $Y=46137 $D=636
M2461 vdd 297 lt_ca<1> vdd hvtpfet l=6e-08 w=1.43e-06 $X=22525 $Y=48197 $D=636
M2462 vdd 298 284 vdd hvtpfet l=6e-08 w=1.2e-06 $X=22775 $Y=32684 $D=636
M2463 lb_ca<0> 299 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=22785 $Y=1506 $D=636
M2464 lb_ca<2> 300 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=22785 $Y=3566 $D=636
M2465 lb_ma<0> 301 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=22785 $Y=7966 $D=636
M2466 lb_ma<2> 302 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=22785 $Y=10026 $D=636
M2467 l_saea_n 303 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=22785 $Y=35277 $D=636
M2468 lt_ma<2> 304 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=22785 $Y=39677 $D=636
M2469 lt_ma<0> 305 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=22785 $Y=41737 $D=636
M2470 lt_ca<2> 306 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=22785 $Y=46137 $D=636
M2471 lt_ca<0> 307 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=22785 $Y=48197 $D=636
M2472 vdd 299 lb_ca<0> vdd hvtpfet l=6e-08 w=1.43e-06 $X=23045 $Y=1506 $D=636
M2473 vdd 300 lb_ca<2> vdd hvtpfet l=6e-08 w=1.43e-06 $X=23045 $Y=3566 $D=636
M2474 vdd 301 lb_ma<0> vdd hvtpfet l=6e-08 w=1.43e-06 $X=23045 $Y=7966 $D=636
M2475 vdd 302 lb_ma<2> vdd hvtpfet l=6e-08 w=1.43e-06 $X=23045 $Y=10026 $D=636
M2476 vdd 303 l_saea_n vdd hvtpfet l=6e-08 w=1.43e-06 $X=23045 $Y=35277 $D=636
M2477 vdd 304 lt_ma<2> vdd hvtpfet l=6e-08 w=1.43e-06 $X=23045 $Y=39677 $D=636
M2478 vdd 305 lt_ma<0> vdd hvtpfet l=6e-08 w=1.43e-06 $X=23045 $Y=41737 $D=636
M2479 vdd 306 lt_ca<2> vdd hvtpfet l=6e-08 w=1.43e-06 $X=23045 $Y=46137 $D=636
M2480 vdd 307 lt_ca<0> vdd hvtpfet l=6e-08 w=1.43e-06 $X=23045 $Y=48197 $D=636
M2481 308 312 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=23289 $Y=15321 $D=636
M2482 1256 308 vdd vdd hvtpfet l=6e-08 w=2.74e-07 $X=23289 $Y=16069 $D=636
M2483 1257 309 vdd vdd hvtpfet l=6e-08 w=2.74e-07 $X=23289 $Y=20589 $D=636
M2484 309 313 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=23289 $Y=21405 $D=636
M2485 310 314 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=23289 $Y=22241 $D=636
M2486 1258 310 vdd vdd hvtpfet l=6e-08 w=2.74e-07 $X=23289 $Y=22989 $D=636
M2487 1259 311 vdd vdd hvtpfet l=6e-08 w=2.74e-07 $X=23289 $Y=27509 $D=636
M2488 311 315 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=23289 $Y=28325 $D=636
M2489 lb_ca<0> 299 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=23305 $Y=1506 $D=636
M2490 lb_ca<2> 300 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=23305 $Y=3566 $D=636
M2491 lb_ma<0> 301 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=23305 $Y=7966 $D=636
M2492 lb_ma<2> 302 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=23305 $Y=10026 $D=636
M2493 l_saea_n 303 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=23305 $Y=35277 $D=636
M2494 lt_ma<2> 304 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=23305 $Y=39677 $D=636
M2495 lt_ma<0> 305 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=23305 $Y=41737 $D=636
M2496 lt_ca<2> 306 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=23305 $Y=46137 $D=636
M2497 lt_ca<0> 307 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=23305 $Y=48197 $D=636
M2498 vdd 312 308 vdd hvtpfet l=6e-08 w=2.06e-07 $X=23549 $Y=15321 $D=636
M2499 312 323 1256 vdd hvtpfet l=6e-08 w=2.74e-07 $X=23549 $Y=16069 $D=636
M2500 313 323 1257 vdd hvtpfet l=6e-08 w=2.74e-07 $X=23549 $Y=20589 $D=636
M2501 vdd 313 309 vdd hvtpfet l=6e-08 w=2.06e-07 $X=23549 $Y=21405 $D=636
M2502 vdd 314 310 vdd hvtpfet l=6e-08 w=2.06e-07 $X=23549 $Y=22241 $D=636
M2503 314 323 1258 vdd hvtpfet l=6e-08 w=2.74e-07 $X=23549 $Y=22989 $D=636
M2504 315 323 1259 vdd hvtpfet l=6e-08 w=2.74e-07 $X=23549 $Y=27509 $D=636
M2505 vdd 315 311 vdd hvtpfet l=6e-08 w=2.06e-07 $X=23549 $Y=28325 $D=636
M2506 vdd 303 l_saea_n vdd hvtpfet l=6e-08 w=1.43e-06 $X=23565 $Y=35277 $D=636
M2507 l_saea_n 303 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=23825 $Y=35277 $D=636
M2508 vdd aa<0> 327 vdd hvtpfet l=6e-08 w=4.11e-07 $X=23864 $Y=14280 $D=636
M2509 vdd 324 331 vdd hvtpfet l=6e-08 w=3.2e-07 $X=24000 $Y=29554 $D=636
M2510 vdd 298 332 vdd hvtpfet l=6e-08 w=3.2e-07 $X=24000 $Y=33942 $D=636
M2511 1261 317 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=24059 $Y=15520 $D=636
M2512 1262 317 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=24059 $Y=20589 $D=636
M2513 1263 317 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=24059 $Y=22440 $D=636
M2514 1264 317 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=24059 $Y=27509 $D=636
M2515 b_pxca_n<7> 318 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=24060 $Y=1941 $D=636
M2516 318 319 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=24060 $Y=5141 $D=636
M2517 319 320 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=24060 $Y=8691 $D=636
M2518 321 320 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=24060 $Y=41842 $D=636
M2519 322 321 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=24060 $Y=44992 $D=636
M2520 t_pxca_n<7> 322 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=24060 $Y=46622 $D=636
M2521 1260 325 709 vdd hvtpfet l=6e-08 w=4.8e-07 $X=24083 $Y=10476 $D=636
M2522 712 340 vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=24260 $Y=29554 $D=636
M2523 713 340 vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=24260 $Y=33942 $D=636
M2524 vdd 318 b_pxca_n<7> vdd hvtpfet l=6e-08 w=2.57e-06 $X=24320 $Y=1941 $D=636
M2525 vdd 319 318 vdd hvtpfet l=6e-08 w=1e-06 $X=24320 $Y=5141 $D=636
M2526 vdd 320 319 vdd hvtpfet l=6e-08 w=6e-07 $X=24320 $Y=8691 $D=636
M2527 vdd 320 321 vdd hvtpfet l=6e-08 w=6e-07 $X=24320 $Y=41842 $D=636
M2528 vdd 321 322 vdd hvtpfet l=6e-08 w=1e-06 $X=24320 $Y=44992 $D=636
M2529 vdd 322 t_pxca_n<7> vdd hvtpfet l=6e-08 w=2.57e-06 $X=24320 $Y=46622 $D=636
M2530 312 328 1261 vdd hvtpfet l=6e-08 w=4.11e-07 $X=24329 $Y=15932 $D=636
M2531 313 328 1262 vdd hvtpfet l=6e-08 w=4.11e-07 $X=24329 $Y=20589 $D=636
M2532 314 329 1263 vdd hvtpfet l=6e-08 w=4.11e-07 $X=24329 $Y=22852 $D=636
M2533 315 329 1264 vdd hvtpfet l=6e-08 w=4.11e-07 $X=24329 $Y=27509 $D=636
M2534 vdd tm<8> 1260 vdd hvtpfet l=6e-08 w=4.8e-07 $X=24343 $Y=10476 $D=636
M2535 334 327 vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=24374 $Y=14280 $D=636
M2536 vdd tm<5> 264 vdd hvtpfet l=6e-08 w=4.11e-07 $X=24518 $Y=40177 $D=636
M2537 324 331 712 vdd hvtpfet l=6e-08 w=3.2e-07 $X=24520 $Y=29554 $D=636
M2538 298 332 713 vdd hvtpfet l=6e-08 w=3.2e-07 $X=24520 $Y=33942 $D=636
M2539 1265 334 312 vdd hvtpfet l=6e-08 w=4.11e-07 $X=24589 $Y=15932 $D=636
M2540 1266 327 313 vdd hvtpfet l=6e-08 w=4.11e-07 $X=24589 $Y=20589 $D=636
M2541 1267 334 314 vdd hvtpfet l=6e-08 w=4.11e-07 $X=24589 $Y=22852 $D=636
M2542 1268 327 315 vdd hvtpfet l=6e-08 w=4.11e-07 $X=24589 $Y=27509 $D=636
M2543 1269 clka 324 vdd hvtpfet l=6e-08 w=4.8e-07 $X=24780 $Y=29394 $D=636
M2544 1270 clka 298 vdd hvtpfet l=6e-08 w=4.8e-07 $X=24780 $Y=33942 $D=636
M2545 b_pxca_n<6> 335 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=24830 $Y=1941 $D=636
M2546 335 336 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=24830 $Y=5141 $D=636
M2547 336 337 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=24830 $Y=8691 $D=636
M2548 338 337 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=24830 $Y=41842 $D=636
M2549 339 338 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=24830 $Y=44992 $D=636
M2550 t_pxca_n<6> 339 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=24830 $Y=46622 $D=636
M2551 1271 tm<8> vdd vdd hvtpfet l=6e-08 w=4.8e-07 $X=24853 $Y=10476 $D=636
M2552 vdd 317 1265 vdd hvtpfet l=6e-08 w=8.23e-07 $X=24859 $Y=15520 $D=636
M2553 vdd 317 1266 vdd hvtpfet l=6e-08 w=8.23e-07 $X=24859 $Y=20589 $D=636
M2554 vdd 317 1267 vdd hvtpfet l=6e-08 w=8.23e-07 $X=24859 $Y=22440 $D=636
M2555 vdd 317 1268 vdd hvtpfet l=6e-08 w=8.23e-07 $X=24859 $Y=27509 $D=636
M2556 1272 264 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=24874 $Y=35907 $D=636
M2557 vdd aa<1> 329 vdd hvtpfet l=6e-08 w=4.11e-07 $X=24884 $Y=14280 $D=636
M2558 vdd aa<4> 1269 vdd hvtpfet l=6e-08 w=4.8e-07 $X=25040 $Y=29394 $D=636
M2559 vdd wena 1270 vdd hvtpfet l=6e-08 w=4.8e-07 $X=25040 $Y=33942 $D=636
M2560 vdd 335 b_pxca_n<6> vdd hvtpfet l=6e-08 w=2.57e-06 $X=25090 $Y=1941 $D=636
M2561 vdd 336 335 vdd hvtpfet l=6e-08 w=1e-06 $X=25090 $Y=5141 $D=636
M2562 vdd 337 336 vdd hvtpfet l=6e-08 w=6e-07 $X=25090 $Y=8691 $D=636
M2563 vdd 337 338 vdd hvtpfet l=6e-08 w=6e-07 $X=25090 $Y=41842 $D=636
M2564 vdd 338 339 vdd hvtpfet l=6e-08 w=1e-06 $X=25090 $Y=44992 $D=636
M2565 vdd 339 t_pxca_n<6> vdd hvtpfet l=6e-08 w=2.57e-06 $X=25090 $Y=46622 $D=636
M2566 718 tm<9> 1271 vdd hvtpfet l=6e-08 w=4.8e-07 $X=25113 $Y=10476 $D=636
M2567 376 wena 1272 vdd hvtpfet l=6e-08 w=8e-07 $X=25134 $Y=35907 $D=636
M2568 328 329 vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=25394 $Y=14280 $D=636
M2569 b_pxca_n<5> 345 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=25600 $Y=1941 $D=636
M2570 345 346 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=25600 $Y=5141 $D=636
M2571 346 347 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=25600 $Y=8691 $D=636
M2572 348 347 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=25600 $Y=41842 $D=636
M2573 349 348 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=25600 $Y=44992 $D=636
M2574 t_pxca_n<5> 349 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=25600 $Y=46622 $D=636
M2575 337 352 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=25609 $Y=15321 $D=636
M2576 1273 337 vdd vdd hvtpfet l=6e-08 w=2.74e-07 $X=25609 $Y=16069 $D=636
M2577 1274 320 vdd vdd hvtpfet l=6e-08 w=2.74e-07 $X=25609 $Y=20589 $D=636
M2578 320 353 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=25609 $Y=21405 $D=636
M2579 350 354 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=25609 $Y=22241 $D=636
M2580 1275 350 vdd vdd hvtpfet l=6e-08 w=2.74e-07 $X=25609 $Y=22989 $D=636
M2581 1276 351 vdd vdd hvtpfet l=6e-08 w=2.74e-07 $X=25609 $Y=27509 $D=636
M2582 351 355 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=25609 $Y=28325 $D=636
M2583 1277 tm<9> 721 vdd hvtpfet l=6e-08 w=4.8e-07 $X=25623 $Y=10476 $D=636
M2584 vdd clka 340 vdd hvtpfet l=6e-08 w=9e-07 $X=25854 $Y=29274 $D=636
M2585 vdd 345 b_pxca_n<5> vdd hvtpfet l=6e-08 w=2.57e-06 $X=25860 $Y=1941 $D=636
M2586 vdd 346 345 vdd hvtpfet l=6e-08 w=1e-06 $X=25860 $Y=5141 $D=636
M2587 vdd 347 346 vdd hvtpfet l=6e-08 w=6e-07 $X=25860 $Y=8691 $D=636
M2588 vdd 347 348 vdd hvtpfet l=6e-08 w=6e-07 $X=25860 $Y=41842 $D=636
M2589 vdd 348 349 vdd hvtpfet l=6e-08 w=1e-06 $X=25860 $Y=44992 $D=636
M2590 vdd 349 t_pxca_n<5> vdd hvtpfet l=6e-08 w=2.57e-06 $X=25860 $Y=46622 $D=636
M2591 vdd 352 337 vdd hvtpfet l=6e-08 w=2.06e-07 $X=25869 $Y=15321 $D=636
M2592 352 323 1273 vdd hvtpfet l=6e-08 w=2.74e-07 $X=25869 $Y=16069 $D=636
M2593 353 323 1274 vdd hvtpfet l=6e-08 w=2.74e-07 $X=25869 $Y=20589 $D=636
M2594 vdd 353 320 vdd hvtpfet l=6e-08 w=2.06e-07 $X=25869 $Y=21405 $D=636
M2595 vdd 354 350 vdd hvtpfet l=6e-08 w=2.06e-07 $X=25869 $Y=22241 $D=636
M2596 354 323 1275 vdd hvtpfet l=6e-08 w=2.74e-07 $X=25869 $Y=22989 $D=636
M2597 355 323 1276 vdd hvtpfet l=6e-08 w=2.74e-07 $X=25869 $Y=27509 $D=636
M2598 vdd 355 351 vdd hvtpfet l=6e-08 w=2.06e-07 $X=25869 $Y=28325 $D=636
M2599 vdd 366 1277 vdd hvtpfet l=6e-08 w=4.8e-07 $X=25883 $Y=10476 $D=636
M2600 vdd 356 363 vdd hvtpfet l=6e-08 w=3.2e-07 $X=26138 $Y=35913 $D=636
M2601 b_pxca_n<4> 357 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=26370 $Y=1941 $D=636
M2602 357 358 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=26370 $Y=5141 $D=636
M2603 358 359 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=26370 $Y=8691 $D=636
M2604 360 359 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=26370 $Y=41842 $D=636
M2605 361 360 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=26370 $Y=44992 $D=636
M2606 t_pxca_n<4> 361 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=26370 $Y=46622 $D=636
M2607 729 123 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=26374 $Y=29274 $D=636
M2608 1279 317 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=26379 $Y=15520 $D=636
M2609 1280 317 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=26379 $Y=20589 $D=636
M2610 1281 317 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=26379 $Y=22440 $D=636
M2611 1282 317 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=26379 $Y=27509 $D=636
M2612 1278 366 vdd vdd hvtpfet l=6e-08 w=4.8e-07 $X=26393 $Y=10476 $D=636
M2613 725 368 vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=26398 $Y=35913 $D=636
M2614 vdd 357 b_pxca_n<4> vdd hvtpfet l=6e-08 w=2.57e-06 $X=26630 $Y=1941 $D=636
M2615 vdd 358 357 vdd hvtpfet l=6e-08 w=1e-06 $X=26630 $Y=5141 $D=636
M2616 vdd 359 358 vdd hvtpfet l=6e-08 w=6e-07 $X=26630 $Y=8691 $D=636
M2617 vdd 359 360 vdd hvtpfet l=6e-08 w=6e-07 $X=26630 $Y=41842 $D=636
M2618 vdd 360 361 vdd hvtpfet l=6e-08 w=1e-06 $X=26630 $Y=44992 $D=636
M2619 vdd 361 t_pxca_n<4> vdd hvtpfet l=6e-08 w=2.57e-06 $X=26630 $Y=46622 $D=636
M2620 vdd 123 729 vdd hvtpfet l=6e-08 w=6e-07 $X=26634 $Y=29274 $D=636
M2621 352 364 1279 vdd hvtpfet l=6e-08 w=4.11e-07 $X=26649 $Y=15932 $D=636
M2622 353 364 1280 vdd hvtpfet l=6e-08 w=4.11e-07 $X=26649 $Y=20589 $D=636
M2623 354 365 1281 vdd hvtpfet l=6e-08 w=4.11e-07 $X=26649 $Y=22852 $D=636
M2624 355 365 1282 vdd hvtpfet l=6e-08 w=4.11e-07 $X=26649 $Y=27509 $D=636
M2625 727 325 1278 vdd hvtpfet l=6e-08 w=4.8e-07 $X=26653 $Y=10476 $D=636
M2626 356 363 725 vdd hvtpfet l=6e-08 w=3.2e-07 $X=26658 $Y=35913 $D=636
M2627 vdd tm<7> 726 vdd hvtpfet l=6e-08 w=4.11e-07 $X=26820 $Y=40177 $D=636
M2628 1283 123 vdd vdd hvtpfet l=6e-08 w=4.8e-07 $X=26839 $Y=33942 $D=636
M2629 729 123 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=26894 $Y=29274 $D=636
M2630 1285 369 352 vdd hvtpfet l=6e-08 w=4.11e-07 $X=26909 $Y=15932 $D=636
M2631 1286 369 353 vdd hvtpfet l=6e-08 w=4.11e-07 $X=26909 $Y=20589 $D=636
M2632 1287 369 354 vdd hvtpfet l=6e-08 w=4.11e-07 $X=26909 $Y=22852 $D=636
M2633 1288 369 355 vdd hvtpfet l=6e-08 w=4.11e-07 $X=26909 $Y=27509 $D=636
M2634 1284 362 356 vdd hvtpfet l=6e-08 w=4.8e-07 $X=26918 $Y=35753 $D=636
M2635 vdd aa<10> 374 vdd hvtpfet l=6e-08 w=4.11e-07 $X=26924 $Y=14280 $D=636
M2636 379 131 1283 vdd hvtpfet l=6e-08 w=4.8e-07 $X=27099 $Y=33942 $D=636
M2637 b_pxca_n<3> 370 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=27140 $Y=1941 $D=636
M2638 370 371 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=27140 $Y=5141 $D=636
M2639 371 351 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=27140 $Y=8691 $D=636
M2640 372 351 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=27140 $Y=41842 $D=636
M2641 373 372 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=27140 $Y=44992 $D=636
M2642 t_pxca_n<3> 373 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=27140 $Y=46622 $D=636
M2643 vdd 123 729 vdd hvtpfet l=6e-08 w=6e-07 $X=27154 $Y=29274 $D=636
M2644 vdd tm<9> 325 vdd hvtpfet l=7e-08 w=4.8e-07 $X=27163 $Y=10476 $D=636
M2645 vdd 376 1284 vdd hvtpfet l=6e-08 w=4.8e-07 $X=27178 $Y=35753 $D=636
M2646 vdd 317 1285 vdd hvtpfet l=6e-08 w=8.23e-07 $X=27179 $Y=15520 $D=636
M2647 vdd 317 1286 vdd hvtpfet l=6e-08 w=8.23e-07 $X=27179 $Y=20589 $D=636
M2648 vdd 317 1287 vdd hvtpfet l=6e-08 w=8.23e-07 $X=27179 $Y=22440 $D=636
M2649 vdd 317 1288 vdd hvtpfet l=6e-08 w=8.23e-07 $X=27179 $Y=27509 $D=636
M2650 375 374 vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=27184 $Y=14280 $D=636
M2651 736 377 379 vdd hvtpfet l=6e-08 w=3.2e-07 $X=27359 $Y=33942 $D=636
M2652 vdd 370 b_pxca_n<3> vdd hvtpfet l=6e-08 w=2.57e-06 $X=27400 $Y=1941 $D=636
M2653 vdd 371 370 vdd hvtpfet l=6e-08 w=1e-06 $X=27400 $Y=5141 $D=636
M2654 vdd 351 371 vdd hvtpfet l=6e-08 w=6e-07 $X=27400 $Y=8691 $D=636
M2655 vdd 351 372 vdd hvtpfet l=6e-08 w=6e-07 $X=27400 $Y=41842 $D=636
M2656 vdd 372 373 vdd hvtpfet l=6e-08 w=1e-06 $X=27400 $Y=44992 $D=636
M2657 vdd 373 t_pxca_n<3> vdd hvtpfet l=6e-08 w=2.57e-06 $X=27400 $Y=46622 $D=636
M2658 366 tm<8> vdd vdd hvtpfet l=7e-08 w=4.8e-07 $X=27433 $Y=10476 $D=636
M2659 vdd 123 736 vdd hvtpfet l=6e-08 w=3.2e-07 $X=27619 $Y=33942 $D=636
M2660 vdd tm<1> 735 vdd hvtpfet l=6e-08 w=4.11e-07 $X=27620 $Y=40177 $D=636
M2661 317 323 vdd vdd hvtpfet l=6e-08 w=7e-07 $X=27664 $Y=29648 $D=636
M2662 1289 374 352 vdd hvtpfet l=6e-08 w=4.11e-07 $X=27689 $Y=15932 $D=636
M2663 1290 375 353 vdd hvtpfet l=6e-08 w=4.11e-07 $X=27689 $Y=20589 $D=636
M2664 1291 374 354 vdd hvtpfet l=6e-08 w=4.11e-07 $X=27689 $Y=22852 $D=636
M2665 1292 375 355 vdd hvtpfet l=6e-08 w=4.11e-07 $X=27689 $Y=27509 $D=636
M2666 vdd 380 369 vdd hvtpfet l=6e-08 w=4.11e-07 $X=27784 $Y=14280 $D=636
M2667 vdd 362 386 vdd hvtpfet l=6e-08 w=4e-07 $X=27858 $Y=35682 $D=636
M2668 377 379 vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=27879 $Y=33942 $D=636
M2669 b_pxca_n<2> 381 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=27910 $Y=1941 $D=636
M2670 381 382 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=27910 $Y=5141 $D=636
M2671 382 350 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=27910 $Y=8691 $D=636
M2672 383 350 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=27910 $Y=41842 $D=636
M2673 384 383 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=27910 $Y=44992 $D=636
M2674 t_pxca_n<2> 384 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=27910 $Y=46622 $D=636
M2675 vdd 323 317 vdd hvtpfet l=6e-08 w=7e-07 $X=27924 $Y=29648 $D=636
M2676 vdd 317 1289 vdd hvtpfet l=6e-08 w=8.23e-07 $X=27959 $Y=15520 $D=636
M2677 vdd 317 1290 vdd hvtpfet l=6e-08 w=8.23e-07 $X=27959 $Y=20589 $D=636
M2678 vdd 317 1291 vdd hvtpfet l=6e-08 w=8.23e-07 $X=27959 $Y=22440 $D=636
M2679 vdd 317 1292 vdd hvtpfet l=6e-08 w=8.23e-07 $X=27959 $Y=27509 $D=636
M2680 380 aa<11> vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=28044 $Y=14280 $D=636
M2681 386 356 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=28118 $Y=35682 $D=636
M2682 vdd 381 b_pxca_n<2> vdd hvtpfet l=6e-08 w=2.57e-06 $X=28170 $Y=1941 $D=636
M2683 vdd 382 381 vdd hvtpfet l=6e-08 w=1e-06 $X=28170 $Y=5141 $D=636
M2684 vdd 350 382 vdd hvtpfet l=6e-08 w=6e-07 $X=28170 $Y=8691 $D=636
M2685 vdd 350 383 vdd hvtpfet l=6e-08 w=6e-07 $X=28170 $Y=41842 $D=636
M2686 vdd 383 384 vdd hvtpfet l=6e-08 w=1e-06 $X=28170 $Y=44992 $D=636
M2687 vdd 384 t_pxca_n<2> vdd hvtpfet l=6e-08 w=2.57e-06 $X=28170 $Y=46622 $D=636
M2688 317 323 vdd vdd hvtpfet l=6e-08 w=7e-07 $X=28184 $Y=29648 $D=636
M2689 1293 317 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=28219 $Y=15520 $D=636
M2690 1294 317 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=28219 $Y=20589 $D=636
M2691 1295 317 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=28219 $Y=22440 $D=636
M2692 1296 317 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=28219 $Y=27509 $D=636
M2693 vdd 323 317 vdd hvtpfet l=6e-08 w=7e-07 $X=28444 $Y=29648 $D=636
M2694 407 374 1293 vdd hvtpfet l=6e-08 w=4.11e-07 $X=28489 $Y=15932 $D=636
M2695 408 375 1294 vdd hvtpfet l=6e-08 w=4.11e-07 $X=28489 $Y=20589 $D=636
M2696 409 374 1295 vdd hvtpfet l=6e-08 w=4.11e-07 $X=28489 $Y=22852 $D=636
M2697 410 375 1296 vdd hvtpfet l=6e-08 w=4.11e-07 $X=28489 $Y=27509 $D=636
M2698 vdd 392 541 vdd hvtpfet l=6e-08 w=4e-07 $X=28514 $Y=10167 $D=636
M2699 vdd 393 544 vdd hvtpfet l=6e-08 w=4e-07 $X=28514 $Y=40566 $D=636
M2700 494 386 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=28628 $Y=35682 $D=636
M2701 b_pxca_n<1> 387 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=28680 $Y=1941 $D=636
M2702 387 388 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=28680 $Y=5141 $D=636
M2703 388 389 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=28680 $Y=8691 $D=636
M2704 390 389 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=28680 $Y=41842 $D=636
M2705 391 390 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=28680 $Y=44992 $D=636
M2706 t_pxca_n<1> 391 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=28680 $Y=46622 $D=636
M2707 742 123 vdd vdd hvtpfet l=6e-08 w=1.2e-06 $X=28704 $Y=29148 $D=636
M2708 vdd 387 b_pxca_n<1> vdd hvtpfet l=6e-08 w=2.57e-06 $X=28940 $Y=1941 $D=636
M2709 vdd 388 387 vdd hvtpfet l=6e-08 w=1e-06 $X=28940 $Y=5141 $D=636
M2710 vdd 389 388 vdd hvtpfet l=6e-08 w=6e-07 $X=28940 $Y=8691 $D=636
M2711 vdd 389 390 vdd hvtpfet l=6e-08 w=6e-07 $X=28940 $Y=41842 $D=636
M2712 vdd 390 391 vdd hvtpfet l=6e-08 w=1e-06 $X=28940 $Y=44992 $D=636
M2713 vdd 391 t_pxca_n<1> vdd hvtpfet l=6e-08 w=2.57e-06 $X=28940 $Y=46622 $D=636
M2714 1297 317 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=28999 $Y=15520 $D=636
M2715 1298 317 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=28999 $Y=20589 $D=636
M2716 1299 317 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=28999 $Y=22440 $D=636
M2717 1300 317 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=28999 $Y=27509 $D=636
M2718 vdd 308 392 vdd hvtpfet l=6e-08 w=4.11e-07 $X=29024 $Y=10156 $D=636
M2719 vdd 308 393 vdd hvtpfet l=6e-08 w=4.11e-07 $X=29024 $Y=40566 $D=636
M2720 vdd aa<12> 365 vdd hvtpfet l=6e-08 w=4.11e-07 $X=29054 $Y=14280 $D=636
M2721 407 380 1297 vdd hvtpfet l=6e-08 w=4.11e-07 $X=29269 $Y=15932 $D=636
M2722 408 380 1298 vdd hvtpfet l=6e-08 w=4.11e-07 $X=29269 $Y=20589 $D=636
M2723 409 380 1299 vdd hvtpfet l=6e-08 w=4.11e-07 $X=29269 $Y=22852 $D=636
M2724 410 380 1300 vdd hvtpfet l=6e-08 w=4.11e-07 $X=29269 $Y=27509 $D=636
M2725 392 dwla<1> vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=29284 $Y=10156 $D=636
M2726 393 dwla<0> vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=29284 $Y=40566 $D=636
M2727 743 395 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=29298 $Y=33468 $D=636
M2728 b_pxca_n<0> 396 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=29450 $Y=1941 $D=636
M2729 396 397 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=29450 $Y=5141 $D=636
M2730 397 398 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=29450 $Y=8691 $D=636
M2731 399 398 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=29450 $Y=41842 $D=636
M2732 400 399 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=29450 $Y=44992 $D=636
M2733 t_pxca_n<0> 400 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=29450 $Y=46622 $D=636
M2734 748 403 456 vdd hvtpfet l=6e-08 w=1e-06 $X=29487 $Y=35707 $D=636
M2735 1301 364 407 vdd hvtpfet l=6e-08 w=4.11e-07 $X=29529 $Y=15932 $D=636
M2736 1302 364 408 vdd hvtpfet l=6e-08 w=4.11e-07 $X=29529 $Y=20589 $D=636
M2737 1303 365 409 vdd hvtpfet l=6e-08 w=4.11e-07 $X=29529 $Y=22852 $D=636
M2738 1304 365 410 vdd hvtpfet l=6e-08 w=4.11e-07 $X=29529 $Y=27509 $D=636
M2739 403 405 743 vdd hvtpfet l=6e-08 w=6e-07 $X=29558 $Y=33468 $D=636
M2740 364 365 vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=29564 $Y=14280 $D=636
M2741 vdd 404 395 vdd hvtpfet l=2.5e-07 w=5e-07 $X=29591 $Y=29813 $D=636
M2742 vdd 396 b_pxca_n<0> vdd hvtpfet l=6e-08 w=2.57e-06 $X=29710 $Y=1941 $D=636
M2743 vdd 397 396 vdd hvtpfet l=6e-08 w=1e-06 $X=29710 $Y=5141 $D=636
M2744 vdd 398 397 vdd hvtpfet l=6e-08 w=6e-07 $X=29710 $Y=8691 $D=636
M2745 vdd 398 399 vdd hvtpfet l=6e-08 w=6e-07 $X=29710 $Y=41842 $D=636
M2746 vdd 399 400 vdd hvtpfet l=6e-08 w=1e-06 $X=29710 $Y=44992 $D=636
M2747 vdd 400 t_pxca_n<0> vdd hvtpfet l=6e-08 w=2.57e-06 $X=29710 $Y=46622 $D=636
M2748 456 403 748 vdd hvtpfet l=6e-08 w=1e-06 $X=29747 $Y=35707 $D=636
M2749 vdd 317 1301 vdd hvtpfet l=6e-08 w=8.23e-07 $X=29799 $Y=15520 $D=636
M2750 vdd 317 1302 vdd hvtpfet l=6e-08 w=8.23e-07 $X=29799 $Y=20589 $D=636
M2751 vdd 317 1303 vdd hvtpfet l=6e-08 w=8.23e-07 $X=29799 $Y=22440 $D=636
M2752 vdd 317 1304 vdd hvtpfet l=6e-08 w=8.23e-07 $X=29799 $Y=27509 $D=636
M2753 748 403 456 vdd hvtpfet l=6e-08 w=1e-06 $X=30007 $Y=35707 $D=636
M2754 404 406 vdd vdd hvtpfet l=6e-08 w=5e-07 $X=30041 $Y=29813 $D=636
M2755 405 tm<7> vdd vdd hvtpfet l=6e-08 w=3e-07 $X=30068 $Y=33468 $D=636
M2756 dbl_pd_n<3> 131 vdd vdd hvtpfet l=6e-08 w=4.28e-07 $X=30204 $Y=14263 $D=636
M2757 b_pxba_n<7> 411 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=30220 $Y=1941 $D=636
M2758 411 412 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=30220 $Y=5141 $D=636
M2759 412 413 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=30220 $Y=8691 $D=636
M2760 414 413 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=30220 $Y=41842 $D=636
M2761 415 414 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=30220 $Y=44992 $D=636
M2762 t_pxba_n<7> 415 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=30220 $Y=46622 $D=636
M2763 753 416 748 vdd hvtpfet l=6e-08 w=1e-06 $X=30267 $Y=35707 $D=636
M2764 359 407 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=30309 $Y=15321 $D=636
M2765 1305 323 407 vdd hvtpfet l=6e-08 w=2.74e-07 $X=30309 $Y=16069 $D=636
M2766 1306 323 408 vdd hvtpfet l=6e-08 w=2.74e-07 $X=30309 $Y=20589 $D=636
M2767 347 408 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=30309 $Y=21405 $D=636
M2768 398 409 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=30309 $Y=22241 $D=636
M2769 1307 323 409 vdd hvtpfet l=6e-08 w=2.74e-07 $X=30309 $Y=22989 $D=636
M2770 1308 323 410 vdd hvtpfet l=6e-08 w=2.74e-07 $X=30309 $Y=27509 $D=636
M2771 389 410 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=30309 $Y=28325 $D=636
M2772 vdd 131 dbl_pd_n<3> vdd hvtpfet l=6e-08 w=4.28e-07 $X=30464 $Y=14263 $D=636
M2773 vdd 411 b_pxba_n<7> vdd hvtpfet l=6e-08 w=2.57e-06 $X=30480 $Y=1941 $D=636
M2774 vdd 412 411 vdd hvtpfet l=6e-08 w=1e-06 $X=30480 $Y=5141 $D=636
M2775 vdd 413 412 vdd hvtpfet l=6e-08 w=6e-07 $X=30480 $Y=8691 $D=636
M2776 vdd 413 414 vdd hvtpfet l=6e-08 w=6e-07 $X=30480 $Y=41842 $D=636
M2777 vdd 414 415 vdd hvtpfet l=6e-08 w=1e-06 $X=30480 $Y=44992 $D=636
M2778 vdd 415 t_pxba_n<7> vdd hvtpfet l=6e-08 w=2.57e-06 $X=30480 $Y=46622 $D=636
M2779 748 416 753 vdd hvtpfet l=6e-08 w=1e-06 $X=30527 $Y=35707 $D=636
M2780 vdd 407 359 vdd hvtpfet l=6e-08 w=2.06e-07 $X=30569 $Y=15321 $D=636
M2781 vdd 359 1305 vdd hvtpfet l=6e-08 w=2.74e-07 $X=30569 $Y=16069 $D=636
M2782 vdd 347 1306 vdd hvtpfet l=6e-08 w=2.74e-07 $X=30569 $Y=20589 $D=636
M2783 vdd 408 347 vdd hvtpfet l=6e-08 w=2.06e-07 $X=30569 $Y=21405 $D=636
M2784 vdd 409 398 vdd hvtpfet l=6e-08 w=2.06e-07 $X=30569 $Y=22241 $D=636
M2785 vdd 398 1307 vdd hvtpfet l=6e-08 w=2.74e-07 $X=30569 $Y=22989 $D=636
M2786 vdd 389 1308 vdd hvtpfet l=6e-08 w=2.74e-07 $X=30569 $Y=27509 $D=636
M2787 vdd 410 389 vdd hvtpfet l=6e-08 w=2.06e-07 $X=30569 $Y=28325 $D=636
M2788 vdd dwla<1> 426 vdd hvtpfet l=6e-08 w=4.11e-07 $X=30584 $Y=10156 $D=636
M2789 vdd dwla<0> 427 vdd hvtpfet l=6e-08 w=4.11e-07 $X=30584 $Y=40566 $D=636
M2790 749 406 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=30644 $Y=33468 $D=636
M2791 vdd 417 406 vdd hvtpfet l=2.5e-07 w=5e-07 $X=30711 $Y=29813 $D=636
M2792 dbl_pd_n<3> 131 vdd vdd hvtpfet l=6e-08 w=4.28e-07 $X=30724 $Y=14263 $D=636
M2793 753 416 748 vdd hvtpfet l=6e-08 w=1e-06 $X=30787 $Y=35707 $D=636
M2794 426 309 vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=30844 $Y=10156 $D=636
M2795 427 309 vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=30844 $Y=40566 $D=636
M2796 416 423 749 vdd hvtpfet l=6e-08 w=6e-07 $X=30904 $Y=33468 $D=636
M2797 b_pxba_n<6> 418 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=30990 $Y=1941 $D=636
M2798 418 419 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=30990 $Y=5141 $D=636
M2799 419 420 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=30990 $Y=8691 $D=636
M2800 421 420 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=30990 $Y=41842 $D=636
M2801 422 421 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=30990 $Y=44992 $D=636
M2802 t_pxba_n<6> 422 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=30990 $Y=46622 $D=636
M2803 vdd 362 753 vdd hvtpfet l=6e-08 w=1e-06 $X=31047 $Y=35707 $D=636
M2804 420 428 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=31079 $Y=15321 $D=636
M2805 1309 420 vdd vdd hvtpfet l=6e-08 w=2.74e-07 $X=31079 $Y=16069 $D=636
M2806 1310 413 vdd vdd hvtpfet l=6e-08 w=2.74e-07 $X=31079 $Y=20589 $D=636
M2807 413 429 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=31079 $Y=21405 $D=636
M2808 424 430 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=31079 $Y=22241 $D=636
M2809 1311 424 vdd vdd hvtpfet l=6e-08 w=2.74e-07 $X=31079 $Y=22989 $D=636
M2810 1312 425 vdd vdd hvtpfet l=6e-08 w=2.74e-07 $X=31079 $Y=27509 $D=636
M2811 425 431 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=31079 $Y=28325 $D=636
M2812 417 368 vdd vdd hvtpfet l=6e-08 w=5e-07 $X=31161 $Y=29813 $D=636
M2813 dbl_pd_n<1> tm<1> vdd vdd hvtpfet l=6e-08 w=4.28e-07 $X=31234 $Y=14263 $D=636
M2814 vdd 418 b_pxba_n<6> vdd hvtpfet l=6e-08 w=2.57e-06 $X=31250 $Y=1941 $D=636
M2815 vdd 419 418 vdd hvtpfet l=6e-08 w=1e-06 $X=31250 $Y=5141 $D=636
M2816 vdd 420 419 vdd hvtpfet l=6e-08 w=6e-07 $X=31250 $Y=8691 $D=636
M2817 vdd 420 421 vdd hvtpfet l=6e-08 w=6e-07 $X=31250 $Y=41842 $D=636
M2818 vdd 421 422 vdd hvtpfet l=6e-08 w=1e-06 $X=31250 $Y=44992 $D=636
M2819 vdd 422 t_pxba_n<6> vdd hvtpfet l=6e-08 w=2.57e-06 $X=31250 $Y=46622 $D=636
M2820 753 362 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=31307 $Y=35707 $D=636
M2821 vdd 428 420 vdd hvtpfet l=6e-08 w=2.06e-07 $X=31339 $Y=15321 $D=636
M2822 428 323 1309 vdd hvtpfet l=6e-08 w=2.74e-07 $X=31339 $Y=16069 $D=636
M2823 429 323 1310 vdd hvtpfet l=6e-08 w=2.74e-07 $X=31339 $Y=20589 $D=636
M2824 vdd 429 413 vdd hvtpfet l=6e-08 w=2.06e-07 $X=31339 $Y=21405 $D=636
M2825 vdd 430 424 vdd hvtpfet l=6e-08 w=2.06e-07 $X=31339 $Y=22241 $D=636
M2826 430 323 1311 vdd hvtpfet l=6e-08 w=2.74e-07 $X=31339 $Y=22989 $D=636
M2827 431 323 1312 vdd hvtpfet l=6e-08 w=2.74e-07 $X=31339 $Y=27509 $D=636
M2828 vdd 431 425 vdd hvtpfet l=6e-08 w=2.06e-07 $X=31339 $Y=28325 $D=636
M2829 556 426 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=31354 $Y=10167 $D=636
M2830 558 427 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=31354 $Y=40566 $D=636
M2831 vdd 173 423 vdd hvtpfet l=6e-08 w=3e-07 $X=31414 $Y=33468 $D=636
M2832 vdd tm<1> dbl_pd_n<1> vdd hvtpfet l=6e-08 w=4.28e-07 $X=31494 $Y=14263 $D=636
M2833 vdd 362 753 vdd hvtpfet l=6e-08 w=1e-06 $X=31567 $Y=35707 $D=636
M2834 dbl_pd_n<1> tm<1> vdd vdd hvtpfet l=6e-08 w=4.28e-07 $X=31754 $Y=14263 $D=636
M2835 b_pxba_n<5> 432 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=31760 $Y=1941 $D=636
M2836 432 433 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=31760 $Y=5141 $D=636
M2837 433 434 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=31760 $Y=8691 $D=636
M2838 435 434 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=31760 $Y=41842 $D=636
M2839 436 435 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=31760 $Y=44992 $D=636
M2840 t_pxba_n<5> 436 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=31760 $Y=46622 $D=636
M2841 vdd 368 362 vdd hvtpfet l=6e-08 w=4e-07 $X=31761 $Y=29948 $D=636
M2842 1313 317 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=31849 $Y=15520 $D=636
M2843 1314 317 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=31849 $Y=20589 $D=636
M2844 1315 317 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=31849 $Y=22440 $D=636
M2845 1316 317 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=31849 $Y=27509 $D=636
M2846 vdd 437 540 vdd hvtpfet l=6e-08 w=4e-07 $X=31864 $Y=10167 $D=636
M2847 vdd 438 545 vdd hvtpfet l=6e-08 w=4e-07 $X=31864 $Y=40566 $D=636
M2848 vdd 432 b_pxba_n<5> vdd hvtpfet l=6e-08 w=2.57e-06 $X=32020 $Y=1941 $D=636
M2849 vdd 433 432 vdd hvtpfet l=6e-08 w=1e-06 $X=32020 $Y=5141 $D=636
M2850 vdd 434 433 vdd hvtpfet l=6e-08 w=6e-07 $X=32020 $Y=8691 $D=636
M2851 vdd 434 435 vdd hvtpfet l=6e-08 w=6e-07 $X=32020 $Y=41842 $D=636
M2852 vdd 435 436 vdd hvtpfet l=6e-08 w=1e-06 $X=32020 $Y=44992 $D=636
M2853 vdd 436 t_pxba_n<5> vdd hvtpfet l=6e-08 w=2.57e-06 $X=32020 $Y=46622 $D=636
M2854 428 439 1313 vdd hvtpfet l=6e-08 w=4.11e-07 $X=32119 $Y=15932 $D=636
M2855 429 439 1314 vdd hvtpfet l=6e-08 w=4.11e-07 $X=32119 $Y=20589 $D=636
M2856 430 440 1315 vdd hvtpfet l=6e-08 w=4.11e-07 $X=32119 $Y=22852 $D=636
M2857 431 440 1316 vdd hvtpfet l=6e-08 w=4.11e-07 $X=32119 $Y=27509 $D=636
M2858 761 442 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=32271 $Y=29348 $D=636
M2859 762 442 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=32271 $Y=35707 $D=636
M2860 vdd 310 437 vdd hvtpfet l=6e-08 w=4.11e-07 $X=32374 $Y=10156 $D=636
M2861 vdd 310 438 vdd hvtpfet l=6e-08 w=4.11e-07 $X=32374 $Y=40566 $D=636
M2862 1317 443 428 vdd hvtpfet l=6e-08 w=4.11e-07 $X=32379 $Y=15932 $D=636
M2863 1318 443 429 vdd hvtpfet l=6e-08 w=4.11e-07 $X=32379 $Y=20589 $D=636
M2864 1319 443 430 vdd hvtpfet l=6e-08 w=4.11e-07 $X=32379 $Y=22852 $D=636
M2865 1320 443 431 vdd hvtpfet l=6e-08 w=4.11e-07 $X=32379 $Y=27509 $D=636
M2866 vdd aa<7> 449 vdd hvtpfet l=6e-08 w=4.11e-07 $X=32394 $Y=14280 $D=636
M2867 vdd 324 442 vdd hvtpfet l=6e-08 w=1e-06 $X=32394 $Y=33493 $D=636
M2868 b_pxba_n<4> 444 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=32530 $Y=1941 $D=636
M2869 444 445 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=32530 $Y=5141 $D=636
M2870 445 446 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=32530 $Y=8691 $D=636
M2871 447 446 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=32530 $Y=41842 $D=636
M2872 448 447 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=32530 $Y=44992 $D=636
M2873 t_pxba_n<4> 448 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=32530 $Y=46622 $D=636
M2874 vdd 442 761 vdd hvtpfet l=6e-08 w=1e-06 $X=32531 $Y=29348 $D=636
M2875 vdd 442 762 vdd hvtpfet l=6e-08 w=1e-06 $X=32531 $Y=35707 $D=636
M2876 437 dwla<1> vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=32634 $Y=10156 $D=636
M2877 438 dwla<0> vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=32634 $Y=40566 $D=636
M2878 vdd 317 1317 vdd hvtpfet l=6e-08 w=8.23e-07 $X=32649 $Y=15520 $D=636
M2879 vdd 317 1318 vdd hvtpfet l=6e-08 w=8.23e-07 $X=32649 $Y=20589 $D=636
M2880 vdd 317 1319 vdd hvtpfet l=6e-08 w=8.23e-07 $X=32649 $Y=22440 $D=636
M2881 vdd 317 1320 vdd hvtpfet l=6e-08 w=8.23e-07 $X=32649 $Y=27509 $D=636
M2882 450 449 vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=32654 $Y=14280 $D=636
M2883 vdd 444 b_pxba_n<4> vdd hvtpfet l=6e-08 w=2.57e-06 $X=32790 $Y=1941 $D=636
M2884 vdd 445 444 vdd hvtpfet l=6e-08 w=1e-06 $X=32790 $Y=5141 $D=636
M2885 vdd 446 445 vdd hvtpfet l=6e-08 w=6e-07 $X=32790 $Y=8691 $D=636
M2886 vdd 446 447 vdd hvtpfet l=6e-08 w=6e-07 $X=32790 $Y=41842 $D=636
M2887 vdd 447 448 vdd hvtpfet l=6e-08 w=1e-06 $X=32790 $Y=44992 $D=636
M2888 vdd 448 t_pxba_n<4> vdd hvtpfet l=6e-08 w=2.57e-06 $X=32790 $Y=46622 $D=636
M2889 dwla<1> 368 761 vdd hvtpfet l=6e-08 w=1e-06 $X=33041 $Y=29348 $D=636
M2890 497 456 762 vdd hvtpfet l=6e-08 w=1e-06 $X=33041 $Y=35707 $D=636
M2891 465 442 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=33094 $Y=33493 $D=636
M2892 vdd dwla<1> 458 vdd hvtpfet l=6e-08 w=4.11e-07 $X=33144 $Y=10156 $D=636
M2893 vdd dwla<0> 459 vdd hvtpfet l=6e-08 w=4.11e-07 $X=33144 $Y=40566 $D=636
M2894 1321 449 428 vdd hvtpfet l=6e-08 w=4.11e-07 $X=33159 $Y=15932 $D=636
M2895 1322 450 429 vdd hvtpfet l=6e-08 w=4.11e-07 $X=33159 $Y=20589 $D=636
M2896 1323 449 430 vdd hvtpfet l=6e-08 w=4.11e-07 $X=33159 $Y=22852 $D=636
M2897 1324 450 431 vdd hvtpfet l=6e-08 w=4.11e-07 $X=33159 $Y=27509 $D=636
M2898 vdd 455 443 vdd hvtpfet l=6e-08 w=4.11e-07 $X=33254 $Y=14280 $D=636
M2899 b_pxba_n<3> 451 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=33300 $Y=1941 $D=636
M2900 451 452 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=33300 $Y=5141 $D=636
M2901 452 425 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=33300 $Y=8691 $D=636
M2902 453 425 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=33300 $Y=41842 $D=636
M2903 454 453 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=33300 $Y=44992 $D=636
M2904 t_pxba_n<3> 454 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=33300 $Y=46622 $D=636
M2905 761 368 dwla<1> vdd hvtpfet l=6e-08 w=1e-06 $X=33301 $Y=29348 $D=636
M2906 762 456 497 vdd hvtpfet l=6e-08 w=1e-06 $X=33301 $Y=35707 $D=636
M2907 458 311 vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=33404 $Y=10156 $D=636
M2908 459 311 vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=33404 $Y=40566 $D=636
M2909 vdd 317 1321 vdd hvtpfet l=6e-08 w=8.23e-07 $X=33429 $Y=15520 $D=636
M2910 vdd 317 1322 vdd hvtpfet l=6e-08 w=8.23e-07 $X=33429 $Y=20589 $D=636
M2911 vdd 317 1323 vdd hvtpfet l=6e-08 w=8.23e-07 $X=33429 $Y=22440 $D=636
M2912 vdd 317 1324 vdd hvtpfet l=6e-08 w=8.23e-07 $X=33429 $Y=27509 $D=636
M2913 455 aa<8> vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=33514 $Y=14280 $D=636
M2914 vdd 451 b_pxba_n<3> vdd hvtpfet l=6e-08 w=2.57e-06 $X=33560 $Y=1941 $D=636
M2915 vdd 452 451 vdd hvtpfet l=6e-08 w=1e-06 $X=33560 $Y=5141 $D=636
M2916 vdd 425 452 vdd hvtpfet l=6e-08 w=6e-07 $X=33560 $Y=8691 $D=636
M2917 vdd 425 453 vdd hvtpfet l=6e-08 w=6e-07 $X=33560 $Y=41842 $D=636
M2918 vdd 453 454 vdd hvtpfet l=6e-08 w=1e-06 $X=33560 $Y=44992 $D=636
M2919 vdd 454 t_pxba_n<3> vdd hvtpfet l=6e-08 w=2.57e-06 $X=33560 $Y=46622 $D=636
M2920 1325 317 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=33689 $Y=15520 $D=636
M2921 1326 317 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=33689 $Y=20589 $D=636
M2922 1327 317 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=33689 $Y=22440 $D=636
M2923 1328 317 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=33689 $Y=27509 $D=636
M2924 dwla<0> 368 765 vdd hvtpfet l=6e-08 w=1e-06 $X=33811 $Y=29348 $D=636
M2925 498 456 766 vdd hvtpfet l=6e-08 w=1e-06 $X=33811 $Y=35707 $D=636
M2926 555 458 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=33914 $Y=10167 $D=636
M2927 559 459 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=33914 $Y=40566 $D=636
M2928 479 449 1325 vdd hvtpfet l=6e-08 w=4.11e-07 $X=33959 $Y=15932 $D=636
M2929 480 450 1326 vdd hvtpfet l=6e-08 w=4.11e-07 $X=33959 $Y=20589 $D=636
M2930 481 449 1327 vdd hvtpfet l=6e-08 w=4.11e-07 $X=33959 $Y=22852 $D=636
M2931 482 450 1328 vdd hvtpfet l=6e-08 w=4.11e-07 $X=33959 $Y=27509 $D=636
M2932 b_pxba_n<2> 460 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=34070 $Y=1941 $D=636
M2933 460 461 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=34070 $Y=5141 $D=636
M2934 461 424 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=34070 $Y=8691 $D=636
M2935 462 424 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=34070 $Y=41842 $D=636
M2936 463 462 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=34070 $Y=44992 $D=636
M2937 t_pxba_n<2> 463 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=34070 $Y=46622 $D=636
M2938 765 368 dwla<0> vdd hvtpfet l=6e-08 w=1e-06 $X=34071 $Y=29348 $D=636
M2939 766 456 498 vdd hvtpfet l=6e-08 w=1e-06 $X=34071 $Y=35707 $D=636
M2940 vdd 460 b_pxba_n<2> vdd hvtpfet l=6e-08 w=2.57e-06 $X=34330 $Y=1941 $D=636
M2941 vdd 461 460 vdd hvtpfet l=6e-08 w=1e-06 $X=34330 $Y=5141 $D=636
M2942 vdd 424 461 vdd hvtpfet l=6e-08 w=6e-07 $X=34330 $Y=8691 $D=636
M2943 vdd 424 462 vdd hvtpfet l=6e-08 w=6e-07 $X=34330 $Y=41842 $D=636
M2944 vdd 462 463 vdd hvtpfet l=6e-08 w=1e-06 $X=34330 $Y=44992 $D=636
M2945 vdd 463 t_pxba_n<2> vdd hvtpfet l=6e-08 w=2.57e-06 $X=34330 $Y=46622 $D=636
M2946 1329 317 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=34469 $Y=15520 $D=636
M2947 1330 317 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=34469 $Y=20589 $D=636
M2948 1331 317 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=34469 $Y=22440 $D=636
M2949 1332 317 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=34469 $Y=27509 $D=636
M2950 vdd aa<9> 440 vdd hvtpfet l=6e-08 w=4.11e-07 $X=34524 $Y=14280 $D=636
M2951 765 465 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=34581 $Y=29348 $D=636
M2952 766 465 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=34581 $Y=35707 $D=636
M2953 vdd vdd 535 vdd hvtpfet l=6e-08 w=6.4e-07 $X=34621 $Y=33468 $D=636
M2954 479 455 1329 vdd hvtpfet l=6e-08 w=4.11e-07 $X=34739 $Y=15932 $D=636
M2955 480 455 1330 vdd hvtpfet l=6e-08 w=4.11e-07 $X=34739 $Y=20589 $D=636
M2956 481 455 1331 vdd hvtpfet l=6e-08 w=4.11e-07 $X=34739 $Y=22852 $D=636
M2957 482 455 1332 vdd hvtpfet l=6e-08 w=4.11e-07 $X=34739 $Y=27509 $D=636
M2958 b_pxba_n<1> 466 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=34840 $Y=1941 $D=636
M2959 466 467 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=34840 $Y=5141 $D=636
M2960 467 468 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=34840 $Y=8691 $D=636
M2961 469 468 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=34840 $Y=41842 $D=636
M2962 470 469 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=34840 $Y=44992 $D=636
M2963 t_pxba_n<1> 470 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=34840 $Y=46622 $D=636
M2964 vdd 465 765 vdd hvtpfet l=6e-08 w=1e-06 $X=34841 $Y=29348 $D=636
M2965 vdd 465 766 vdd hvtpfet l=6e-08 w=1e-06 $X=34841 $Y=35707 $D=636
M2966 535 471 vdd vdd hvtpfet l=6e-08 w=6.4e-07 $X=34881 $Y=33468 $D=636
M2967 vdd 123 131 vdd hvtpfet l=6e-08 w=2e-07 $X=34906 $Y=10756 $D=636
M2968 1333 439 479 vdd hvtpfet l=6e-08 w=4.11e-07 $X=34999 $Y=15932 $D=636
M2969 1334 439 480 vdd hvtpfet l=6e-08 w=4.11e-07 $X=34999 $Y=20589 $D=636
M2970 1335 440 481 vdd hvtpfet l=6e-08 w=4.11e-07 $X=34999 $Y=22852 $D=636
M2971 1336 440 482 vdd hvtpfet l=6e-08 w=4.11e-07 $X=34999 $Y=27509 $D=636
M2972 439 440 vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=35034 $Y=14280 $D=636
M2973 vdd 466 b_pxba_n<1> vdd hvtpfet l=6e-08 w=2.57e-06 $X=35100 $Y=1941 $D=636
M2974 vdd 467 466 vdd hvtpfet l=6e-08 w=1e-06 $X=35100 $Y=5141 $D=636
M2975 vdd 468 467 vdd hvtpfet l=6e-08 w=6e-07 $X=35100 $Y=8691 $D=636
M2976 vdd 468 469 vdd hvtpfet l=6e-08 w=6e-07 $X=35100 $Y=41842 $D=636
M2977 vdd 469 470 vdd hvtpfet l=6e-08 w=1e-06 $X=35100 $Y=44992 $D=636
M2978 vdd 470 t_pxba_n<1> vdd hvtpfet l=6e-08 w=2.57e-06 $X=35100 $Y=46622 $D=636
M2979 vdd 317 1333 vdd hvtpfet l=6e-08 w=8.23e-07 $X=35269 $Y=15520 $D=636
M2980 vdd 317 1334 vdd hvtpfet l=6e-08 w=8.23e-07 $X=35269 $Y=20589 $D=636
M2981 vdd 317 1335 vdd hvtpfet l=6e-08 w=8.23e-07 $X=35269 $Y=22440 $D=636
M2982 vdd 317 1336 vdd hvtpfet l=6e-08 w=8.23e-07 $X=35269 $Y=27509 $D=636
M2983 vdd 473 484 vdd hvtpfet l=6e-08 w=3e-07 $X=35351 $Y=36377 $D=636
M2984 vdd 472 471 vdd hvtpfet l=2.5e-07 w=5e-07 $X=35416 $Y=33503 $D=636
M2985 b_pxba_n<0> 474 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=35610 $Y=1941 $D=636
M2986 474 475 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=35610 $Y=5141 $D=636
M2987 475 476 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=35610 $Y=8691 $D=636
M2988 477 476 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=35610 $Y=41842 $D=636
M2989 478 477 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=35610 $Y=44992 $D=636
M2990 t_pxba_n<0> 478 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=35610 $Y=46622 $D=636
M2991 446 479 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=35779 $Y=15321 $D=636
M2992 1337 323 479 vdd hvtpfet l=6e-08 w=2.74e-07 $X=35779 $Y=16069 $D=636
M2993 1338 323 480 vdd hvtpfet l=6e-08 w=2.74e-07 $X=35779 $Y=20589 $D=636
M2994 434 480 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=35779 $Y=21405 $D=636
M2995 476 481 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=35779 $Y=22241 $D=636
M2996 1339 323 481 vdd hvtpfet l=6e-08 w=2.74e-07 $X=35779 $Y=22989 $D=636
M2997 1340 323 482 vdd hvtpfet l=6e-08 w=2.74e-07 $X=35779 $Y=27509 $D=636
M2998 468 482 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=35779 $Y=28325 $D=636
M2999 473 484 vdd vdd hvtpfet l=1.2e-07 w=3e-07 $X=35861 $Y=36382 $D=636
M3000 472 483 vdd vdd hvtpfet l=6e-08 w=5e-07 $X=35866 $Y=33503 $D=636
M3001 vdd 474 b_pxba_n<0> vdd hvtpfet l=6e-08 w=2.57e-06 $X=35870 $Y=1941 $D=636
M3002 vdd 475 474 vdd hvtpfet l=6e-08 w=1e-06 $X=35870 $Y=5141 $D=636
M3003 vdd 476 475 vdd hvtpfet l=6e-08 w=6e-07 $X=35870 $Y=8691 $D=636
M3004 vdd 476 477 vdd hvtpfet l=6e-08 w=6e-07 $X=35870 $Y=41842 $D=636
M3005 vdd 477 478 vdd hvtpfet l=6e-08 w=1e-06 $X=35870 $Y=44992 $D=636
M3006 vdd 478 t_pxba_n<0> vdd hvtpfet l=6e-08 w=2.57e-06 $X=35870 $Y=46622 $D=636
M3007 368 495 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=35945 $Y=29548 $D=636
M3008 vdd 479 446 vdd hvtpfet l=6e-08 w=2.06e-07 $X=36039 $Y=15321 $D=636
M3009 vdd 446 1337 vdd hvtpfet l=6e-08 w=2.74e-07 $X=36039 $Y=16069 $D=636
M3010 vdd 434 1338 vdd hvtpfet l=6e-08 w=2.74e-07 $X=36039 $Y=20589 $D=636
M3011 vdd 480 434 vdd hvtpfet l=6e-08 w=2.06e-07 $X=36039 $Y=21405 $D=636
M3012 vdd 481 476 vdd hvtpfet l=6e-08 w=2.06e-07 $X=36039 $Y=22241 $D=636
M3013 vdd 476 1339 vdd hvtpfet l=6e-08 w=2.74e-07 $X=36039 $Y=22989 $D=636
M3014 vdd 468 1340 vdd hvtpfet l=6e-08 w=2.74e-07 $X=36039 $Y=27509 $D=636
M3015 vdd 482 468 vdd hvtpfet l=6e-08 w=2.06e-07 $X=36039 $Y=28325 $D=636
M3016 vdd 495 368 vdd hvtpfet l=6e-08 w=8e-07 $X=36205 $Y=29548 $D=636
M3017 vdd 491 509 vdd hvtpfet l=6e-08 w=4.11e-07 $X=36254 $Y=14280 $D=636
M3018 b_pxaa<3> 485 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=36380 $Y=1941 $D=636
M3019 485 486 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=36380 $Y=5141 $D=636
M3020 486 487 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=36380 $Y=8691 $D=636
M3021 vdd 492 487 vdd hvtpfet l=6e-08 w=4.11e-07 $X=36380 $Y=10156 $D=636
M3022 vdd 492 488 vdd hvtpfet l=6e-08 w=4.11e-07 $X=36380 $Y=40566 $D=636
M3023 489 488 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=36380 $Y=41842 $D=636
M3024 490 489 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=36380 $Y=44992 $D=636
M3025 t_pxaa<3> 490 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=36380 $Y=46622 $D=636
M3026 vdd 493 473 vdd hvtpfet l=6e-08 w=6.4e-07 $X=36431 $Y=35802 $D=636
M3027 vdd 496 483 vdd hvtpfet l=6e-08 w=6.4e-07 $X=36466 $Y=33468 $D=636
M3028 vdd 485 b_pxaa<3> vdd hvtpfet l=6e-08 w=2.57e-06 $X=36640 $Y=1941 $D=636
M3029 vdd 486 485 vdd hvtpfet l=6e-08 w=1e-06 $X=36640 $Y=5141 $D=636
M3030 vdd 487 486 vdd hvtpfet l=6e-08 w=6e-07 $X=36640 $Y=8691 $D=636
M3031 487 497 vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=36640 $Y=10156 $D=636
M3032 488 498 vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=36640 $Y=40566 $D=636
M3033 vdd 488 489 vdd hvtpfet l=6e-08 w=6e-07 $X=36640 $Y=41842 $D=636
M3034 vdd 489 490 vdd hvtpfet l=6e-08 w=1e-06 $X=36640 $Y=44992 $D=636
M3035 vdd 490 t_pxaa<3> vdd hvtpfet l=6e-08 w=2.57e-06 $X=36640 $Y=46622 $D=636
M3036 368 clka vdd vdd hvtpfet l=6e-08 w=8e-07 $X=36715 $Y=29548 $D=636
M3037 491 aa<6> vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=36764 $Y=14280 $D=636
M3038 1341 317 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=36789 $Y=15520 $D=636
M3039 1342 317 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=36789 $Y=20589 $D=636
M3040 1343 317 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=36789 $Y=22440 $D=636
M3041 1344 317 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=36789 $Y=27509 $D=636
M3042 vdd clka 368 vdd hvtpfet l=6e-08 w=8e-07 $X=36975 $Y=29548 $D=636
M3043 vdd 473 496 vdd hvtpfet l=6e-08 w=6.4e-07 $X=36976 $Y=33693 $D=636
M3044 519 501 1341 vdd hvtpfet l=6e-08 w=4.11e-07 $X=37059 $Y=15932 $D=636
M3045 520 502 1342 vdd hvtpfet l=6e-08 w=4.11e-07 $X=37059 $Y=20589 $D=636
M3046 521 501 1343 vdd hvtpfet l=6e-08 w=4.11e-07 $X=37059 $Y=22852 $D=636
M3047 522 502 1344 vdd hvtpfet l=6e-08 w=4.11e-07 $X=37059 $Y=27509 $D=636
M3048 b_pxaa<2> 503 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=37150 $Y=1941 $D=636
M3049 503 504 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=37150 $Y=5141 $D=636
M3050 504 505 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=37150 $Y=8691 $D=636
M3051 vdd 497 505 vdd hvtpfet l=6e-08 w=4.11e-07 $X=37150 $Y=10156 $D=636
M3052 vdd 498 506 vdd hvtpfet l=6e-08 w=4.11e-07 $X=37150 $Y=40566 $D=636
M3053 507 506 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=37150 $Y=41842 $D=636
M3054 508 507 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=37150 $Y=44992 $D=636
M3055 t_pxaa<2> 508 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=37150 $Y=46622 $D=636
M3056 776 ddqa_n vdd vdd hvtpfet l=6e-08 w=6.4e-07 $X=37161 $Y=35802 $D=636
M3057 vdd 502 501 vdd hvtpfet l=6e-08 w=4.11e-07 $X=37274 $Y=14280 $D=636
M3058 1345 509 519 vdd hvtpfet l=6e-08 w=4.11e-07 $X=37319 $Y=15932 $D=636
M3059 1346 509 520 vdd hvtpfet l=6e-08 w=4.11e-07 $X=37319 $Y=20589 $D=636
M3060 1347 491 521 vdd hvtpfet l=6e-08 w=4.11e-07 $X=37319 $Y=22852 $D=636
M3061 1348 491 522 vdd hvtpfet l=6e-08 w=4.11e-07 $X=37319 $Y=27509 $D=636
M3062 vdd 503 b_pxaa<2> vdd hvtpfet l=6e-08 w=2.57e-06 $X=37410 $Y=1941 $D=636
M3063 vdd 504 503 vdd hvtpfet l=6e-08 w=1e-06 $X=37410 $Y=5141 $D=636
M3064 vdd 505 504 vdd hvtpfet l=6e-08 w=6e-07 $X=37410 $Y=8691 $D=636
M3065 505 510 vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=37410 $Y=10156 $D=636
M3066 506 510 vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=37410 $Y=40566 $D=636
M3067 vdd 506 507 vdd hvtpfet l=6e-08 w=6e-07 $X=37410 $Y=41842 $D=636
M3068 vdd 507 508 vdd hvtpfet l=6e-08 w=1e-06 $X=37410 $Y=44992 $D=636
M3069 vdd 508 t_pxaa<2> vdd hvtpfet l=6e-08 w=2.57e-06 $X=37410 $Y=46622 $D=636
M3070 493 ddqa 776 vdd hvtpfet l=6e-08 w=6.4e-07 $X=37421 $Y=35802 $D=636
M3071 vdd clka 524 vdd hvtpfet l=6e-08 w=1.2e-06 $X=37485 $Y=29148 $D=636
M3072 vdd 317 1345 vdd hvtpfet l=6e-08 w=8.23e-07 $X=37589 $Y=15520 $D=636
M3073 vdd 317 1346 vdd hvtpfet l=6e-08 w=8.23e-07 $X=37589 $Y=20589 $D=636
M3074 vdd 317 1347 vdd hvtpfet l=6e-08 w=8.23e-07 $X=37589 $Y=22440 $D=636
M3075 vdd 317 1348 vdd hvtpfet l=6e-08 w=8.23e-07 $X=37589 $Y=27509 $D=636
M3076 vdd 496 557 vdd hvtpfet l=6e-08 w=6.4e-07 $X=37661 $Y=33693 $D=636
M3077 502 aa<5> vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=37784 $Y=14280 $D=636
M3078 b_pxaa<1> 512 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=37920 $Y=1941 $D=636
M3079 512 513 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=37920 $Y=5141 $D=636
M3080 513 514 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=37920 $Y=8691 $D=636
M3081 vdd 523 514 vdd hvtpfet l=6e-08 w=4.11e-07 $X=37920 $Y=10156 $D=636
M3082 vdd 523 515 vdd hvtpfet l=6e-08 w=4.11e-07 $X=37920 $Y=40566 $D=636
M3083 516 515 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=37920 $Y=41842 $D=636
M3084 517 516 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=37920 $Y=44992 $D=636
M3085 t_pxaa<1> 517 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=37920 $Y=46622 $D=636
M3086 557 386 vdd vdd hvtpfet l=6e-08 w=6.4e-07 $X=37921 $Y=33693 $D=636
M3087 492 519 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=38099 $Y=15321 $D=636
M3088 1349 323 519 vdd hvtpfet l=6e-08 w=2.74e-07 $X=38099 $Y=16069 $D=636
M3089 1350 323 520 vdd hvtpfet l=6e-08 w=2.74e-07 $X=38099 $Y=20589 $D=636
M3090 510 520 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=38099 $Y=21405 $D=636
M3091 523 521 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=38099 $Y=22241 $D=636
M3092 1351 323 521 vdd hvtpfet l=6e-08 w=2.74e-07 $X=38099 $Y=22989 $D=636
M3093 1352 323 522 vdd hvtpfet l=6e-08 w=2.74e-07 $X=38099 $Y=27509 $D=636
M3094 525 522 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=38099 $Y=28325 $D=636
M3095 vdd 493 526 vdd hvtpfet l=1.4e-07 w=6.4e-07 $X=38141 $Y=36067 $D=636
M3096 vdd 512 b_pxaa<1> vdd hvtpfet l=6e-08 w=2.57e-06 $X=38180 $Y=1941 $D=636
M3097 vdd 513 512 vdd hvtpfet l=6e-08 w=1e-06 $X=38180 $Y=5141 $D=636
M3098 vdd 514 513 vdd hvtpfet l=6e-08 w=6e-07 $X=38180 $Y=8691 $D=636
M3099 514 497 vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=38180 $Y=10156 $D=636
M3100 515 498 vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=38180 $Y=40566 $D=636
M3101 vdd 515 516 vdd hvtpfet l=6e-08 w=6e-07 $X=38180 $Y=41842 $D=636
M3102 vdd 516 517 vdd hvtpfet l=6e-08 w=1e-06 $X=38180 $Y=44992 $D=636
M3103 vdd 517 t_pxaa<1> vdd hvtpfet l=6e-08 w=2.57e-06 $X=38180 $Y=46622 $D=636
M3104 1353 524 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=38255 $Y=29525 $D=636
M3105 vdd 519 492 vdd hvtpfet l=6e-08 w=2.06e-07 $X=38359 $Y=15321 $D=636
M3106 vdd 492 1349 vdd hvtpfet l=6e-08 w=2.74e-07 $X=38359 $Y=16069 $D=636
M3107 vdd 510 1350 vdd hvtpfet l=6e-08 w=2.74e-07 $X=38359 $Y=20589 $D=636
M3108 vdd 520 510 vdd hvtpfet l=6e-08 w=2.06e-07 $X=38359 $Y=21405 $D=636
M3109 vdd 521 523 vdd hvtpfet l=6e-08 w=2.06e-07 $X=38359 $Y=22241 $D=636
M3110 vdd 523 1351 vdd hvtpfet l=6e-08 w=2.74e-07 $X=38359 $Y=22989 $D=636
M3111 vdd 525 1352 vdd hvtpfet l=6e-08 w=2.74e-07 $X=38359 $Y=27509 $D=636
M3112 vdd 522 525 vdd hvtpfet l=6e-08 w=2.06e-07 $X=38359 $Y=28325 $D=636
M3113 779 494 vdd vdd hvtpfet l=6e-08 w=6.4e-07 $X=38431 $Y=33468 $D=636
M3114 780 526 vdd vdd hvtpfet l=1.4e-07 w=6.4e-07 $X=38481 $Y=36067 $D=636
M3115 534 495 1353 vdd hvtpfet l=6e-08 w=8.23e-07 $X=38515 $Y=29525 $D=636
M3116 vdd 533 546 vdd hvtpfet l=6e-08 w=4.11e-07 $X=38574 $Y=14280 $D=636
M3117 b_pxaa<0> 527 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=38690 $Y=1941 $D=636
M3118 527 528 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=38690 $Y=5141 $D=636
M3119 528 529 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=38690 $Y=8691 $D=636
M3120 vdd 497 529 vdd hvtpfet l=6e-08 w=4.11e-07 $X=38690 $Y=10156 $D=636
M3121 vdd 498 530 vdd hvtpfet l=6e-08 w=4.11e-07 $X=38690 $Y=40566 $D=636
M3122 531 530 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=38690 $Y=41842 $D=636
M3123 532 531 vdd vdd hvtpfet l=6e-08 w=1e-06 $X=38690 $Y=44992 $D=636
M3124 t_pxaa<0> 532 vdd vdd hvtpfet l=6e-08 w=2.57e-06 $X=38690 $Y=46622 $D=636
M3125 vdd 527 b_pxaa<0> vdd hvtpfet l=6e-08 w=2.57e-06 $X=38950 $Y=1941 $D=636
M3126 vdd 528 527 vdd hvtpfet l=6e-08 w=1e-06 $X=38950 $Y=5141 $D=636
M3127 vdd 529 528 vdd hvtpfet l=6e-08 w=6e-07 $X=38950 $Y=8691 $D=636
M3128 529 525 vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=38950 $Y=10156 $D=636
M3129 530 525 vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=38950 $Y=40566 $D=636
M3130 vdd 530 531 vdd hvtpfet l=6e-08 w=6e-07 $X=38950 $Y=41842 $D=636
M3131 vdd 531 532 vdd hvtpfet l=6e-08 w=1e-06 $X=38950 $Y=44992 $D=636
M3132 vdd 532 t_pxaa<0> vdd hvtpfet l=6e-08 w=2.57e-06 $X=38950 $Y=46622 $D=636
M3133 1354 534 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=39025 $Y=29525 $D=636
M3134 533 aa<3> vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=39084 $Y=14280 $D=636
M3135 1355 317 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=39109 $Y=15520 $D=636
M3136 1356 317 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=39109 $Y=20589 $D=636
M3137 1357 317 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=39109 $Y=22440 $D=636
M3138 1358 317 vdd vdd hvtpfet l=6e-08 w=8.23e-07 $X=39109 $Y=27509 $D=636
M3139 vdd clka 323 vdd hvtpfet l=6e-08 w=6e-07 $X=39174 $Y=33747 $D=636
M3140 293 535 vdd vdd hvtpfet l=6e-08 w=1.2e-06 $X=39185 $Y=35277 $D=636
M3141 495 539 1354 vdd hvtpfet l=6e-08 w=8.23e-07 $X=39285 $Y=29525 $D=636
M3142 549 537 1355 vdd hvtpfet l=6e-08 w=4.11e-07 $X=39379 $Y=15932 $D=636
M3143 550 538 1356 vdd hvtpfet l=6e-08 w=4.11e-07 $X=39379 $Y=20589 $D=636
M3144 551 537 1357 vdd hvtpfet l=6e-08 w=4.11e-07 $X=39379 $Y=22852 $D=636
M3145 552 538 1358 vdd hvtpfet l=6e-08 w=4.11e-07 $X=39379 $Y=27509 $D=636
M3146 323 clka vdd vdd hvtpfet l=6e-08 w=6e-07 $X=39434 $Y=33747 $D=636
M3147 vdd 538 537 vdd hvtpfet l=6e-08 w=4.11e-07 $X=39594 $Y=14280 $D=636
M3148 1359 546 549 vdd hvtpfet l=6e-08 w=4.11e-07 $X=39639 $Y=15932 $D=636
M3149 1360 546 550 vdd hvtpfet l=6e-08 w=4.11e-07 $X=39639 $Y=20589 $D=636
M3150 1361 533 551 vdd hvtpfet l=6e-08 w=4.11e-07 $X=39639 $Y=22852 $D=636
M3151 1362 533 552 vdd hvtpfet l=6e-08 w=4.11e-07 $X=39639 $Y=27509 $D=636
M3152 vdd clka 323 vdd hvtpfet l=6e-08 w=6e-07 $X=39694 $Y=33747 $D=636
M3153 r_sa_prea_n 293 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=39695 $Y=35277 $D=636
M3154 289 540 vdd vdd hvtpfet l=6e-08 w=1.2e-06 $X=39705 $Y=1736 $D=636
M3155 290 541 vdd vdd hvtpfet l=6e-08 w=1.2e-06 $X=39705 $Y=3566 $D=636
M3156 291 542 vdd vdd hvtpfet l=6e-08 w=1.2e-06 $X=39705 $Y=8196 $D=636
M3157 292 543 vdd vdd hvtpfet l=6e-08 w=1.2e-06 $X=39705 $Y=10026 $D=636
M3158 294 543 vdd vdd hvtpfet l=6e-08 w=1.2e-06 $X=39705 $Y=39907 $D=636
M3159 295 542 vdd vdd hvtpfet l=6e-08 w=1.2e-06 $X=39705 $Y=41737 $D=636
M3160 296 544 vdd vdd hvtpfet l=6e-08 w=1.2e-06 $X=39705 $Y=46367 $D=636
M3161 297 545 vdd vdd hvtpfet l=6e-08 w=1.2e-06 $X=39705 $Y=48197 $D=636
M3162 vdd stclka 539 vdd hvtpfet l=6e-08 w=4.11e-07 $X=39795 $Y=29937 $D=636
M3163 vdd 317 1359 vdd hvtpfet l=6e-08 w=8.23e-07 $X=39909 $Y=15520 $D=636
M3164 vdd 317 1360 vdd hvtpfet l=6e-08 w=8.23e-07 $X=39909 $Y=20589 $D=636
M3165 vdd 317 1361 vdd hvtpfet l=6e-08 w=8.23e-07 $X=39909 $Y=22440 $D=636
M3166 vdd 317 1362 vdd hvtpfet l=6e-08 w=8.23e-07 $X=39909 $Y=27509 $D=636
M3167 323 clka vdd vdd hvtpfet l=6e-08 w=6e-07 $X=39954 $Y=33747 $D=636
M3168 vdd 293 r_sa_prea_n vdd hvtpfet l=6e-08 w=1.43e-06 $X=39955 $Y=35277 $D=636
M3169 538 aa<2> vdd vdd hvtpfet l=6e-08 w=4.11e-07 $X=40104 $Y=14280 $D=636
M3170 rb_ca<1> 289 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=40215 $Y=1506 $D=636
M3171 rb_ca<3> 290 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=40215 $Y=3566 $D=636
M3172 rb_ma<1> 291 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=40215 $Y=7966 $D=636
M3173 rb_ma<3> 292 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=40215 $Y=10026 $D=636
M3174 r_sa_prea_n 293 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=40215 $Y=35277 $D=636
M3175 rt_ma<3> 294 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=40215 $Y=39677 $D=636
M3176 rt_ma<1> 295 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=40215 $Y=41737 $D=636
M3177 rt_ca<3> 296 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=40215 $Y=46137 $D=636
M3178 rt_ca<1> 297 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=40215 $Y=48197 $D=636
M3179 543 549 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=40419 $Y=15321 $D=636
M3180 1363 323 549 vdd hvtpfet l=6e-08 w=2.74e-07 $X=40419 $Y=16069 $D=636
M3181 1364 323 550 vdd hvtpfet l=6e-08 w=2.74e-07 $X=40419 $Y=20589 $D=636
M3182 553 550 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=40419 $Y=21405 $D=636
M3183 542 551 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=40419 $Y=22241 $D=636
M3184 1365 323 551 vdd hvtpfet l=6e-08 w=2.74e-07 $X=40419 $Y=22989 $D=636
M3185 1366 323 552 vdd hvtpfet l=6e-08 w=2.74e-07 $X=40419 $Y=27509 $D=636
M3186 554 552 vdd vdd hvtpfet l=6e-08 w=2.06e-07 $X=40419 $Y=28325 $D=636
M3187 vdd 289 rb_ca<1> vdd hvtpfet l=6e-08 w=1.43e-06 $X=40475 $Y=1506 $D=636
M3188 vdd 290 rb_ca<3> vdd hvtpfet l=6e-08 w=1.43e-06 $X=40475 $Y=3566 $D=636
M3189 vdd 291 rb_ma<1> vdd hvtpfet l=6e-08 w=1.43e-06 $X=40475 $Y=7966 $D=636
M3190 vdd 292 rb_ma<3> vdd hvtpfet l=6e-08 w=1.43e-06 $X=40475 $Y=10026 $D=636
M3191 vdd 294 rt_ma<3> vdd hvtpfet l=6e-08 w=1.43e-06 $X=40475 $Y=39677 $D=636
M3192 vdd 295 rt_ma<1> vdd hvtpfet l=6e-08 w=1.43e-06 $X=40475 $Y=41737 $D=636
M3193 vdd 296 rt_ca<3> vdd hvtpfet l=6e-08 w=1.43e-06 $X=40475 $Y=46137 $D=636
M3194 vdd 297 rt_ca<1> vdd hvtpfet l=6e-08 w=1.43e-06 $X=40475 $Y=48197 $D=636
M3195 vdd 549 543 vdd hvtpfet l=6e-08 w=2.06e-07 $X=40679 $Y=15321 $D=636
M3196 vdd 543 1363 vdd hvtpfet l=6e-08 w=2.74e-07 $X=40679 $Y=16069 $D=636
M3197 vdd 553 1364 vdd hvtpfet l=6e-08 w=2.74e-07 $X=40679 $Y=20589 $D=636
M3198 vdd 550 553 vdd hvtpfet l=6e-08 w=2.06e-07 $X=40679 $Y=21405 $D=636
M3199 vdd 551 542 vdd hvtpfet l=6e-08 w=2.06e-07 $X=40679 $Y=22241 $D=636
M3200 vdd 542 1365 vdd hvtpfet l=6e-08 w=2.74e-07 $X=40679 $Y=22989 $D=636
M3201 vdd 554 1366 vdd hvtpfet l=6e-08 w=2.74e-07 $X=40679 $Y=27509 $D=636
M3202 vdd 552 554 vdd hvtpfet l=6e-08 w=2.06e-07 $X=40679 $Y=28325 $D=636
M3203 vdd 303 r_saea_n vdd hvtpfet l=6e-08 w=1.43e-06 $X=40725 $Y=35277 $D=636
M3204 rb_ca<1> 289 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=40735 $Y=1506 $D=636
M3205 rb_ca<3> 290 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=40735 $Y=3566 $D=636
M3206 rb_ma<1> 291 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=40735 $Y=7966 $D=636
M3207 rb_ma<3> 292 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=40735 $Y=10026 $D=636
M3208 rt_ma<3> 294 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=40735 $Y=39677 $D=636
M3209 rt_ma<1> 295 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=40735 $Y=41737 $D=636
M3210 rt_ca<3> 296 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=40735 $Y=46137 $D=636
M3211 rt_ca<1> 297 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=40735 $Y=48197 $D=636
M3212 r_saea_n 303 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=40985 $Y=35277 $D=636
M3213 vdd 299 rb_ca<0> vdd hvtpfet l=6e-08 w=1.43e-06 $X=41245 $Y=1506 $D=636
M3214 vdd 300 rb_ca<2> vdd hvtpfet l=6e-08 w=1.43e-06 $X=41245 $Y=3566 $D=636
M3215 vdd 301 rb_ma<0> vdd hvtpfet l=6e-08 w=1.43e-06 $X=41245 $Y=7966 $D=636
M3216 vdd 302 rb_ma<2> vdd hvtpfet l=6e-08 w=1.43e-06 $X=41245 $Y=10026 $D=636
M3217 vdd 303 r_saea_n vdd hvtpfet l=6e-08 w=1.43e-06 $X=41245 $Y=35277 $D=636
M3218 vdd 304 rt_ma<2> vdd hvtpfet l=6e-08 w=1.43e-06 $X=41245 $Y=39677 $D=636
M3219 vdd 305 rt_ma<0> vdd hvtpfet l=6e-08 w=1.43e-06 $X=41245 $Y=41737 $D=636
M3220 vdd 306 rt_ca<2> vdd hvtpfet l=6e-08 w=1.43e-06 $X=41245 $Y=46137 $D=636
M3221 vdd 307 rt_ca<0> vdd hvtpfet l=6e-08 w=1.43e-06 $X=41245 $Y=48197 $D=636
M3222 vdd clka 287 vdd hvtpfet l=6e-08 w=2.1e-06 $X=41495 $Y=23621 $D=636
M3223 vdd 340 288 vdd hvtpfet l=6e-08 w=2.1e-06 $X=41495 $Y=26587 $D=636
M3224 rb_ca<0> 299 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=41505 $Y=1506 $D=636
M3225 rb_ca<2> 300 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=41505 $Y=3566 $D=636
M3226 rb_ma<0> 301 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=41505 $Y=7966 $D=636
M3227 rb_ma<2> 302 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=41505 $Y=10026 $D=636
M3228 285 497 vdd vdd hvtpfet l=6e-08 w=1.2e-06 $X=41505 $Y=15067 $D=636
M3229 286 498 vdd vdd hvtpfet l=6e-08 w=1.2e-06 $X=41505 $Y=18424 $D=636
M3230 r_saea_n 303 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=41505 $Y=35277 $D=636
M3231 rt_ma<2> 304 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=41505 $Y=39677 $D=636
M3232 rt_ma<0> 305 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=41505 $Y=41737 $D=636
M3233 rt_ca<2> 306 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=41505 $Y=46137 $D=636
M3234 rt_ca<0> 307 vdd vdd hvtpfet l=6e-08 w=1.43e-06 $X=41505 $Y=48197 $D=636
M3235 r_clk_dqa 287 vdd vdd hvtpfet l=6e-08 w=2.1e-06 $X=41755 $Y=23621 $D=636
M3236 r_clk_dqa_n 288 vdd vdd hvtpfet l=6e-08 w=2.1e-06 $X=41755 $Y=26587 $D=636
M3237 vdd 299 rb_ca<0> vdd hvtpfet l=6e-08 w=1.43e-06 $X=41765 $Y=1506 $D=636
M3238 vdd 300 rb_ca<2> vdd hvtpfet l=6e-08 w=1.43e-06 $X=41765 $Y=3566 $D=636
M3239 vdd 301 rb_ma<0> vdd hvtpfet l=6e-08 w=1.43e-06 $X=41765 $Y=7966 $D=636
M3240 vdd 302 rb_ma<2> vdd hvtpfet l=6e-08 w=1.43e-06 $X=41765 $Y=10026 $D=636
M3241 vdd 303 r_saea_n vdd hvtpfet l=6e-08 w=1.43e-06 $X=41765 $Y=35277 $D=636
M3242 vdd 304 rt_ma<2> vdd hvtpfet l=6e-08 w=1.43e-06 $X=41765 $Y=39677 $D=636
M3243 vdd 305 rt_ma<0> vdd hvtpfet l=6e-08 w=1.43e-06 $X=41765 $Y=41737 $D=636
M3244 vdd 306 rt_ca<2> vdd hvtpfet l=6e-08 w=1.43e-06 $X=41765 $Y=46137 $D=636
M3245 vdd 307 rt_ca<0> vdd hvtpfet l=6e-08 w=1.43e-06 $X=41765 $Y=48197 $D=636
M3246 rb_tm_prea_n 285 vdd vdd hvtpfet l=6e-08 w=2.145e-06 $X=42015 $Y=14887 $D=636
M3247 rt_tm_prea_n 286 vdd vdd hvtpfet l=6e-08 w=2.145e-06 $X=42015 $Y=17659 $D=636
M3248 vdd 287 r_clk_dqa vdd hvtpfet l=6e-08 w=2.1e-06 $X=42015 $Y=23621 $D=636
M3249 vdd 288 r_clk_dqa_n vdd hvtpfet l=6e-08 w=2.1e-06 $X=42015 $Y=26587 $D=636
M3250 r_lwea 284 vdd vdd hvtpfet l=6e-08 w=2.145e-06 $X=42015 $Y=32504 $D=636
M3251 vdd 555 299 vdd hvtpfet l=6e-08 w=1.2e-06 $X=42275 $Y=1736 $D=636
M3252 vdd 556 300 vdd hvtpfet l=6e-08 w=1.2e-06 $X=42275 $Y=3566 $D=636
M3253 vdd 554 301 vdd hvtpfet l=6e-08 w=1.2e-06 $X=42275 $Y=8196 $D=636
M3254 vdd 553 302 vdd hvtpfet l=6e-08 w=1.2e-06 $X=42275 $Y=10026 $D=636
M3255 vdd 285 rb_tm_prea_n vdd hvtpfet l=6e-08 w=2.145e-06 $X=42275 $Y=14887 $D=636
M3256 vdd 286 rt_tm_prea_n vdd hvtpfet l=6e-08 w=2.145e-06 $X=42275 $Y=17659 $D=636
M3257 r_clk_dqa 287 vdd vdd hvtpfet l=6e-08 w=2.1e-06 $X=42275 $Y=23621 $D=636
M3258 r_clk_dqa_n 288 vdd vdd hvtpfet l=6e-08 w=2.1e-06 $X=42275 $Y=26587 $D=636
M3259 vdd 284 r_lwea vdd hvtpfet l=6e-08 w=2.145e-06 $X=42275 $Y=32504 $D=636
M3260 vdd 557 303 vdd hvtpfet l=6e-08 w=1.2e-06 $X=42275 $Y=35277 $D=636
M3261 vdd 553 304 vdd hvtpfet l=6e-08 w=1.2e-06 $X=42275 $Y=39907 $D=636
M3262 vdd 554 305 vdd hvtpfet l=6e-08 w=1.2e-06 $X=42275 $Y=41737 $D=636
M3263 vdd 558 306 vdd hvtpfet l=6e-08 w=1.2e-06 $X=42275 $Y=46367 $D=636
M3264 vdd 559 307 vdd hvtpfet l=6e-08 w=1.2e-06 $X=42275 $Y=48197 $D=636
M3265 303 557 vdd vdd hvtpfet l=6e-08 w=1.2e-06 $X=42535 $Y=35277 $D=636
.ends

************************************************************************
* Library Name: XMC55_DPS
* Cell Name:    xmc55_dps_localc4io_bw
************************************************************************
.SUBCKT xmc55_dps_localc4io_bw b_bla<3> b_bla<2> b_bla<1> b_bla<0> b_bla_n<3> 
+ b_bla_n<2> b_bla_n<1> b_bla_n<0> b_blb<3> b_blb<2> b_blb<1> b_blb<0> 
+ b_blb_n<3> b_blb_n<2> b_blb_n<1> b_blb_n<0> b_ca<3> b_ca<2> b_ca<1> b_ca<0> 
+ b_cb<3> b_cb<2> b_cb<1> b_cb<0> b_ma<3> b_ma<2> b_ma<1> b_ma<0> b_mb<3> 
+ b_mb<2> b_mb<1> b_mb<0> b_tm_prea_n b_tm_preb_n bwena bwenb clk_dqa 
+ clk_dqa_n clk_dqb clk_dqb_n da db ddqa ddqa_n ddqb ddqb_n lwea lweb qa qb 
+ sa_prea_n sa_preb_n saea_n saeb_n t_bla<3> t_bla<2> t_bla<1> t_bla<0> 
+ t_bla_n<3> t_bla_n<2> t_bla_n<1> t_bla_n<0> t_blb<3> t_blb<2> t_blb<1> 
+ t_blb<0> t_blb_n<3> t_blb_n<2> t_blb_n<1> t_blb_n<0> t_ca<3> t_ca<2> t_ca<1> 
+ t_ca<0> t_cb<3> t_cb<2> t_cb<1> t_cb<0> t_ma<3> t_ma<2> t_ma<1> t_ma<0> 
+ t_mb<3> t_mb<2> t_mb<1> t_mb<0> t_tm_prea_n t_tm_preb_n vdd vss
** N=5219 EP=90 IP=0 FDC=654
M0 143 11 b_blb<3> vss hvtnfet l=6e-08 w=6e-07 $X=210 $Y=2941 $D=616
M1 143 11 b_blb<3> vss hvtnfet l=6e-08 w=6e-07 $X=210 $Y=3201 $D=616
M2 148 24 b_bla_n<3> vss hvtnfet l=6e-08 w=6e-07 $X=210 $Y=3881 $D=616
M3 148 24 b_bla_n<3> vss hvtnfet l=6e-08 w=6e-07 $X=210 $Y=4141 $D=616
M4 t_bla_n<3> 25 148 vss hvtnfet l=6e-08 w=6e-07 $X=210 $Y=46932 $D=616
M5 148 25 t_bla_n<3> vss hvtnfet l=6e-08 w=6e-07 $X=210 $Y=47192 $D=616
M6 t_blb<3> 12 143 vss hvtnfet l=6e-08 w=6e-07 $X=210 $Y=47872 $D=616
M7 143 12 t_blb<3> vss hvtnfet l=6e-08 w=6e-07 $X=210 $Y=48132 $D=616
M8 148 23 vss vss hvtnfet l=6e-08 w=6e-07 $X=423 $Y=26159 $D=616
M9 11 5 vss vss hvtnfet l=6e-08 w=4e-07 $X=535 $Y=4836 $D=616
M10 311 b_cb<3> 5 vss hvtnfet l=6e-08 w=4e-07 $X=535 $Y=11331 $D=616
M11 312 5 2 vss hvtnfet l=6e-08 w=4e-07 $X=535 $Y=12191 $D=616
M12 313 6 3 vss hvtnfet l=6e-08 w=4e-07 $X=535 $Y=38542 $D=616
M13 314 t_cb<3> 6 vss hvtnfet l=6e-08 w=4e-07 $X=535 $Y=39402 $D=616
M14 12 6 vss vss hvtnfet l=6e-08 w=4e-07 $X=535 $Y=45897 $D=616
M15 vss vdd 152 vss hvtnfet l=6e-08 w=3e-07 $X=573 $Y=31223 $D=616
M16 vss bwena 26 vss hvtnfet l=1.4e-07 w=2.1e-07 $X=605 $Y=14555 $D=616
M17 vss 13 43 vss hvtnfet l=1.4e-07 w=2.1e-07 $X=605 $Y=16755 $D=616
M18 vss 14 ddqa_n vss hvtnfet l=7e-08 w=3.2e-07 $X=610 $Y=33798 $D=616
M19 174 vdd vss vss hvtnfet l=6e-08 w=3e-07 $X=630 $Y=17670 $D=616
M20 14 16 196 vss hvtnfet l=1.4e-07 w=7.5e-07 $X=650 $Y=34593 $D=616
M21 vss 23 148 vss hvtnfet l=6e-08 w=6e-07 $X=683 $Y=26159 $D=616
M22 vss 18 11 vss hvtnfet l=6e-08 w=4e-07 $X=795 $Y=4836 $D=616
M23 vss b_mb<0> 311 vss hvtnfet l=6e-08 w=4e-07 $X=795 $Y=11331 $D=616
M24 vss 20 312 vss hvtnfet l=6e-08 w=4e-07 $X=795 $Y=12191 $D=616
M25 vss 21 313 vss hvtnfet l=6e-08 w=4e-07 $X=795 $Y=38542 $D=616
M26 vss t_mb<0> 314 vss hvtnfet l=6e-08 w=4e-07 $X=795 $Y=39402 $D=616
M27 vss 18 12 vss hvtnfet l=6e-08 w=4e-07 $X=795 $Y=45897 $D=616
M28 vss vdd 174 vss hvtnfet l=6e-08 w=3e-07 $X=890 $Y=17670 $D=616
M29 196 17 vss vss hvtnfet l=8e-08 w=3.75e-07 $X=890 $Y=33798 $D=616
M30 39 26 vss vss hvtnfet l=1.4e-07 w=2.1e-07 $X=945 $Y=14555 $D=616
M31 13 42 vss vss hvtnfet l=1.4e-07 w=2.1e-07 $X=945 $Y=16755 $D=616
M32 196 16 14 vss hvtnfet l=1.4e-07 w=7.5e-07 $X=990 $Y=34593 $D=616
M33 24 29 vss vss hvtnfet l=6e-08 w=4e-07 $X=1055 $Y=4836 $D=616
M34 315 b_ma<0> vss vss hvtnfet l=6e-08 w=4e-07 $X=1055 $Y=11331 $D=616
M35 316 31 vss vss hvtnfet l=6e-08 w=4e-07 $X=1055 $Y=12191 $D=616
M36 317 32 vss vss hvtnfet l=6e-08 w=4e-07 $X=1055 $Y=38542 $D=616
M37 318 t_ma<0> vss vss hvtnfet l=6e-08 w=4e-07 $X=1055 $Y=39402 $D=616
M38 25 29 vss vss hvtnfet l=6e-08 w=4e-07 $X=1055 $Y=45897 $D=616
M39 319 17 vss vss hvtnfet l=6e-08 w=3e-07 $X=1083 $Y=31223 $D=616
M40 159 11 b_blb_n<3> vss hvtnfet l=6e-08 w=6e-07 $X=1100 $Y=2941 $D=616
M41 159 11 b_blb_n<3> vss hvtnfet l=6e-08 w=6e-07 $X=1100 $Y=3201 $D=616
M42 b_bla<3> 24 169 vss hvtnfet l=6e-08 w=6e-07 $X=1100 $Y=3881 $D=616
M43 b_bla<3> 24 169 vss hvtnfet l=6e-08 w=6e-07 $X=1100 $Y=4141 $D=616
M44 169 25 t_bla<3> vss hvtnfet l=6e-08 w=6e-07 $X=1100 $Y=46932 $D=616
M45 t_bla<3> 25 169 vss hvtnfet l=6e-08 w=6e-07 $X=1100 $Y=47192 $D=616
M46 t_blb_n<3> 12 159 vss hvtnfet l=6e-08 w=6e-07 $X=1100 $Y=47872 $D=616
M47 159 12 t_blb_n<3> vss hvtnfet l=6e-08 w=6e-07 $X=1100 $Y=48132 $D=616
M48 174 vdd vss vss hvtnfet l=6e-08 w=3e-07 $X=1150 $Y=17670 $D=616
M49 vss 17 196 vss hvtnfet l=8e-08 w=3.75e-07 $X=1170 $Y=33798 $D=616
M50 vss 35 179 vss hvtnfet l=6e-08 w=8e-07 $X=1193 $Y=26159 $D=616
M51 49 14 319 vss hvtnfet l=6e-08 w=3e-07 $X=1273 $Y=31223 $D=616
M52 vss 27 24 vss hvtnfet l=6e-08 w=4e-07 $X=1315 $Y=4836 $D=616
M53 27 b_ca<3> 315 vss hvtnfet l=6e-08 w=4e-07 $X=1315 $Y=11331 $D=616
M54 36 27 316 vss hvtnfet l=6e-08 w=4e-07 $X=1315 $Y=12191 $D=616
M55 37 28 317 vss hvtnfet l=6e-08 w=4e-07 $X=1315 $Y=38542 $D=616
M56 28 t_ca<3> 318 vss hvtnfet l=6e-08 w=4e-07 $X=1315 $Y=39402 $D=616
M57 vss 28 25 vss hvtnfet l=6e-08 w=4e-07 $X=1315 $Y=45897 $D=616
M58 16 14 196 vss hvtnfet l=1.4e-07 w=7.5e-07 $X=1330 $Y=34593 $D=616
M59 vss vdd 174 vss hvtnfet l=6e-08 w=3e-07 $X=1410 $Y=17670 $D=616
M60 196 17 vss vss hvtnfet l=8e-08 w=3.75e-07 $X=1450 $Y=33798 $D=616
M61 179 35 vss vss hvtnfet l=6e-08 w=8e-07 $X=1453 $Y=26159 $D=616
M62 320 34 49 vss hvtnfet l=6e-08 w=3e-07 $X=1533 $Y=31223 $D=616
M63 vss 39 52 vss hvtnfet l=1.4e-07 w=2.1e-07 $X=1535 $Y=14555 $D=616
M64 vss 47 42 vss hvtnfet l=1.4e-07 w=2.1e-07 $X=1535 $Y=16755 $D=616
M65 qa 34 vss vss hvtnfet l=6e-08 w=4.5e-07 $X=1615 $Y=19812 $D=616
M66 vss 34 qa vss hvtnfet l=6e-08 w=4.5e-07 $X=1615 $Y=20072 $D=616
M67 321 43 vss vss hvtnfet l=6e-08 w=3.2e-07 $X=1615 $Y=21012 $D=616
M68 321 38 40 vss hvtnfet l=6e-08 w=3.2e-07 $X=1615 $Y=21202 $D=616
M69 322 10 40 vss hvtnfet l=6e-08 w=1.4e-07 $X=1615 $Y=21477 $D=616
M70 vss 8 322 vss hvtnfet l=6e-08 w=1.4e-07 $X=1615 $Y=21667 $D=616
M71 10 40 vss vss hvtnfet l=6e-08 w=2.1e-07 $X=1615 $Y=21942 $D=616
M72 vss 40 23 vss hvtnfet l=6e-08 w=3.2e-07 $X=1615 $Y=22762 $D=616
M73 323 44 vss vss hvtnfet l=6e-08 w=3.2e-07 $X=1615 $Y=23729 $D=616
M74 323 38 41 vss hvtnfet l=6e-08 w=3.2e-07 $X=1615 $Y=23919 $D=616
M75 324 9 41 vss hvtnfet l=6e-08 w=1.4e-07 $X=1615 $Y=24194 $D=616
M76 vss 8 324 vss hvtnfet l=6e-08 w=1.4e-07 $X=1615 $Y=24384 $D=616
M77 9 41 vss vss hvtnfet l=6e-08 w=2.1e-07 $X=1615 $Y=24659 $D=616
M78 174 vdd vss vss hvtnfet l=6e-08 w=3e-07 $X=1670 $Y=17670 $D=616
M79 196 14 16 vss hvtnfet l=1.4e-07 w=7.5e-07 $X=1670 $Y=34593 $D=616
M80 29 lwea 179 vss hvtnfet l=6e-08 w=8e-07 $X=1713 $Y=26159 $D=616
M81 vss saea_n 320 vss hvtnfet l=6e-08 w=3e-07 $X=1723 $Y=31223 $D=616
M82 vss 17 196 vss hvtnfet l=8e-08 w=3.75e-07 $X=1730 $Y=33798 $D=616
M83 44 52 vss vss hvtnfet l=1.4e-07 w=2.1e-07 $X=1875 $Y=14555 $D=616
M84 47 da vss vss hvtnfet l=1.4e-07 w=2.1e-07 $X=1875 $Y=16755 $D=616
M85 vss vdd 174 vss hvtnfet l=6e-08 w=3e-07 $X=1930 $Y=17670 $D=616
M86 179 lwea 29 vss hvtnfet l=6e-08 w=8e-07 $X=1973 $Y=26159 $D=616
M87 196 17 vss vss hvtnfet l=8e-08 w=3.75e-07 $X=2010 $Y=33798 $D=616
M88 14 16 196 vss hvtnfet l=1.4e-07 w=7.5e-07 $X=2010 $Y=34593 $D=616
M89 159 68 b_blb_n<2> vss hvtnfet l=6e-08 w=6e-07 $X=2120 $Y=2941 $D=616
M90 159 68 b_blb_n<2> vss hvtnfet l=6e-08 w=6e-07 $X=2120 $Y=3201 $D=616
M91 b_bla<2> 61 169 vss hvtnfet l=6e-08 w=6e-07 $X=2120 $Y=3881 $D=616
M92 b_bla<2> 61 169 vss hvtnfet l=6e-08 w=6e-07 $X=2120 $Y=4141 $D=616
M93 169 62 t_bla<2> vss hvtnfet l=6e-08 w=6e-07 $X=2120 $Y=46932 $D=616
M94 t_bla<2> 62 169 vss hvtnfet l=6e-08 w=6e-07 $X=2120 $Y=47192 $D=616
M95 t_blb_n<2> 69 159 vss hvtnfet l=6e-08 w=6e-07 $X=2120 $Y=47872 $D=616
M96 159 69 t_blb_n<2> vss hvtnfet l=6e-08 w=6e-07 $X=2120 $Y=48132 $D=616
M97 vss 17 196 vss hvtnfet l=8e-08 w=3.75e-07 $X=2290 $Y=33798 $D=616
M98 196 16 14 vss hvtnfet l=1.4e-07 w=7.5e-07 $X=2350 $Y=34593 $D=616
M99 31 b_tm_prea_n vss vss hvtnfet l=6e-08 w=2.5e-07 $X=2440 $Y=17720 $D=616
M100 61 55 vss vss hvtnfet l=6e-08 w=4e-07 $X=2445 $Y=4836 $D=616
M101 325 b_ca<2> 55 vss hvtnfet l=6e-08 w=4e-07 $X=2445 $Y=11331 $D=616
M102 326 55 58 vss hvtnfet l=6e-08 w=4e-07 $X=2445 $Y=12191 $D=616
M103 327 56 59 vss hvtnfet l=6e-08 w=4e-07 $X=2445 $Y=38542 $D=616
M104 328 t_ca<2> 56 vss hvtnfet l=6e-08 w=4e-07 $X=2445 $Y=39402 $D=616
M105 62 56 vss vss hvtnfet l=6e-08 w=4e-07 $X=2445 $Y=45897 $D=616
M106 169 40 vss vss hvtnfet l=6e-08 w=6e-07 $X=2493 $Y=26159 $D=616
M107 196 17 vss vss hvtnfet l=8e-08 w=3.75e-07 $X=2570 $Y=33798 $D=616
M108 vss 49 34 vss hvtnfet l=6e-08 w=3e-07 $X=2633 $Y=31223 $D=616
M109 38 clk_dqa vss vss hvtnfet l=6e-08 w=2e-07 $X=2645 $Y=21427 $D=616
M110 8 clk_dqa_n vss vss hvtnfet l=6e-08 w=2e-07 $X=2645 $Y=23694 $D=616
M111 65 41 vss vss hvtnfet l=6e-08 w=2e-07 $X=2645 $Y=24394 $D=616
M112 35 65 vss vss hvtnfet l=6e-08 w=2e-07 $X=2645 $Y=24904 $D=616
M113 16 14 196 vss hvtnfet l=1.4e-07 w=7.5e-07 $X=2690 $Y=34593 $D=616
M114 vss b_tm_prea_n 31 vss hvtnfet l=6e-08 w=2.5e-07 $X=2700 $Y=17720 $D=616
M115 vss 29 61 vss hvtnfet l=6e-08 w=4e-07 $X=2705 $Y=4836 $D=616
M116 vss b_ma<0> 325 vss hvtnfet l=6e-08 w=4e-07 $X=2705 $Y=11331 $D=616
M117 vss 31 326 vss hvtnfet l=6e-08 w=4e-07 $X=2705 $Y=12191 $D=616
M118 vss 32 327 vss hvtnfet l=6e-08 w=4e-07 $X=2705 $Y=38542 $D=616
M119 vss t_ma<0> 328 vss hvtnfet l=6e-08 w=4e-07 $X=2705 $Y=39402 $D=616
M120 vss 29 62 vss hvtnfet l=6e-08 w=4e-07 $X=2705 $Y=45897 $D=616
M121 vss 40 169 vss hvtnfet l=6e-08 w=6e-07 $X=2753 $Y=26159 $D=616
M122 vss 17 196 vss hvtnfet l=8e-08 w=3.75e-07 $X=2850 $Y=33798 $D=616
M123 17 saea_n vss vss hvtnfet l=6e-08 w=3e-07 $X=2893 $Y=31223 $D=616
M124 32 t_tm_prea_n vss vss hvtnfet l=6e-08 w=2.5e-07 $X=2960 $Y=17720 $D=616
M125 68 18 vss vss hvtnfet l=6e-08 w=4e-07 $X=2965 $Y=4836 $D=616
M126 329 b_mb<0> vss vss hvtnfet l=6e-08 w=4e-07 $X=2965 $Y=11331 $D=616
M127 330 20 vss vss hvtnfet l=6e-08 w=4e-07 $X=2965 $Y=12191 $D=616
M128 331 21 vss vss hvtnfet l=6e-08 w=4e-07 $X=2965 $Y=38542 $D=616
M129 332 t_mb<0> vss vss hvtnfet l=6e-08 w=4e-07 $X=2965 $Y=39402 $D=616
M130 69 18 vss vss hvtnfet l=6e-08 w=4e-07 $X=2965 $Y=45897 $D=616
M131 143 68 b_blb<2> vss hvtnfet l=6e-08 w=6e-07 $X=3010 $Y=2941 $D=616
M132 143 68 b_blb<2> vss hvtnfet l=6e-08 w=6e-07 $X=3010 $Y=3201 $D=616
M133 148 61 b_bla_n<2> vss hvtnfet l=6e-08 w=6e-07 $X=3010 $Y=3881 $D=616
M134 148 61 b_bla_n<2> vss hvtnfet l=6e-08 w=6e-07 $X=3010 $Y=4141 $D=616
M135 t_bla_n<2> 62 148 vss hvtnfet l=6e-08 w=6e-07 $X=3010 $Y=46932 $D=616
M136 148 62 t_bla_n<2> vss hvtnfet l=6e-08 w=6e-07 $X=3010 $Y=47192 $D=616
M137 t_blb<2> 69 143 vss hvtnfet l=6e-08 w=6e-07 $X=3010 $Y=47872 $D=616
M138 143 69 t_blb<2> vss hvtnfet l=6e-08 w=6e-07 $X=3010 $Y=48132 $D=616
M139 196 14 16 vss hvtnfet l=1.4e-07 w=7.5e-07 $X=3030 $Y=34593 $D=616
M140 ddqa 16 vss vss hvtnfet l=7e-08 w=3.2e-07 $X=3140 $Y=33798 $D=616
M141 vss t_tm_prea_n 32 vss hvtnfet l=6e-08 w=2.5e-07 $X=3220 $Y=17720 $D=616
M142 vss 66 68 vss hvtnfet l=6e-08 w=4e-07 $X=3225 $Y=4836 $D=616
M143 66 b_cb<2> 329 vss hvtnfet l=6e-08 w=4e-07 $X=3225 $Y=11331 $D=616
M144 70 66 330 vss hvtnfet l=6e-08 w=4e-07 $X=3225 $Y=12191 $D=616
M145 71 67 331 vss hvtnfet l=6e-08 w=4e-07 $X=3225 $Y=38542 $D=616
M146 67 t_cb<2> 332 vss hvtnfet l=6e-08 w=4e-07 $X=3225 $Y=39402 $D=616
M147 vss 67 69 vss hvtnfet l=6e-08 w=4e-07 $X=3225 $Y=45897 $D=616
M148 202 16 vss vss hvtnfet l=6e-08 w=3e-07 $X=3403 $Y=31223 $D=616
M149 143 83 b_blb<1> vss hvtnfet l=6e-08 w=6e-07 $X=4030 $Y=2941 $D=616
M150 143 83 b_blb<1> vss hvtnfet l=6e-08 w=6e-07 $X=4030 $Y=3201 $D=616
M151 148 91 b_bla_n<1> vss hvtnfet l=6e-08 w=6e-07 $X=4030 $Y=3881 $D=616
M152 148 91 b_bla_n<1> vss hvtnfet l=6e-08 w=6e-07 $X=4030 $Y=4141 $D=616
M153 t_bla_n<1> 92 148 vss hvtnfet l=6e-08 w=6e-07 $X=4030 $Y=46932 $D=616
M154 148 92 t_bla_n<1> vss hvtnfet l=6e-08 w=6e-07 $X=4030 $Y=47192 $D=616
M155 t_blb<1> 84 143 vss hvtnfet l=6e-08 w=6e-07 $X=4030 $Y=47872 $D=616
M156 143 84 t_blb<1> vss hvtnfet l=6e-08 w=6e-07 $X=4030 $Y=48132 $D=616
M157 vss 75 209 vss hvtnfet l=6e-08 w=3e-07 $X=4177 $Y=31223 $D=616
M158 83 79 vss vss hvtnfet l=6e-08 w=4e-07 $X=4355 $Y=4836 $D=616
M159 333 b_cb<1> 79 vss hvtnfet l=6e-08 w=4e-07 $X=4355 $Y=11331 $D=616
M160 334 79 76 vss hvtnfet l=6e-08 w=4e-07 $X=4355 $Y=12191 $D=616
M161 335 80 77 vss hvtnfet l=6e-08 w=4e-07 $X=4355 $Y=38542 $D=616
M162 336 t_cb<1> 80 vss hvtnfet l=6e-08 w=4e-07 $X=4355 $Y=39402 $D=616
M163 84 80 vss vss hvtnfet l=6e-08 w=4e-07 $X=4355 $Y=45897 $D=616
M164 21 t_tm_preb_n vss vss hvtnfet l=6e-08 w=2.5e-07 $X=4360 $Y=17720 $D=616
M165 vss 75 ddqb vss hvtnfet l=7e-08 w=3.2e-07 $X=4430 $Y=33798 $D=616
M166 75 85 252 vss hvtnfet l=1.4e-07 w=7.5e-07 $X=4470 $Y=34593 $D=616
M167 vss 18 83 vss hvtnfet l=6e-08 w=4e-07 $X=4615 $Y=4836 $D=616
M168 vss b_mb<0> 333 vss hvtnfet l=6e-08 w=4e-07 $X=4615 $Y=11331 $D=616
M169 vss 20 334 vss hvtnfet l=6e-08 w=4e-07 $X=4615 $Y=12191 $D=616
M170 vss 21 335 vss hvtnfet l=6e-08 w=4e-07 $X=4615 $Y=38542 $D=616
M171 vss t_mb<0> 336 vss hvtnfet l=6e-08 w=4e-07 $X=4615 $Y=39402 $D=616
M172 vss 18 84 vss hvtnfet l=6e-08 w=4e-07 $X=4615 $Y=45897 $D=616
M173 vss t_tm_preb_n 21 vss hvtnfet l=6e-08 w=2.5e-07 $X=4620 $Y=17720 $D=616
M174 vss saeb_n 86 vss hvtnfet l=6e-08 w=3e-07 $X=4687 $Y=31223 $D=616
M175 252 86 vss vss hvtnfet l=8e-08 w=3.75e-07 $X=4710 $Y=33798 $D=616
M176 107 clk_dqb vss vss hvtnfet l=6e-08 w=2e-07 $X=4795 $Y=21427 $D=616
M177 105 clk_dqb_n vss vss hvtnfet l=6e-08 w=2e-07 $X=4795 $Y=23694 $D=616
M178 89 88 vss vss hvtnfet l=6e-08 w=2e-07 $X=4795 $Y=24394 $D=616
M179 117 89 vss vss hvtnfet l=6e-08 w=2e-07 $X=4795 $Y=24904 $D=616
M180 252 85 75 vss hvtnfet l=1.4e-07 w=7.5e-07 $X=4810 $Y=34593 $D=616
M181 143 93 vss vss hvtnfet l=6e-08 w=6e-07 $X=4827 $Y=26159 $D=616
M182 91 29 vss vss hvtnfet l=6e-08 w=4e-07 $X=4875 $Y=4836 $D=616
M183 337 b_ma<0> vss vss hvtnfet l=6e-08 w=4e-07 $X=4875 $Y=11331 $D=616
M184 338 31 vss vss hvtnfet l=6e-08 w=4e-07 $X=4875 $Y=12191 $D=616
M185 339 32 vss vss hvtnfet l=6e-08 w=4e-07 $X=4875 $Y=38542 $D=616
M186 340 t_ma<0> vss vss hvtnfet l=6e-08 w=4e-07 $X=4875 $Y=39402 $D=616
M187 92 29 vss vss hvtnfet l=6e-08 w=4e-07 $X=4875 $Y=45897 $D=616
M188 20 b_tm_preb_n vss vss hvtnfet l=6e-08 w=2.5e-07 $X=4880 $Y=17720 $D=616
M189 159 83 b_blb_n<1> vss hvtnfet l=6e-08 w=6e-07 $X=4920 $Y=2941 $D=616
M190 159 83 b_blb_n<1> vss hvtnfet l=6e-08 w=6e-07 $X=4920 $Y=3201 $D=616
M191 b_bla<1> 91 169 vss hvtnfet l=6e-08 w=6e-07 $X=4920 $Y=3881 $D=616
M192 b_bla<1> 91 169 vss hvtnfet l=6e-08 w=6e-07 $X=4920 $Y=4141 $D=616
M193 169 92 t_bla<1> vss hvtnfet l=6e-08 w=6e-07 $X=4920 $Y=46932 $D=616
M194 t_bla<1> 92 169 vss hvtnfet l=6e-08 w=6e-07 $X=4920 $Y=47192 $D=616
M195 t_blb_n<1> 84 159 vss hvtnfet l=6e-08 w=6e-07 $X=4920 $Y=47872 $D=616
M196 159 84 t_blb_n<1> vss hvtnfet l=6e-08 w=6e-07 $X=4920 $Y=48132 $D=616
M197 104 109 vss vss hvtnfet l=6e-08 w=3e-07 $X=4947 $Y=31223 $D=616
M198 vss 86 252 vss hvtnfet l=8e-08 w=3.75e-07 $X=4990 $Y=33798 $D=616
M199 vss 93 143 vss hvtnfet l=6e-08 w=6e-07 $X=5087 $Y=26159 $D=616
M200 vss 94 91 vss hvtnfet l=6e-08 w=4e-07 $X=5135 $Y=4836 $D=616
M201 94 b_ca<1> 337 vss hvtnfet l=6e-08 w=4e-07 $X=5135 $Y=11331 $D=616
M202 97 94 338 vss hvtnfet l=6e-08 w=4e-07 $X=5135 $Y=12191 $D=616
M203 98 95 339 vss hvtnfet l=6e-08 w=4e-07 $X=5135 $Y=38542 $D=616
M204 95 t_ca<1> 340 vss hvtnfet l=6e-08 w=4e-07 $X=5135 $Y=39402 $D=616
M205 vss 95 92 vss hvtnfet l=6e-08 w=4e-07 $X=5135 $Y=45897 $D=616
M206 vss b_tm_preb_n 20 vss hvtnfet l=6e-08 w=2.5e-07 $X=5140 $Y=17720 $D=616
M207 85 75 252 vss hvtnfet l=1.4e-07 w=7.5e-07 $X=5150 $Y=34593 $D=616
M208 252 86 vss vss hvtnfet l=8e-08 w=3.75e-07 $X=5270 $Y=33798 $D=616
M209 252 75 85 vss hvtnfet l=1.4e-07 w=7.5e-07 $X=5490 $Y=34593 $D=616
M210 vss 86 252 vss hvtnfet l=8e-08 w=3.75e-07 $X=5550 $Y=33798 $D=616
M211 qb 104 vss vss hvtnfet l=6e-08 w=4.5e-07 $X=5575 $Y=19812 $D=616
M212 vss 104 qb vss hvtnfet l=6e-08 w=4.5e-07 $X=5575 $Y=20072 $D=616
M213 18 lweb 240 vss hvtnfet l=6e-08 w=8e-07 $X=5607 $Y=26159 $D=616
M214 vss 106 119 vss hvtnfet l=1.4e-07 w=2.1e-07 $X=5625 $Y=14555 $D=616
M215 vss db 110 vss hvtnfet l=1.4e-07 w=2.1e-07 $X=5625 $Y=16755 $D=616
M216 245 vdd vss vss hvtnfet l=6e-08 w=3e-07 $X=5650 $Y=17670 $D=616
M217 341 118 vss vss hvtnfet l=6e-08 w=3.2e-07 $X=5705 $Y=21012 $D=616
M218 341 107 93 vss hvtnfet l=6e-08 w=3.2e-07 $X=5705 $Y=21202 $D=616
M219 vss 93 125 vss hvtnfet l=6e-08 w=3.2e-07 $X=5705 $Y=22762 $D=616
M220 342 119 vss vss hvtnfet l=6e-08 w=3.2e-07 $X=5705 $Y=23729 $D=616
M221 342 107 88 vss hvtnfet l=6e-08 w=3.2e-07 $X=5705 $Y=23919 $D=616
M222 134 93 vss vss hvtnfet l=6e-08 w=2.1e-07 $X=5815 $Y=21942 $D=616
M223 137 88 vss vss hvtnfet l=6e-08 w=2.1e-07 $X=5815 $Y=24659 $D=616
M224 252 86 vss vss hvtnfet l=8e-08 w=3.75e-07 $X=5830 $Y=33798 $D=616
M225 75 85 252 vss hvtnfet l=1.4e-07 w=7.5e-07 $X=5830 $Y=34593 $D=616
M226 345 saeb_n vss vss hvtnfet l=6e-08 w=3e-07 $X=5857 $Y=31223 $D=616
M227 240 lweb 18 vss hvtnfet l=6e-08 w=8e-07 $X=5867 $Y=26159 $D=616
M228 343 134 93 vss hvtnfet l=6e-08 w=1.4e-07 $X=5885 $Y=21477 $D=616
M229 vss 105 343 vss hvtnfet l=6e-08 w=1.4e-07 $X=5885 $Y=21667 $D=616
M230 344 137 88 vss hvtnfet l=6e-08 w=1.4e-07 $X=5885 $Y=24194 $D=616
M231 vss 105 344 vss hvtnfet l=6e-08 w=1.4e-07 $X=5885 $Y=24384 $D=616
M232 vss vdd 245 vss hvtnfet l=6e-08 w=3e-07 $X=5910 $Y=17670 $D=616
M233 159 128 b_blb_n<0> vss hvtnfet l=6e-08 w=6e-07 $X=5940 $Y=2941 $D=616
M234 159 128 b_blb_n<0> vss hvtnfet l=6e-08 w=6e-07 $X=5940 $Y=3201 $D=616
M235 b_bla<0> 122 169 vss hvtnfet l=6e-08 w=6e-07 $X=5940 $Y=3881 $D=616
M236 b_bla<0> 122 169 vss hvtnfet l=6e-08 w=6e-07 $X=5940 $Y=4141 $D=616
M237 169 123 t_bla<0> vss hvtnfet l=6e-08 w=6e-07 $X=5940 $Y=46932 $D=616
M238 t_bla<0> 123 169 vss hvtnfet l=6e-08 w=6e-07 $X=5940 $Y=47192 $D=616
M239 t_blb_n<0> 129 159 vss hvtnfet l=6e-08 w=6e-07 $X=5940 $Y=47872 $D=616
M240 159 129 t_blb_n<0> vss hvtnfet l=6e-08 w=6e-07 $X=5940 $Y=48132 $D=616
M241 106 121 vss vss hvtnfet l=1.4e-07 w=2.1e-07 $X=5965 $Y=14555 $D=616
M242 120 110 vss vss hvtnfet l=1.4e-07 w=2.1e-07 $X=5965 $Y=16755 $D=616
M243 109 104 345 vss hvtnfet l=6e-08 w=3e-07 $X=6047 $Y=31223 $D=616
M244 vss 86 252 vss hvtnfet l=8e-08 w=3.75e-07 $X=6110 $Y=33798 $D=616
M245 vss 117 240 vss hvtnfet l=6e-08 w=8e-07 $X=6127 $Y=26159 $D=616
M246 245 vdd vss vss hvtnfet l=6e-08 w=3e-07 $X=6170 $Y=17670 $D=616
M247 252 85 75 vss hvtnfet l=1.4e-07 w=7.5e-07 $X=6170 $Y=34593 $D=616
M248 122 112 vss vss hvtnfet l=6e-08 w=4e-07 $X=6265 $Y=4836 $D=616
M249 346 b_ca<0> 112 vss hvtnfet l=6e-08 w=4e-07 $X=6265 $Y=11331 $D=616
M250 347 112 115 vss hvtnfet l=6e-08 w=4e-07 $X=6265 $Y=12191 $D=616
M251 348 113 116 vss hvtnfet l=6e-08 w=4e-07 $X=6265 $Y=38542 $D=616
M252 349 t_ca<0> 113 vss hvtnfet l=6e-08 w=4e-07 $X=6265 $Y=39402 $D=616
M253 123 113 vss vss hvtnfet l=6e-08 w=4e-07 $X=6265 $Y=45897 $D=616
M254 350 85 109 vss hvtnfet l=6e-08 w=3e-07 $X=6307 $Y=31223 $D=616
M255 240 117 vss vss hvtnfet l=6e-08 w=8e-07 $X=6387 $Y=26159 $D=616
M256 252 86 vss vss hvtnfet l=8e-08 w=3.75e-07 $X=6390 $Y=33798 $D=616
M257 vss vdd 245 vss hvtnfet l=6e-08 w=3e-07 $X=6430 $Y=17670 $D=616
M258 vss 86 350 vss hvtnfet l=6e-08 w=3e-07 $X=6497 $Y=31223 $D=616
M259 85 75 252 vss hvtnfet l=1.4e-07 w=7.5e-07 $X=6510 $Y=34593 $D=616
M260 vss 29 122 vss hvtnfet l=6e-08 w=4e-07 $X=6525 $Y=4836 $D=616
M261 vss b_ma<0> 346 vss hvtnfet l=6e-08 w=4e-07 $X=6525 $Y=11331 $D=616
M262 vss 31 347 vss hvtnfet l=6e-08 w=4e-07 $X=6525 $Y=12191 $D=616
M263 vss 32 348 vss hvtnfet l=6e-08 w=4e-07 $X=6525 $Y=38542 $D=616
M264 vss t_ma<0> 349 vss hvtnfet l=6e-08 w=4e-07 $X=6525 $Y=39402 $D=616
M265 vss 29 123 vss hvtnfet l=6e-08 w=4e-07 $X=6525 $Y=45897 $D=616
M266 vss 124 121 vss hvtnfet l=1.4e-07 w=2.1e-07 $X=6555 $Y=14555 $D=616
M267 vss 120 133 vss hvtnfet l=1.4e-07 w=2.1e-07 $X=6555 $Y=16755 $D=616
M268 vss 86 252 vss hvtnfet l=8e-08 w=3.75e-07 $X=6670 $Y=33798 $D=616
M269 245 vdd vss vss hvtnfet l=6e-08 w=3e-07 $X=6690 $Y=17670 $D=616
M270 128 18 vss vss hvtnfet l=6e-08 w=4e-07 $X=6785 $Y=4836 $D=616
M271 351 b_mb<0> vss vss hvtnfet l=6e-08 w=4e-07 $X=6785 $Y=11331 $D=616
M272 352 20 vss vss hvtnfet l=6e-08 w=4e-07 $X=6785 $Y=12191 $D=616
M273 353 21 vss vss hvtnfet l=6e-08 w=4e-07 $X=6785 $Y=38542 $D=616
M274 354 t_mb<0> vss vss hvtnfet l=6e-08 w=4e-07 $X=6785 $Y=39402 $D=616
M275 129 18 vss vss hvtnfet l=6e-08 w=4e-07 $X=6785 $Y=45897 $D=616
M276 143 128 b_blb<0> vss hvtnfet l=6e-08 w=6e-07 $X=6830 $Y=2941 $D=616
M277 143 128 b_blb<0> vss hvtnfet l=6e-08 w=6e-07 $X=6830 $Y=3201 $D=616
M278 148 122 b_bla_n<0> vss hvtnfet l=6e-08 w=6e-07 $X=6830 $Y=3881 $D=616
M279 148 122 b_bla_n<0> vss hvtnfet l=6e-08 w=6e-07 $X=6830 $Y=4141 $D=616
M280 t_bla_n<0> 123 148 vss hvtnfet l=6e-08 w=6e-07 $X=6830 $Y=46932 $D=616
M281 148 123 t_bla_n<0> vss hvtnfet l=6e-08 w=6e-07 $X=6830 $Y=47192 $D=616
M282 t_blb<0> 129 143 vss hvtnfet l=6e-08 w=6e-07 $X=6830 $Y=47872 $D=616
M283 143 129 t_blb<0> vss hvtnfet l=6e-08 w=6e-07 $X=6830 $Y=48132 $D=616
M284 252 75 85 vss hvtnfet l=1.4e-07 w=7.5e-07 $X=6850 $Y=34593 $D=616
M285 124 bwenb vss vss hvtnfet l=1.4e-07 w=2.1e-07 $X=6895 $Y=14555 $D=616
M286 118 133 vss vss hvtnfet l=1.4e-07 w=2.1e-07 $X=6895 $Y=16755 $D=616
M287 159 125 vss vss hvtnfet l=6e-08 w=6e-07 $X=6897 $Y=26159 $D=616
M288 vss vdd 245 vss hvtnfet l=6e-08 w=3e-07 $X=6950 $Y=17670 $D=616
M289 ddqb_n 85 vss vss hvtnfet l=7e-08 w=3.2e-07 $X=6960 $Y=33798 $D=616
M290 256 vdd vss vss hvtnfet l=6e-08 w=3e-07 $X=7007 $Y=31223 $D=616
M291 vss 126 128 vss hvtnfet l=6e-08 w=4e-07 $X=7045 $Y=4836 $D=616
M292 126 b_cb<0> 351 vss hvtnfet l=6e-08 w=4e-07 $X=7045 $Y=11331 $D=616
M293 131 126 352 vss hvtnfet l=6e-08 w=4e-07 $X=7045 $Y=12191 $D=616
M294 132 127 353 vss hvtnfet l=6e-08 w=4e-07 $X=7045 $Y=38542 $D=616
M295 127 t_cb<0> 354 vss hvtnfet l=6e-08 w=4e-07 $X=7045 $Y=39402 $D=616
M296 vss 127 129 vss hvtnfet l=6e-08 w=4e-07 $X=7045 $Y=45897 $D=616
M297 vss 125 159 vss hvtnfet l=6e-08 w=6e-07 $X=7157 $Y=26159 $D=616
M298 b_blb_n<3> 2 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=187 $Y=-170 $D=636
M299 t_blb_n<3> 3 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=187 $Y=50503 $D=636
M300 vdd vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=205 $Y=35893 $D=636
M301 140 5 b_blb<3> vdd hvtpfet l=6e-08 w=3e-07 $X=210 $Y=1094 $D=636
M302 b_blb<3> 5 140 vdd hvtpfet l=6e-08 w=3e-07 $X=210 $Y=1354 $D=636
M303 b_blb_n<3> 5 141 vdd hvtpfet l=6e-08 w=3e-07 $X=210 $Y=1864 $D=636
M304 141 5 b_blb_n<3> vdd hvtpfet l=6e-08 w=3e-07 $X=210 $Y=2124 $D=636
M305 t_blb_n<3> 6 141 vdd hvtpfet l=6e-08 w=3e-07 $X=210 $Y=48949 $D=636
M306 141 6 t_blb_n<3> vdd hvtpfet l=6e-08 w=3e-07 $X=210 $Y=49209 $D=636
M307 140 6 t_blb<3> vdd hvtpfet l=6e-08 w=3e-07 $X=210 $Y=49719 $D=636
M308 t_blb<3> 6 140 vdd hvtpfet l=6e-08 w=3e-07 $X=210 $Y=49979 $D=636
M309 qa 34 vdd vdd hvtpfet l=6e-08 w=9e-07 $X=298 $Y=19812 $D=636
M310 qa 34 vdd vdd hvtpfet l=6e-08 w=9e-07 $X=298 $Y=20072 $D=636
M311 b_blb<3> 2 b_blb_n<3> vdd hvtpfet l=6e-08 w=8e-07 $X=447 $Y=-170 $D=636
M312 t_blb<3> 3 t_blb_n<3> vdd hvtpfet l=6e-08 w=8e-07 $X=447 $Y=50503 $D=636
M313 359 5 11 vdd hvtpfet l=6e-08 w=8e-07 $X=535 $Y=5556 $D=636
M314 5 b_cb<3> vdd vdd hvtpfet l=6e-08 w=4e-07 $X=535 $Y=10611 $D=636
M315 2 5 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=535 $Y=12911 $D=636
M316 3 6 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=535 $Y=37822 $D=636
M317 6 t_cb<3> vdd vdd hvtpfet l=6e-08 w=4e-07 $X=535 $Y=40122 $D=636
M318 360 6 12 vdd hvtpfet l=6e-08 w=8e-07 $X=535 $Y=44777 $D=636
M319 vdd vdd 152 vdd hvtpfet l=6e-08 w=6e-07 $X=573 $Y=29008 $D=636
M320 vdd bwena 26 vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=605 $Y=15085 $D=636
M321 vdd 13 43 vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=605 $Y=16115 $D=636
M322 174 vdd vdd vdd hvtpfet l=6e-08 w=6e-07 $X=630 $Y=18290 $D=636
M323 14 16 vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=650 $Y=35893 $D=636
M324 361 43 vdd vdd hvtpfet l=6e-08 w=4.8e-07 $X=653 $Y=21012 $D=636
M325 361 8 40 vdd hvtpfet l=6e-08 w=4.8e-07 $X=653 $Y=21202 $D=636
M326 23 40 vdd vdd hvtpfet l=6e-08 w=4.8e-07 $X=653 $Y=22762 $D=636
M327 362 44 vdd vdd hvtpfet l=6e-08 w=4.8e-07 $X=653 $Y=23729 $D=636
M328 362 8 41 vdd hvtpfet l=6e-08 w=4.8e-07 $X=653 $Y=23919 $D=636
M329 vdd 23 148 vdd hvtpfet l=6e-08 w=6e-07 $X=683 $Y=27488 $D=636
M330 14 17 166 vdd hvtpfet l=1e-07 w=2e-07 $X=685 $Y=36723 $D=636
M331 vdd 2 b_blb<3> vdd hvtpfet l=6e-08 w=8e-07 $X=707 $Y=-170 $D=636
M332 vdd 3 t_blb<3> vdd hvtpfet l=6e-08 w=8e-07 $X=707 $Y=50503 $D=636
M333 vdd 18 359 vdd hvtpfet l=6e-08 w=8e-07 $X=795 $Y=5556 $D=636
M334 vdd b_mb<0> 5 vdd hvtpfet l=6e-08 w=4e-07 $X=795 $Y=10611 $D=636
M335 vdd 20 2 vdd hvtpfet l=6e-08 w=4e-07 $X=795 $Y=12911 $D=636
M336 vdd 21 3 vdd hvtpfet l=6e-08 w=4e-07 $X=795 $Y=37822 $D=636
M337 vdd t_mb<0> 6 vdd hvtpfet l=6e-08 w=4e-07 $X=795 $Y=40122 $D=636
M338 vdd 18 360 vdd hvtpfet l=6e-08 w=8e-07 $X=795 $Y=44777 $D=636
M339 vdd 40 10 vdd hvtpfet l=6e-08 w=3.2e-07 $X=813 $Y=21942 $D=636
M340 vdd 41 9 vdd hvtpfet l=6e-08 w=3.2e-07 $X=813 $Y=24659 $D=636
M341 vdd vdd 174 vdd hvtpfet l=6e-08 w=6e-07 $X=890 $Y=18290 $D=636
M342 363 10 40 vdd hvtpfet l=6e-08 w=2.1e-07 $X=923 $Y=21477 $D=636
M343 363 38 vdd vdd hvtpfet l=6e-08 w=2.1e-07 $X=923 $Y=21667 $D=636
M344 364 9 41 vdd hvtpfet l=6e-08 w=2.1e-07 $X=923 $Y=24194 $D=636
M345 364 38 vdd vdd hvtpfet l=6e-08 w=2.1e-07 $X=923 $Y=24384 $D=636
M346 39 26 vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=945 $Y=15085 $D=636
M347 13 42 vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=945 $Y=16115 $D=636
M348 166 17 14 vdd hvtpfet l=1e-07 w=2e-07 $X=985 $Y=36723 $D=636
M349 ddqa_n 14 vdd vdd hvtpfet l=7e-08 w=3.2e-07 $X=990 $Y=32628 $D=636
M350 vdd 16 14 vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=990 $Y=35893 $D=636
M351 365 29 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=1055 $Y=5556 $D=636
M352 27 b_ma<0> vdd vdd hvtpfet l=6e-08 w=4e-07 $X=1055 $Y=10611 $D=636
M353 36 31 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=1055 $Y=12911 $D=636
M354 37 32 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=1055 $Y=37822 $D=636
M355 28 t_ma<0> vdd vdd hvtpfet l=6e-08 w=4e-07 $X=1055 $Y=40122 $D=636
M356 366 29 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=1055 $Y=44777 $D=636
M357 367 17 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=1083 $Y=29008 $D=636
M358 b_bla_n<3> 36 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=1143 $Y=-170 $D=636
M359 t_bla_n<3> 37 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=1143 $Y=50503 $D=636
M360 174 vdd vdd vdd hvtpfet l=6e-08 w=6e-07 $X=1150 $Y=18290 $D=636
M361 29 35 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=1193 $Y=27288 $D=636
M362 49 34 367 vdd hvtpfet l=6e-08 w=6e-07 $X=1273 $Y=29008 $D=636
M363 vdd 14 ddqa_n vdd hvtpfet l=7e-08 w=3.2e-07 $X=1280 $Y=32628 $D=636
M364 14 17 166 vdd hvtpfet l=1e-07 w=2e-07 $X=1285 $Y=36723 $D=636
M365 24 27 365 vdd hvtpfet l=6e-08 w=8e-07 $X=1315 $Y=5556 $D=636
M366 vdd b_ca<3> 27 vdd hvtpfet l=6e-08 w=4e-07 $X=1315 $Y=10611 $D=636
M367 vdd 27 36 vdd hvtpfet l=6e-08 w=4e-07 $X=1315 $Y=12911 $D=636
M368 vdd 28 37 vdd hvtpfet l=6e-08 w=4e-07 $X=1315 $Y=37822 $D=636
M369 vdd t_ca<3> 28 vdd hvtpfet l=6e-08 w=4e-07 $X=1315 $Y=40122 $D=636
M370 25 28 366 vdd hvtpfet l=6e-08 w=8e-07 $X=1315 $Y=44777 $D=636
M371 16 14 vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=1330 $Y=35893 $D=636
M372 166 27 b_bla<3> vdd hvtpfet l=6e-08 w=3e-07 $X=1400 $Y=1094 $D=636
M373 b_bla<3> 27 166 vdd hvtpfet l=6e-08 w=3e-07 $X=1400 $Y=1354 $D=636
M374 b_bla_n<3> 27 167 vdd hvtpfet l=6e-08 w=3e-07 $X=1400 $Y=1864 $D=636
M375 167 27 b_bla_n<3> vdd hvtpfet l=6e-08 w=3e-07 $X=1400 $Y=2124 $D=636
M376 t_bla_n<3> 28 167 vdd hvtpfet l=6e-08 w=3e-07 $X=1400 $Y=48949 $D=636
M377 167 28 t_bla_n<3> vdd hvtpfet l=6e-08 w=3e-07 $X=1400 $Y=49209 $D=636
M378 166 28 t_bla<3> vdd hvtpfet l=6e-08 w=3e-07 $X=1400 $Y=49719 $D=636
M379 t_bla<3> 28 166 vdd hvtpfet l=6e-08 w=3e-07 $X=1400 $Y=49979 $D=636
M380 b_bla<3> 36 b_bla_n<3> vdd hvtpfet l=6e-08 w=8e-07 $X=1403 $Y=-170 $D=636
M381 t_bla<3> 37 t_bla_n<3> vdd hvtpfet l=6e-08 w=8e-07 $X=1403 $Y=50503 $D=636
M382 vdd vdd 174 vdd hvtpfet l=6e-08 w=6e-07 $X=1410 $Y=18290 $D=636
M383 vdd 35 29 vdd hvtpfet l=6e-08 w=8e-07 $X=1453 $Y=27288 $D=636
M384 368 14 49 vdd hvtpfet l=6e-08 w=6e-07 $X=1533 $Y=29008 $D=636
M385 vdd 39 52 vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=1535 $Y=15085 $D=636
M386 vdd 47 42 vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=1535 $Y=16115 $D=636
M387 14 sa_prea_n vdd vdd hvtpfet l=1e-07 w=6e-07 $X=1560 $Y=32628 $D=636
M388 166 17 14 vdd hvtpfet l=1e-07 w=2e-07 $X=1585 $Y=36723 $D=636
M389 vdd 36 b_bla<3> vdd hvtpfet l=6e-08 w=8e-07 $X=1663 $Y=-170 $D=636
M390 vdd 37 t_bla<3> vdd hvtpfet l=6e-08 w=8e-07 $X=1663 $Y=50503 $D=636
M391 174 vdd vdd vdd hvtpfet l=6e-08 w=6e-07 $X=1670 $Y=18290 $D=636
M392 vdd 14 16 vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=1670 $Y=35893 $D=636
M393 29 lwea vdd vdd hvtpfet l=6e-08 w=8e-07 $X=1713 $Y=27288 $D=636
M394 vdd saea_n 368 vdd hvtpfet l=6e-08 w=6e-07 $X=1723 $Y=29008 $D=636
M395 16 sa_prea_n 14 vdd hvtpfet l=1e-07 w=6e-07 $X=1860 $Y=32628 $D=636
M396 44 52 vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=1875 $Y=15085 $D=636
M397 47 da vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=1875 $Y=16115 $D=636
M398 vdd vdd 174 vdd hvtpfet l=6e-08 w=6e-07 $X=1930 $Y=18290 $D=636
M399 vdd lwea 29 vdd hvtpfet l=6e-08 w=8e-07 $X=1973 $Y=27288 $D=636
M400 14 16 vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=2010 $Y=35893 $D=636
M401 b_bla<2> 58 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=2097 $Y=-170 $D=636
M402 t_bla<2> 59 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=2097 $Y=50503 $D=636
M403 166 55 b_bla<2> vdd hvtpfet l=6e-08 w=3e-07 $X=2120 $Y=1094 $D=636
M404 b_bla<2> 55 166 vdd hvtpfet l=6e-08 w=3e-07 $X=2120 $Y=1354 $D=636
M405 b_bla_n<2> 55 167 vdd hvtpfet l=6e-08 w=3e-07 $X=2120 $Y=1864 $D=636
M406 167 55 b_bla_n<2> vdd hvtpfet l=6e-08 w=3e-07 $X=2120 $Y=2124 $D=636
M407 t_bla_n<2> 56 167 vdd hvtpfet l=6e-08 w=3e-07 $X=2120 $Y=48949 $D=636
M408 167 56 t_bla_n<2> vdd hvtpfet l=6e-08 w=3e-07 $X=2120 $Y=49209 $D=636
M409 166 56 t_bla<2> vdd hvtpfet l=6e-08 w=3e-07 $X=2120 $Y=49719 $D=636
M410 t_bla<2> 56 166 vdd hvtpfet l=6e-08 w=3e-07 $X=2120 $Y=49979 $D=636
M411 16 17 167 vdd hvtpfet l=1e-07 w=2e-07 $X=2135 $Y=36723 $D=636
M412 vdd sa_prea_n 16 vdd hvtpfet l=1e-07 w=6e-07 $X=2160 $Y=32628 $D=636
M413 vdd 16 14 vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=2350 $Y=35893 $D=636
M414 b_bla_n<2> 58 b_bla<2> vdd hvtpfet l=6e-08 w=8e-07 $X=2357 $Y=-170 $D=636
M415 t_bla_n<2> 59 t_bla<2> vdd hvtpfet l=6e-08 w=8e-07 $X=2357 $Y=50503 $D=636
M416 167 17 16 vdd hvtpfet l=1e-07 w=2e-07 $X=2435 $Y=36723 $D=636
M417 31 b_tm_prea_n vdd vdd hvtpfet l=6e-08 w=5e-07 $X=2440 $Y=18290 $D=636
M418 373 55 61 vdd hvtpfet l=6e-08 w=8e-07 $X=2445 $Y=5556 $D=636
M419 55 b_ca<2> vdd vdd hvtpfet l=6e-08 w=4e-07 $X=2445 $Y=10611 $D=636
M420 58 55 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=2445 $Y=12911 $D=636
M421 59 56 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=2445 $Y=37822 $D=636
M422 56 t_ca<2> vdd vdd hvtpfet l=6e-08 w=4e-07 $X=2445 $Y=40122 $D=636
M423 374 56 62 vdd hvtpfet l=6e-08 w=8e-07 $X=2445 $Y=44777 $D=636
M424 ddqa 16 vdd vdd hvtpfet l=7e-08 w=3.2e-07 $X=2470 $Y=32628 $D=636
M425 169 40 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=2493 $Y=27488 $D=636
M426 vdd 58 b_bla_n<2> vdd hvtpfet l=6e-08 w=8e-07 $X=2617 $Y=-170 $D=636
M427 vdd 59 t_bla_n<2> vdd hvtpfet l=6e-08 w=8e-07 $X=2617 $Y=50503 $D=636
M428 vdd 49 34 vdd hvtpfet l=6e-08 w=6e-07 $X=2633 $Y=29008 $D=636
M429 16 14 vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=2690 $Y=35893 $D=636
M430 vdd b_tm_prea_n 31 vdd hvtpfet l=6e-08 w=5e-07 $X=2700 $Y=18290 $D=636
M431 vdd 29 373 vdd hvtpfet l=6e-08 w=8e-07 $X=2705 $Y=5556 $D=636
M432 vdd b_ma<0> 55 vdd hvtpfet l=6e-08 w=4e-07 $X=2705 $Y=10611 $D=636
M433 vdd 31 58 vdd hvtpfet l=6e-08 w=4e-07 $X=2705 $Y=12911 $D=636
M434 vdd 32 59 vdd hvtpfet l=6e-08 w=4e-07 $X=2705 $Y=37822 $D=636
M435 vdd t_ma<0> 56 vdd hvtpfet l=6e-08 w=4e-07 $X=2705 $Y=40122 $D=636
M436 vdd 29 374 vdd hvtpfet l=6e-08 w=8e-07 $X=2705 $Y=44777 $D=636
M437 16 17 167 vdd hvtpfet l=1e-07 w=2e-07 $X=2735 $Y=36723 $D=636
M438 vdd 16 ddqa vdd hvtpfet l=7e-08 w=3.2e-07 $X=2760 $Y=32628 $D=636
M439 17 saea_n vdd vdd hvtpfet l=6e-08 w=6e-07 $X=2893 $Y=29008 $D=636
M440 32 t_tm_prea_n vdd vdd hvtpfet l=6e-08 w=5e-07 $X=2960 $Y=18290 $D=636
M441 375 18 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=2965 $Y=5556 $D=636
M442 66 b_mb<0> vdd vdd hvtpfet l=6e-08 w=4e-07 $X=2965 $Y=10611 $D=636
M443 70 20 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=2965 $Y=12911 $D=636
M444 71 21 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=2965 $Y=37822 $D=636
M445 67 t_mb<0> vdd vdd hvtpfet l=6e-08 w=4e-07 $X=2965 $Y=40122 $D=636
M446 376 18 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=2965 $Y=44777 $D=636
M447 vdd 14 16 vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=3030 $Y=35893 $D=636
M448 167 17 16 vdd hvtpfet l=1e-07 w=2e-07 $X=3035 $Y=36723 $D=636
M449 b_blb<2> 70 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=3053 $Y=-170 $D=636
M450 t_blb<2> 71 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=3053 $Y=50503 $D=636
M451 38 clk_dqa vdd vdd hvtpfet l=6e-08 w=4e-07 $X=3165 $Y=21427 $D=636
M452 8 clk_dqa_n vdd vdd hvtpfet l=6e-08 w=4e-07 $X=3165 $Y=23694 $D=636
M453 65 41 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=3165 $Y=24394 $D=636
M454 35 65 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=3165 $Y=24904 $D=636
M455 vdd t_tm_prea_n 32 vdd hvtpfet l=6e-08 w=5e-07 $X=3220 $Y=18290 $D=636
M456 68 66 375 vdd hvtpfet l=6e-08 w=8e-07 $X=3225 $Y=5556 $D=636
M457 vdd b_cb<2> 66 vdd hvtpfet l=6e-08 w=4e-07 $X=3225 $Y=10611 $D=636
M458 vdd 66 70 vdd hvtpfet l=6e-08 w=4e-07 $X=3225 $Y=12911 $D=636
M459 vdd 67 71 vdd hvtpfet l=6e-08 w=4e-07 $X=3225 $Y=37822 $D=636
M460 vdd t_cb<2> 67 vdd hvtpfet l=6e-08 w=4e-07 $X=3225 $Y=40122 $D=636
M461 69 67 376 vdd hvtpfet l=6e-08 w=8e-07 $X=3225 $Y=44777 $D=636
M462 140 66 b_blb<2> vdd hvtpfet l=6e-08 w=3e-07 $X=3310 $Y=1094 $D=636
M463 b_blb<2> 66 140 vdd hvtpfet l=6e-08 w=3e-07 $X=3310 $Y=1354 $D=636
M464 b_blb_n<2> 66 141 vdd hvtpfet l=6e-08 w=3e-07 $X=3310 $Y=1864 $D=636
M465 141 66 b_blb_n<2> vdd hvtpfet l=6e-08 w=3e-07 $X=3310 $Y=2124 $D=636
M466 t_blb_n<2> 67 141 vdd hvtpfet l=6e-08 w=3e-07 $X=3310 $Y=48949 $D=636
M467 141 67 t_blb_n<2> vdd hvtpfet l=6e-08 w=3e-07 $X=3310 $Y=49209 $D=636
M468 140 67 t_blb<2> vdd hvtpfet l=6e-08 w=3e-07 $X=3310 $Y=49719 $D=636
M469 t_blb<2> 67 140 vdd hvtpfet l=6e-08 w=3e-07 $X=3310 $Y=49979 $D=636
M470 b_blb_n<2> 70 b_blb<2> vdd hvtpfet l=6e-08 w=8e-07 $X=3313 $Y=-170 $D=636
M471 t_blb_n<2> 71 t_blb<2> vdd hvtpfet l=6e-08 w=8e-07 $X=3313 $Y=50503 $D=636
M472 202 16 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=3403 $Y=29008 $D=636
M473 vdd vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=3475 $Y=35893 $D=636
M474 vdd 70 b_blb_n<2> vdd hvtpfet l=6e-08 w=8e-07 $X=3573 $Y=-170 $D=636
M475 vdd 71 t_blb_n<2> vdd hvtpfet l=6e-08 w=8e-07 $X=3573 $Y=50503 $D=636
M476 b_blb_n<1> 76 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=4007 $Y=-170 $D=636
M477 t_blb_n<1> 77 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=4007 $Y=50503 $D=636
M478 vdd vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=4025 $Y=35893 $D=636
M479 140 79 b_blb<1> vdd hvtpfet l=6e-08 w=3e-07 $X=4030 $Y=1094 $D=636
M480 b_blb<1> 79 140 vdd hvtpfet l=6e-08 w=3e-07 $X=4030 $Y=1354 $D=636
M481 b_blb_n<1> 79 141 vdd hvtpfet l=6e-08 w=3e-07 $X=4030 $Y=1864 $D=636
M482 141 79 b_blb_n<1> vdd hvtpfet l=6e-08 w=3e-07 $X=4030 $Y=2124 $D=636
M483 t_blb_n<1> 80 141 vdd hvtpfet l=6e-08 w=3e-07 $X=4030 $Y=48949 $D=636
M484 141 80 t_blb_n<1> vdd hvtpfet l=6e-08 w=3e-07 $X=4030 $Y=49209 $D=636
M485 140 80 t_blb<1> vdd hvtpfet l=6e-08 w=3e-07 $X=4030 $Y=49719 $D=636
M486 t_blb<1> 80 140 vdd hvtpfet l=6e-08 w=3e-07 $X=4030 $Y=49979 $D=636
M487 107 clk_dqb vdd vdd hvtpfet l=6e-08 w=4e-07 $X=4075 $Y=21427 $D=636
M488 105 clk_dqb_n vdd vdd hvtpfet l=6e-08 w=4e-07 $X=4075 $Y=23694 $D=636
M489 89 88 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=4075 $Y=24394 $D=636
M490 117 89 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=4075 $Y=24904 $D=636
M491 vdd 75 209 vdd hvtpfet l=6e-08 w=6e-07 $X=4177 $Y=29008 $D=636
M492 b_blb<1> 76 b_blb_n<1> vdd hvtpfet l=6e-08 w=8e-07 $X=4267 $Y=-170 $D=636
M493 t_blb<1> 77 t_blb_n<1> vdd hvtpfet l=6e-08 w=8e-07 $X=4267 $Y=50503 $D=636
M494 381 79 83 vdd hvtpfet l=6e-08 w=8e-07 $X=4355 $Y=5556 $D=636
M495 79 b_cb<1> vdd vdd hvtpfet l=6e-08 w=4e-07 $X=4355 $Y=10611 $D=636
M496 76 79 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=4355 $Y=12911 $D=636
M497 77 80 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=4355 $Y=37822 $D=636
M498 80 t_cb<1> vdd vdd hvtpfet l=6e-08 w=4e-07 $X=4355 $Y=40122 $D=636
M499 382 80 84 vdd hvtpfet l=6e-08 w=8e-07 $X=4355 $Y=44777 $D=636
M500 21 t_tm_preb_n vdd vdd hvtpfet l=6e-08 w=5e-07 $X=4360 $Y=18290 $D=636
M501 75 85 vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=4470 $Y=35893 $D=636
M502 75 86 141 vdd hvtpfet l=1e-07 w=2e-07 $X=4505 $Y=36723 $D=636
M503 vdd 76 b_blb<1> vdd hvtpfet l=6e-08 w=8e-07 $X=4527 $Y=-170 $D=636
M504 vdd 77 t_blb<1> vdd hvtpfet l=6e-08 w=8e-07 $X=4527 $Y=50503 $D=636
M505 vdd 18 381 vdd hvtpfet l=6e-08 w=8e-07 $X=4615 $Y=5556 $D=636
M506 vdd b_mb<0> 79 vdd hvtpfet l=6e-08 w=4e-07 $X=4615 $Y=10611 $D=636
M507 vdd 20 76 vdd hvtpfet l=6e-08 w=4e-07 $X=4615 $Y=12911 $D=636
M508 vdd 21 77 vdd hvtpfet l=6e-08 w=4e-07 $X=4615 $Y=37822 $D=636
M509 vdd t_mb<0> 80 vdd hvtpfet l=6e-08 w=4e-07 $X=4615 $Y=40122 $D=636
M510 vdd 18 382 vdd hvtpfet l=6e-08 w=8e-07 $X=4615 $Y=44777 $D=636
M511 vdd t_tm_preb_n 21 vdd hvtpfet l=6e-08 w=5e-07 $X=4620 $Y=18290 $D=636
M512 vdd saeb_n 86 vdd hvtpfet l=6e-08 w=6e-07 $X=4687 $Y=29008 $D=636
M513 141 86 75 vdd hvtpfet l=1e-07 w=2e-07 $X=4805 $Y=36723 $D=636
M514 ddqb 75 vdd vdd hvtpfet l=7e-08 w=3.2e-07 $X=4810 $Y=32628 $D=636
M515 vdd 85 75 vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=4810 $Y=35893 $D=636
M516 383 29 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=4875 $Y=5556 $D=636
M517 94 b_ma<0> vdd vdd hvtpfet l=6e-08 w=4e-07 $X=4875 $Y=10611 $D=636
M518 97 31 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=4875 $Y=12911 $D=636
M519 98 32 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=4875 $Y=37822 $D=636
M520 95 t_ma<0> vdd vdd hvtpfet l=6e-08 w=4e-07 $X=4875 $Y=40122 $D=636
M521 384 29 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=4875 $Y=44777 $D=636
M522 20 b_tm_preb_n vdd vdd hvtpfet l=6e-08 w=5e-07 $X=4880 $Y=18290 $D=636
M523 104 109 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=4947 $Y=29008 $D=636
M524 b_bla_n<1> 97 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=4963 $Y=-170 $D=636
M525 t_bla_n<1> 98 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=4963 $Y=50503 $D=636
M526 vdd 93 143 vdd hvtpfet l=6e-08 w=6e-07 $X=5087 $Y=27488 $D=636
M527 vdd 75 ddqb vdd hvtpfet l=7e-08 w=3.2e-07 $X=5100 $Y=32628 $D=636
M528 75 86 141 vdd hvtpfet l=1e-07 w=2e-07 $X=5105 $Y=36723 $D=636
M529 91 94 383 vdd hvtpfet l=6e-08 w=8e-07 $X=5135 $Y=5556 $D=636
M530 vdd b_ca<1> 94 vdd hvtpfet l=6e-08 w=4e-07 $X=5135 $Y=10611 $D=636
M531 vdd 94 97 vdd hvtpfet l=6e-08 w=4e-07 $X=5135 $Y=12911 $D=636
M532 vdd 95 98 vdd hvtpfet l=6e-08 w=4e-07 $X=5135 $Y=37822 $D=636
M533 vdd t_ca<1> 95 vdd hvtpfet l=6e-08 w=4e-07 $X=5135 $Y=40122 $D=636
M534 92 95 384 vdd hvtpfet l=6e-08 w=8e-07 $X=5135 $Y=44777 $D=636
M535 vdd b_tm_preb_n 20 vdd hvtpfet l=6e-08 w=5e-07 $X=5140 $Y=18290 $D=636
M536 85 75 vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=5150 $Y=35893 $D=636
M537 166 94 b_bla<1> vdd hvtpfet l=6e-08 w=3e-07 $X=5220 $Y=1094 $D=636
M538 b_bla<1> 94 166 vdd hvtpfet l=6e-08 w=3e-07 $X=5220 $Y=1354 $D=636
M539 b_bla_n<1> 94 167 vdd hvtpfet l=6e-08 w=3e-07 $X=5220 $Y=1864 $D=636
M540 167 94 b_bla_n<1> vdd hvtpfet l=6e-08 w=3e-07 $X=5220 $Y=2124 $D=636
M541 t_bla_n<1> 95 167 vdd hvtpfet l=6e-08 w=3e-07 $X=5220 $Y=48949 $D=636
M542 167 95 t_bla_n<1> vdd hvtpfet l=6e-08 w=3e-07 $X=5220 $Y=49209 $D=636
M543 166 95 t_bla<1> vdd hvtpfet l=6e-08 w=3e-07 $X=5220 $Y=49719 $D=636
M544 t_bla<1> 95 166 vdd hvtpfet l=6e-08 w=3e-07 $X=5220 $Y=49979 $D=636
M545 b_bla<1> 97 b_bla_n<1> vdd hvtpfet l=6e-08 w=8e-07 $X=5223 $Y=-170 $D=636
M546 t_bla<1> 98 t_bla_n<1> vdd hvtpfet l=6e-08 w=8e-07 $X=5223 $Y=50503 $D=636
M547 75 sa_preb_n vdd vdd hvtpfet l=1e-07 w=6e-07 $X=5380 $Y=32628 $D=636
M548 141 86 75 vdd hvtpfet l=1e-07 w=2e-07 $X=5405 $Y=36723 $D=636
M549 vdd 97 b_bla<1> vdd hvtpfet l=6e-08 w=8e-07 $X=5483 $Y=-170 $D=636
M550 vdd 98 t_bla<1> vdd hvtpfet l=6e-08 w=8e-07 $X=5483 $Y=50503 $D=636
M551 vdd 75 85 vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=5490 $Y=35893 $D=636
M552 18 lweb vdd vdd hvtpfet l=6e-08 w=8e-07 $X=5607 $Y=27288 $D=636
M553 vdd 106 119 vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=5625 $Y=15085 $D=636
M554 vdd db 110 vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=5625 $Y=16115 $D=636
M555 245 vdd vdd vdd hvtpfet l=6e-08 w=6e-07 $X=5650 $Y=18290 $D=636
M556 85 sa_preb_n 75 vdd hvtpfet l=1e-07 w=6e-07 $X=5680 $Y=32628 $D=636
M557 75 85 vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=5830 $Y=35893 $D=636
M558 385 saeb_n vdd vdd hvtpfet l=6e-08 w=6e-07 $X=5857 $Y=29008 $D=636
M559 vdd lweb 18 vdd hvtpfet l=6e-08 w=8e-07 $X=5867 $Y=27288 $D=636
M560 vdd vdd 245 vdd hvtpfet l=6e-08 w=6e-07 $X=5910 $Y=18290 $D=636
M561 b_bla<0> 115 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=5917 $Y=-170 $D=636
M562 t_bla<0> 116 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=5917 $Y=50503 $D=636
M563 166 112 b_bla<0> vdd hvtpfet l=6e-08 w=3e-07 $X=5940 $Y=1094 $D=636
M564 b_bla<0> 112 166 vdd hvtpfet l=6e-08 w=3e-07 $X=5940 $Y=1354 $D=636
M565 b_bla_n<0> 112 167 vdd hvtpfet l=6e-08 w=3e-07 $X=5940 $Y=1864 $D=636
M566 167 112 b_bla_n<0> vdd hvtpfet l=6e-08 w=3e-07 $X=5940 $Y=2124 $D=636
M567 t_bla_n<0> 113 167 vdd hvtpfet l=6e-08 w=3e-07 $X=5940 $Y=48949 $D=636
M568 167 113 t_bla_n<0> vdd hvtpfet l=6e-08 w=3e-07 $X=5940 $Y=49209 $D=636
M569 166 113 t_bla<0> vdd hvtpfet l=6e-08 w=3e-07 $X=5940 $Y=49719 $D=636
M570 t_bla<0> 113 166 vdd hvtpfet l=6e-08 w=3e-07 $X=5940 $Y=49979 $D=636
M571 85 86 140 vdd hvtpfet l=1e-07 w=2e-07 $X=5955 $Y=36723 $D=636
M572 106 121 vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=5965 $Y=15085 $D=636
M573 120 110 vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=5965 $Y=16115 $D=636
M574 vdd sa_preb_n 85 vdd hvtpfet l=1e-07 w=6e-07 $X=5980 $Y=32628 $D=636
M575 109 85 385 vdd hvtpfet l=6e-08 w=6e-07 $X=6047 $Y=29008 $D=636
M576 18 117 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=6127 $Y=27288 $D=636
M577 245 vdd vdd vdd hvtpfet l=6e-08 w=6e-07 $X=6170 $Y=18290 $D=636
M578 vdd 85 75 vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=6170 $Y=35893 $D=636
M579 b_bla_n<0> 115 b_bla<0> vdd hvtpfet l=6e-08 w=8e-07 $X=6177 $Y=-170 $D=636
M580 t_bla_n<0> 116 t_bla<0> vdd hvtpfet l=6e-08 w=8e-07 $X=6177 $Y=50503 $D=636
M581 140 86 85 vdd hvtpfet l=1e-07 w=2e-07 $X=6255 $Y=36723 $D=636
M582 390 112 122 vdd hvtpfet l=6e-08 w=8e-07 $X=6265 $Y=5556 $D=636
M583 112 b_ca<0> vdd vdd hvtpfet l=6e-08 w=4e-07 $X=6265 $Y=10611 $D=636
M584 115 112 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=6265 $Y=12911 $D=636
M585 116 113 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=6265 $Y=37822 $D=636
M586 113 t_ca<0> vdd vdd hvtpfet l=6e-08 w=4e-07 $X=6265 $Y=40122 $D=636
M587 391 113 123 vdd hvtpfet l=6e-08 w=8e-07 $X=6265 $Y=44777 $D=636
M588 ddqb_n 85 vdd vdd hvtpfet l=7e-08 w=3.2e-07 $X=6290 $Y=32628 $D=636
M589 392 104 109 vdd hvtpfet l=6e-08 w=6e-07 $X=6307 $Y=29008 $D=636
M590 vdd 117 18 vdd hvtpfet l=6e-08 w=8e-07 $X=6387 $Y=27288 $D=636
M591 vdd vdd 245 vdd hvtpfet l=6e-08 w=6e-07 $X=6430 $Y=18290 $D=636
M592 vdd 115 b_bla_n<0> vdd hvtpfet l=6e-08 w=8e-07 $X=6437 $Y=-170 $D=636
M593 vdd 116 t_bla_n<0> vdd hvtpfet l=6e-08 w=8e-07 $X=6437 $Y=50503 $D=636
M594 qb 104 vdd vdd hvtpfet l=6e-08 w=9e-07 $X=6442 $Y=19812 $D=636
M595 qb 104 vdd vdd hvtpfet l=6e-08 w=9e-07 $X=6442 $Y=20072 $D=636
M596 vdd 86 392 vdd hvtpfet l=6e-08 w=6e-07 $X=6497 $Y=29008 $D=636
M597 393 118 vdd vdd hvtpfet l=6e-08 w=4.8e-07 $X=6507 $Y=21012 $D=636
M598 393 105 93 vdd hvtpfet l=6e-08 w=4.8e-07 $X=6507 $Y=21202 $D=636
M599 394 134 93 vdd hvtpfet l=6e-08 w=2.1e-07 $X=6507 $Y=21477 $D=636
M600 394 107 vdd vdd hvtpfet l=6e-08 w=2.1e-07 $X=6507 $Y=21667 $D=636
M601 vdd 93 134 vdd hvtpfet l=6e-08 w=3.2e-07 $X=6507 $Y=21942 $D=636
M602 125 93 vdd vdd hvtpfet l=6e-08 w=4.8e-07 $X=6507 $Y=22762 $D=636
M603 395 119 vdd vdd hvtpfet l=6e-08 w=4.8e-07 $X=6507 $Y=23729 $D=636
M604 395 105 88 vdd hvtpfet l=6e-08 w=4.8e-07 $X=6507 $Y=23919 $D=636
M605 396 137 88 vdd hvtpfet l=6e-08 w=2.1e-07 $X=6507 $Y=24194 $D=636
M606 396 107 vdd vdd hvtpfet l=6e-08 w=2.1e-07 $X=6507 $Y=24384 $D=636
M607 vdd 88 137 vdd hvtpfet l=6e-08 w=3.2e-07 $X=6507 $Y=24659 $D=636
M608 85 75 vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=6510 $Y=35893 $D=636
M609 vdd 29 390 vdd hvtpfet l=6e-08 w=8e-07 $X=6525 $Y=5556 $D=636
M610 vdd b_ma<0> 112 vdd hvtpfet l=6e-08 w=4e-07 $X=6525 $Y=10611 $D=636
M611 vdd 31 115 vdd hvtpfet l=6e-08 w=4e-07 $X=6525 $Y=12911 $D=636
M612 vdd 32 116 vdd hvtpfet l=6e-08 w=4e-07 $X=6525 $Y=37822 $D=636
M613 vdd t_ma<0> 113 vdd hvtpfet l=6e-08 w=4e-07 $X=6525 $Y=40122 $D=636
M614 vdd 29 391 vdd hvtpfet l=6e-08 w=8e-07 $X=6525 $Y=44777 $D=636
M615 vdd 124 121 vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=6555 $Y=15085 $D=636
M616 vdd 120 133 vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=6555 $Y=16115 $D=636
M617 85 86 140 vdd hvtpfet l=1e-07 w=2e-07 $X=6555 $Y=36723 $D=636
M618 vdd 85 ddqb_n vdd hvtpfet l=7e-08 w=3.2e-07 $X=6580 $Y=32628 $D=636
M619 245 vdd vdd vdd hvtpfet l=6e-08 w=6e-07 $X=6690 $Y=18290 $D=636
M620 397 18 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=6785 $Y=5556 $D=636
M621 126 b_mb<0> vdd vdd hvtpfet l=6e-08 w=4e-07 $X=6785 $Y=10611 $D=636
M622 131 20 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=6785 $Y=12911 $D=636
M623 132 21 vdd vdd hvtpfet l=6e-08 w=4e-07 $X=6785 $Y=37822 $D=636
M624 127 t_mb<0> vdd vdd hvtpfet l=6e-08 w=4e-07 $X=6785 $Y=40122 $D=636
M625 398 18 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=6785 $Y=44777 $D=636
M626 vdd 75 85 vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=6850 $Y=35893 $D=636
M627 140 86 85 vdd hvtpfet l=1e-07 w=2e-07 $X=6855 $Y=36723 $D=636
M628 b_blb<0> 131 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=6873 $Y=-170 $D=636
M629 t_blb<0> 132 vdd vdd hvtpfet l=6e-08 w=8e-07 $X=6873 $Y=50503 $D=636
M630 124 bwenb vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=6895 $Y=15085 $D=636
M631 118 133 vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=6895 $Y=16115 $D=636
M632 159 125 vdd vdd hvtpfet l=6e-08 w=6e-07 $X=6897 $Y=27488 $D=636
M633 vdd vdd 245 vdd hvtpfet l=6e-08 w=6e-07 $X=6950 $Y=18290 $D=636
M634 256 vdd vdd vdd hvtpfet l=6e-08 w=6e-07 $X=7007 $Y=29008 $D=636
M635 128 126 397 vdd hvtpfet l=6e-08 w=8e-07 $X=7045 $Y=5556 $D=636
M636 vdd b_cb<0> 126 vdd hvtpfet l=6e-08 w=4e-07 $X=7045 $Y=10611 $D=636
M637 vdd 126 131 vdd hvtpfet l=6e-08 w=4e-07 $X=7045 $Y=12911 $D=636
M638 vdd 127 132 vdd hvtpfet l=6e-08 w=4e-07 $X=7045 $Y=37822 $D=636
M639 vdd t_cb<0> 127 vdd hvtpfet l=6e-08 w=4e-07 $X=7045 $Y=40122 $D=636
M640 129 127 398 vdd hvtpfet l=6e-08 w=8e-07 $X=7045 $Y=44777 $D=636
M641 140 126 b_blb<0> vdd hvtpfet l=6e-08 w=3e-07 $X=7130 $Y=1094 $D=636
M642 b_blb<0> 126 140 vdd hvtpfet l=6e-08 w=3e-07 $X=7130 $Y=1354 $D=636
M643 b_blb_n<0> 126 141 vdd hvtpfet l=6e-08 w=3e-07 $X=7130 $Y=1864 $D=636
M644 141 126 b_blb_n<0> vdd hvtpfet l=6e-08 w=3e-07 $X=7130 $Y=2124 $D=636
M645 t_blb_n<0> 127 141 vdd hvtpfet l=6e-08 w=3e-07 $X=7130 $Y=48949 $D=636
M646 141 127 t_blb_n<0> vdd hvtpfet l=6e-08 w=3e-07 $X=7130 $Y=49209 $D=636
M647 140 127 t_blb<0> vdd hvtpfet l=6e-08 w=3e-07 $X=7130 $Y=49719 $D=636
M648 t_blb<0> 127 140 vdd hvtpfet l=6e-08 w=3e-07 $X=7130 $Y=49979 $D=636
M649 b_blb_n<0> 131 b_blb<0> vdd hvtpfet l=6e-08 w=8e-07 $X=7133 $Y=-170 $D=636
M650 t_blb_n<0> 132 t_blb<0> vdd hvtpfet l=6e-08 w=8e-07 $X=7133 $Y=50503 $D=636
M651 vdd vdd vdd vdd hvtpfet l=1.4e-07 w=3.2e-07 $X=7295 $Y=35893 $D=636
M652 vdd 131 b_blb_n<0> vdd hvtpfet l=6e-08 w=8e-07 $X=7393 $Y=-170 $D=636
M653 vdd 132 t_blb_n<0> vdd hvtpfet l=6e-08 w=8e-07 $X=7393 $Y=50503 $D=636
.ends

************************************************************************
* Library Name: XMC55_DPS
* Cell Name:    xmc55_dps_localc4io_dummy
************************************************************************
.SUBCKT xmc55_dps_localc4io_dummy b_dbl b_dwl b_tie_low dbl_pd_n<3> 
+ dbl_pd_n<2> dbl_pd_n<1> dbl_pd_n<0> stclk t_dbl t_dwl t_tie_low vdd vss
** N=889 EP=13 IP=0 FDC=76
M0 vss 2 17 vss hvtnfet l=6e-08 w=2e-07 $X=265 $Y=2781 $D=616
M1 vss 3 18 vss hvtnfet l=6e-08 w=2e-07 $X=265 $Y=48152 $D=616
M2 28 t_dbl vss vss hvtnfet l=6e-08 w=4e-07 $X=340 $Y=26568 $D=616
M3 vss 8 stclk vss hvtnfet l=6e-08 w=3e-07 $X=340 $Y=29928 $D=616
M4 49 b_dwl vss vss hvtnfet l=6e-08 w=4e-07 $X=535 $Y=2781 $D=616
M5 50 t_dwl vss vss hvtnfet l=6e-08 w=4e-07 $X=535 $Y=47952 $D=616
M6 b_tie_low 15 vss vss hvtnfet l=7e-08 w=3.2e-07 $X=540 $Y=4916 $D=616
M7 t_tie_low 16 vss vss hvtnfet l=7e-08 w=3.2e-07 $X=540 $Y=45897 $D=616
M8 8 b_dbl 28 vss hvtnfet l=6e-08 w=4e-07 $X=600 $Y=26568 $D=616
M9 vss dbl_pd_n<2> 12 vss hvtnfet l=6e-08 w=3e-07 $X=630 $Y=19039 $D=616
M10 vss dbl_pd_n<1> 14 vss hvtnfet l=6e-08 w=3e-07 $X=630 $Y=21399 $D=616
M11 vss dbl_pd_n<0> 13 vss hvtnfet l=6e-08 w=3e-07 $X=630 $Y=22329 $D=616
M12 vss dbl_pd_n<3> 21 vss hvtnfet l=6e-08 w=3e-07 $X=630 $Y=24794 $D=616
M13 2 21 49 vss hvtnfet l=6e-08 w=4e-07 $X=795 $Y=2781 $D=616
M14 3 21 50 vss hvtnfet l=6e-08 w=4e-07 $X=795 $Y=47952 $D=616
M15 vdd vdd vdd vdd hvtpfet l=6e-08 w=8e-07 $X=187 $Y=-170 $D=636
M16 vdd vdd vdd vdd hvtpfet l=6e-08 w=8e-07 $X=187 $Y=50503 $D=636
M17 vdd 2 17 vdd hvtpfet l=6e-08 w=4e-07 $X=265 $Y=2061 $D=636
M18 vdd 3 18 vdd hvtpfet l=6e-08 w=4e-07 $X=265 $Y=48672 $D=636
M19 8 t_dbl vdd vdd hvtpfet l=6e-08 w=4e-07 $X=340 $Y=27288 $D=636
M20 vdd 8 stclk vdd hvtpfet l=6e-08 w=6e-07 $X=340 $Y=29008 $D=636
M21 b_dbl vdd vdd vdd hvtpfet l=6e-08 w=8e-07 $X=447 $Y=-170 $D=636
M22 t_dbl vdd vdd vdd hvtpfet l=6e-08 w=8e-07 $X=447 $Y=50503 $D=636
M23 2 b_dwl vdd vdd hvtpfet l=6e-08 w=4e-07 $X=535 $Y=2061 $D=636
M24 3 t_dwl vdd vdd hvtpfet l=6e-08 w=4e-07 $X=535 $Y=48672 $D=636
M25 15 15 vdd vdd hvtpfet l=7e-08 w=6.4e-07 $X=540 $Y=5556 $D=636
M26 16 16 vdd vdd hvtpfet l=7e-08 w=6.4e-07 $X=540 $Y=44937 $D=636
M27 vdd b_dbl 8 vdd hvtpfet l=6e-08 w=4e-07 $X=600 $Y=27288 $D=636
M28 vdd dbl_pd_n<2> 12 vdd hvtpfet l=6e-08 w=5e-07 $X=630 $Y=19659 $D=636
M29 vdd dbl_pd_n<1> 14 vdd hvtpfet l=6e-08 w=5e-07 $X=630 $Y=20579 $D=636
M30 vdd dbl_pd_n<0> 13 vdd hvtpfet l=6e-08 w=5e-07 $X=630 $Y=22949 $D=636
M31 vdd dbl_pd_n<3> 21 vdd hvtpfet l=6e-08 w=5e-07 $X=630 $Y=23974 $D=636
M32 vdd b_dwl b_dbl vdd hvtpfet l=6e-08 w=8e-07 $X=707 $Y=-170 $D=636
M33 vdd t_dwl t_dbl vdd hvtpfet l=6e-08 w=8e-07 $X=707 $Y=50503 $D=636
M34 vdd 21 2 vdd hvtpfet l=6e-08 w=4e-07 $X=795 $Y=2061 $D=636
M35 vdd 21 3 vdd hvtpfet l=6e-08 w=4e-07 $X=795 $Y=48672 $D=636
M36 vss t_tie_low 29 vss srpddnfet l=6e-08 w=3.15e-07 $X=670 $Y=7281 $D=778
M37 vss t_tie_low 30 vss srpddnfet l=6e-08 w=3.15e-07 $X=670 $Y=7876 $D=778
M38 vss t_tie_low 31 vss srpddnfet l=6e-08 w=3.15e-07 $X=670 $Y=9246 $D=778
M39 vss 12 32 vss srpddnfet l=6e-08 w=3.15e-07 $X=670 $Y=10871 $D=778
M40 vss 12 33 vss srpddnfet l=6e-08 w=3.15e-07 $X=670 $Y=11466 $D=778
M41 vss 12 34 vss srpddnfet l=6e-08 w=3.15e-07 $X=670 $Y=13091 $D=778
M42 vss 12 35 vss srpddnfet l=6e-08 w=3.15e-07 $X=670 $Y=13686 $D=778
M43 vss 13 36 vss srpddnfet l=6e-08 w=3.15e-07 $X=670 $Y=15311 $D=778
M44 vss 14 37 vss srpddnfet l=6e-08 w=3.15e-07 $X=670 $Y=16681 $D=778
M45 vss 14 38 vss srpddnfet l=6e-08 w=3.15e-07 $X=670 $Y=17276 $D=778
M46 vss 14 39 vss srpddnfet l=6e-08 w=3.15e-07 $X=670 $Y=33542 $D=778
M47 vss 14 40 vss srpddnfet l=6e-08 w=3.15e-07 $X=670 $Y=34137 $D=778
M48 vss 13 41 vss srpddnfet l=6e-08 w=3.15e-07 $X=670 $Y=35507 $D=778
M49 vss 12 42 vss srpddnfet l=6e-08 w=3.15e-07 $X=670 $Y=37132 $D=778
M50 vss 12 43 vss srpddnfet l=6e-08 w=3.15e-07 $X=670 $Y=37727 $D=778
M51 vss 12 44 vss srpddnfet l=6e-08 w=3.15e-07 $X=670 $Y=39352 $D=778
M52 vss 12 45 vss srpddnfet l=6e-08 w=3.15e-07 $X=670 $Y=39947 $D=778
M53 vss t_tie_low 46 vss srpddnfet l=6e-08 w=3.15e-07 $X=670 $Y=41572 $D=778
M54 vss t_tie_low 47 vss srpddnfet l=6e-08 w=3.15e-07 $X=670 $Y=42942 $D=778
M55 vss t_tie_low 48 vss srpddnfet l=6e-08 w=3.15e-07 $X=670 $Y=43537 $D=778
M56 b_dbl 17 29 vss srpgdnfet l=7.5e-08 w=1.05e-07 $X=655 $Y=6816 $D=780
M57 b_dbl 17 30 vss srpgdnfet l=7.5e-08 w=1.05e-07 $X=655 $Y=8551 $D=780
M58 b_dbl 17 31 vss srpgdnfet l=7.5e-08 w=1.05e-07 $X=655 $Y=9921 $D=780
M59 b_dbl 17 32 vss srpgdnfet l=7.5e-08 w=1.05e-07 $X=655 $Y=10406 $D=780
M60 b_dbl 17 33 vss srpgdnfet l=7.5e-08 w=1.05e-07 $X=655 $Y=12141 $D=780
M61 b_dbl 17 34 vss srpgdnfet l=7.5e-08 w=1.05e-07 $X=655 $Y=12626 $D=780
M62 b_dbl 17 35 vss srpgdnfet l=7.5e-08 w=1.05e-07 $X=655 $Y=14361 $D=780
M63 b_dbl 17 36 vss srpgdnfet l=7.5e-08 w=1.05e-07 $X=655 $Y=14846 $D=780
M64 b_dbl 17 37 vss srpgdnfet l=7.5e-08 w=1.05e-07 $X=655 $Y=16216 $D=780
M65 b_dbl 17 38 vss srpgdnfet l=7.5e-08 w=1.05e-07 $X=655 $Y=17951 $D=780
M66 t_dbl 18 39 vss srpgdnfet l=7.5e-08 w=1.05e-07 $X=655 $Y=33077 $D=780
M67 t_dbl 18 40 vss srpgdnfet l=7.5e-08 w=1.05e-07 $X=655 $Y=34812 $D=780
M68 t_dbl 18 41 vss srpgdnfet l=7.5e-08 w=1.05e-07 $X=655 $Y=36182 $D=780
M69 t_dbl 18 42 vss srpgdnfet l=7.5e-08 w=1.05e-07 $X=655 $Y=36667 $D=780
M70 t_dbl 18 43 vss srpgdnfet l=7.5e-08 w=1.05e-07 $X=655 $Y=38402 $D=780
M71 t_dbl 18 44 vss srpgdnfet l=7.5e-08 w=1.05e-07 $X=655 $Y=38887 $D=780
M72 t_dbl 18 45 vss srpgdnfet l=7.5e-08 w=1.05e-07 $X=655 $Y=40622 $D=780
M73 t_dbl 18 46 vss srpgdnfet l=7.5e-08 w=1.05e-07 $X=655 $Y=41107 $D=780
M74 t_dbl 18 47 vss srpgdnfet l=7.5e-08 w=1.05e-07 $X=655 $Y=42477 $D=780
M75 t_dbl 18 48 vss srpgdnfet l=7.5e-08 w=1.05e-07 $X=655 $Y=44212 $D=780
.ends

************************************************************************
* Library Name: XMC55_DPS
* Cell Name:    xmc55_dps_localc4io_edge
************************************************************************
.SUBCKT xmc55_dps_localc4io_edge tie_low vdd vss
** N=1093 EP=3 IP=0 FDC=59
M0 vss vss vss vss hvtnfet l=6e-08 w=4e-07 $X=970 $Y=2941 $D=616
M1 vss vss vss vss hvtnfet l=6e-08 w=4e-07 $X=970 $Y=3201 $D=616
M2 vss vss vss vss hvtnfet l=6e-08 w=4e-07 $X=970 $Y=3881 $D=616
M3 vss vss vss vss hvtnfet l=6e-08 w=4e-07 $X=970 $Y=4141 $D=616
M4 vss vss vss vss hvtnfet l=6e-08 w=4e-07 $X=970 $Y=46932 $D=616
M5 vss vss vss vss hvtnfet l=6e-08 w=4e-07 $X=970 $Y=47192 $D=616
M6 vss vss vss vss hvtnfet l=6e-08 w=4e-07 $X=970 $Y=47872 $D=616
M7 vss vss vss vss hvtnfet l=6e-08 w=4e-07 $X=970 $Y=48132 $D=616
M8 18 tie_low vss vss hvtnfet l=6e-08 w=2.1e-07 $X=1025 $Y=14555 $D=616
M9 19 tie_low vss vss hvtnfet l=6e-08 w=2.1e-07 $X=1025 $Y=16755 $D=616
M10 20 tie_low vss vss hvtnfet l=6e-08 w=2.1e-07 $X=1025 $Y=17760 $D=616
M11 5 5 vss vss hvtnfet l=6e-08 w=3.2e-07 $X=1025 $Y=26624 $D=616
M12 vss 2 tie_low vss hvtnfet l=6e-08 w=2.1e-07 $X=1025 $Y=33548 $D=616
M13 vss tie_low 10 vss hvtnfet l=6e-08 w=4e-07 $X=1130 $Y=4836 $D=616
M14 vss tie_low 11 vss hvtnfet l=6e-08 w=4e-07 $X=1130 $Y=11331 $D=616
M15 vss tie_low 12 vss hvtnfet l=6e-08 w=4e-07 $X=1130 $Y=12191 $D=616
M16 vss tie_low 13 vss hvtnfet l=6e-08 w=4e-07 $X=1130 $Y=38542 $D=616
M17 vss tie_low 14 vss hvtnfet l=6e-08 w=4e-07 $X=1130 $Y=39402 $D=616
M18 vss tie_low 15 vss hvtnfet l=6e-08 w=4e-07 $X=1130 $Y=45897 $D=616
M19 vss 5 5 vss hvtnfet l=6e-08 w=3.2e-07 $X=1285 $Y=26624 $D=616
M20 vdd vdd vdd vdd hvtpfet l=6e-08 w=3e-07 $X=975 $Y=19812 $D=636
M21 vdd vdd vdd vdd hvtpfet l=6e-08 w=3e-07 $X=975 $Y=20072 $D=636
M22 vdd vdd vdd vdd hvtpfet l=6e-08 w=3e-07 $X=975 $Y=20902 $D=636
M23 vdd vdd vdd vdd hvtpfet l=6e-08 w=3e-07 $X=975 $Y=21162 $D=636
M24 vdd vdd vdd vdd hvtpfet l=6e-08 w=3e-07 $X=975 $Y=21422 $D=636
M25 vdd vdd vdd vdd hvtpfet l=6e-08 w=3e-07 $X=975 $Y=21682 $D=636
M26 vdd vdd vdd vdd hvtpfet l=6e-08 w=3e-07 $X=975 $Y=21942 $D=636
M27 vdd vdd vdd vdd hvtpfet l=6e-08 w=3e-07 $X=975 $Y=22762 $D=636
M28 vdd vdd vdd vdd hvtpfet l=6e-08 w=3e-07 $X=975 $Y=23729 $D=636
M29 vdd vdd vdd vdd hvtpfet l=6e-08 w=3e-07 $X=975 $Y=23989 $D=636
M30 vdd vdd vdd vdd hvtpfet l=6e-08 w=3e-07 $X=975 $Y=24249 $D=636
M31 vdd vdd vdd vdd hvtpfet l=6e-08 w=3e-07 $X=975 $Y=24509 $D=636
M32 vdd vdd vdd vdd hvtpfet l=6e-08 w=3e-07 $X=975 $Y=24769 $D=636
M33 18 tie_low vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=1025 $Y=15085 $D=636
M34 19 tie_low vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=1025 $Y=16115 $D=636
M35 20 tie_low vdd vdd hvtpfet l=6e-08 w=3.2e-07 $X=1025 $Y=18290 $D=636
M36 21 5 2 vdd hvtpfet l=6e-08 w=4.8e-07 $X=1025 $Y=27313 $D=636
M37 22 5 2 vdd hvtpfet l=6e-08 w=4.8e-07 $X=1025 $Y=29008 $D=636
M38 vdd 2 tie_low vdd hvtpfet l=6e-08 w=3.2e-07 $X=1025 $Y=32908 $D=636
M39 vdd vdd vdd vdd hvtpfet l=6e-08 w=3e-07 $X=1070 $Y=1094 $D=636
M40 vdd vdd vdd vdd hvtpfet l=6e-08 w=3e-07 $X=1070 $Y=1354 $D=636
M41 vdd vdd vdd vdd hvtpfet l=6e-08 w=3e-07 $X=1070 $Y=1864 $D=636
M42 vdd vdd vdd vdd hvtpfet l=6e-08 w=3e-07 $X=1070 $Y=2124 $D=636
M43 vdd vdd vdd vdd hvtpfet l=6e-08 w=3e-07 $X=1070 $Y=48949 $D=636
M44 vdd vdd vdd vdd hvtpfet l=6e-08 w=3e-07 $X=1070 $Y=49209 $D=636
M45 vdd vdd vdd vdd hvtpfet l=6e-08 w=3e-07 $X=1070 $Y=49719 $D=636
M46 vdd vdd vdd vdd hvtpfet l=6e-08 w=3e-07 $X=1070 $Y=49979 $D=636
M47 vdd vdd vdd vdd hvtpfet l=6e-08 w=8e-07 $X=1073 $Y=-170 $D=636
M48 vdd vdd vdd vdd hvtpfet l=6e-08 w=8e-07 $X=1073 $Y=50503 $D=636
M49 vdd tie_low 10 vdd hvtpfet l=6e-08 w=8e-07 $X=1130 $Y=5556 $D=636
M50 vdd tie_low 11 vdd hvtpfet l=6e-08 w=4e-07 $X=1130 $Y=10611 $D=636
M51 vdd tie_low 12 vdd hvtpfet l=6e-08 w=4e-07 $X=1130 $Y=12911 $D=636
M52 vdd tie_low 13 vdd hvtpfet l=6e-08 w=4e-07 $X=1130 $Y=37822 $D=636
M53 vdd tie_low 14 vdd hvtpfet l=6e-08 w=4e-07 $X=1130 $Y=40122 $D=636
M54 vdd tie_low 15 vdd hvtpfet l=6e-08 w=8e-07 $X=1130 $Y=44777 $D=636
M55 vdd 5 21 vdd hvtpfet l=6e-08 w=4.8e-07 $X=1285 $Y=27313 $D=636
M56 vdd 5 22 vdd hvtpfet l=6e-08 w=4.8e-07 $X=1285 $Y=29008 $D=636
M57 vdd vdd vdd vdd hvtpfet l=6e-08 w=8e-07 $X=1333 $Y=-170 $D=636
M58 vdd vdd vdd vdd hvtpfet l=6e-08 w=8e-07 $X=1333 $Y=50503 $D=636
.ends

************************************************************************
* Library Name: XMC55_DPS
* Cell Name:    xmc55_dps_collar_dq_4_bw
************************************************************************
.SUBCKT xmc55_dps_collar_dq_4_bw bwena bwena_int bwenb bwenb_int da da_int db 
+ db_int qa qa_int qb qb_int vdd vss
** N=376 EP=14 IP=0 FDC=40
D0 vss bwena diodenx AREA=7.04e-14 $X=367 $Y=130 $D=2
D1 vss da diodenx AREA=7.04e-14 $X=2272 $Y=130 $D=2
D2 vss db diodenx AREA=7.04e-14 $X=4190 $Y=130 $D=2
D3 vss bwenb diodenx AREA=7.04e-14 $X=6095 $Y=130 $D=2
M4 2 bwena vss vss hvtnfet l=6e-08 w=6e-07 $X=580 $Y=1420 $D=616
M5 bwena_int 2 vss vss hvtnfet l=6e-08 w=9e-07 $X=1090 $Y=1120 $D=616
M6 vss 2 bwena_int vss hvtnfet l=6e-08 w=9e-07 $X=1350 $Y=1120 $D=616
M7 qa qa_int vss vss hvtnfet l=6e-08 w=9e-07 $X=1610 $Y=1120 $D=616
M8 vss qa_int qa vss hvtnfet l=6e-08 w=9e-07 $X=1870 $Y=1120 $D=616
M9 vss vdd 14 vss hvtnfet l=6e-08 w=6e-07 $X=2380 $Y=1420 $D=616
M10 6 da vss vss hvtnfet l=6e-08 w=6e-07 $X=2890 $Y=1420 $D=616
M11 da_int 6 vss vss hvtnfet l=6e-08 w=9e-07 $X=3400 $Y=1120 $D=616
M12 vss 6 da_int vss hvtnfet l=6e-08 w=9e-07 $X=3660 $Y=1120 $D=616
M13 db_int 7 vss vss hvtnfet l=6e-08 w=9e-07 $X=3920 $Y=1120 $D=616
M14 vss 7 db_int vss hvtnfet l=6e-08 w=9e-07 $X=4180 $Y=1120 $D=616
M15 vss db 7 vss hvtnfet l=6e-08 w=6e-07 $X=4690 $Y=1420 $D=616
M16 18 vdd vss vss hvtnfet l=6e-08 w=6e-07 $X=5200 $Y=1420 $D=616
M17 qb qb_int vss vss hvtnfet l=6e-08 w=9e-07 $X=5710 $Y=1120 $D=616
M18 vss qb_int qb vss hvtnfet l=6e-08 w=9e-07 $X=5970 $Y=1120 $D=616
M19 bwenb_int 10 vss vss hvtnfet l=6e-08 w=9e-07 $X=6230 $Y=1120 $D=616
M20 vss 10 bwenb_int vss hvtnfet l=6e-08 w=9e-07 $X=6490 $Y=1120 $D=616
M21 vss bwenb 10 vss hvtnfet l=6e-08 w=6e-07 $X=7000 $Y=1420 $D=616
M22 2 bwena vdd vdd hvtpfet l=6e-08 w=1.2e-06 $X=580 $Y=2685 $D=636
M23 bwena_int 2 vdd vdd hvtpfet l=6e-08 w=1.8e-06 $X=1090 $Y=2340 $D=636
M24 vdd 2 bwena_int vdd hvtpfet l=6e-08 w=1.8e-06 $X=1350 $Y=2340 $D=636
M25 qa qa_int vdd vdd hvtpfet l=6e-08 w=1.8e-06 $X=1610 $Y=2340 $D=636
M26 vdd qa_int qa vdd hvtpfet l=6e-08 w=1.8e-06 $X=1870 $Y=2340 $D=636
M27 vdd vdd 14 vdd hvtpfet l=6e-08 w=1.2e-06 $X=2380 $Y=2685 $D=636
M28 6 da vdd vdd hvtpfet l=6e-08 w=1.2e-06 $X=2890 $Y=2685 $D=636
M29 da_int 6 vdd vdd hvtpfet l=6e-08 w=1.8e-06 $X=3400 $Y=2340 $D=636
M30 vdd 6 da_int vdd hvtpfet l=6e-08 w=1.8e-06 $X=3660 $Y=2340 $D=636
M31 db_int 7 vdd vdd hvtpfet l=6e-08 w=1.8e-06 $X=3920 $Y=2340 $D=636
M32 vdd 7 db_int vdd hvtpfet l=6e-08 w=1.8e-06 $X=4180 $Y=2340 $D=636
M33 vdd db 7 vdd hvtpfet l=6e-08 w=1.2e-06 $X=4690 $Y=2685 $D=636
M34 18 vdd vdd vdd hvtpfet l=6e-08 w=1.2e-06 $X=5200 $Y=2685 $D=636
M35 qb qb_int vdd vdd hvtpfet l=6e-08 w=1.8e-06 $X=5710 $Y=2340 $D=636
M36 vdd qb_int qb vdd hvtpfet l=6e-08 w=1.8e-06 $X=5970 $Y=2340 $D=636
M37 bwenb_int 10 vdd vdd hvtpfet l=6e-08 w=1.8e-06 $X=6230 $Y=2340 $D=636
M38 vdd 10 bwenb_int vdd hvtpfet l=6e-08 w=1.8e-06 $X=6490 $Y=2340 $D=636
M39 vdd bwenb 10 vdd hvtpfet l=6e-08 w=1.2e-06 $X=7000 $Y=2685 $D=636
.ends

************************************************************************
* Library Name: XMC55_DPS
* Cell Name:    xmc55_dps_xdec4
************************************************************************
.SUBCKT xmc55_dps_xdec4 pxaa<3> pxaa<2> pxaa<1> pxaa<0> pxab<3> pxab<2> 
+ pxab<1> pxab<0> pxba_n pxbb_n pxca_n pxcb_n vdd vss wla<3> wla<2> wla<1> 
+ wla<0> wlb<3> wlb<2> wlb<1> wlb<0>
** N=963 EP=22 IP=0 FDC=80
M0 wlb<3> 1 vss vss hvtnfet l=6e-08 w=2e-06 $X=5555 $Y=100 $D=616
M1 vss 1 wlb<3> vss hvtnfet l=6e-08 w=2e-06 $X=5555 $Y=365 $D=616
M2 wlb<1> 2 vss vss hvtnfet l=6e-08 w=2e-06 $X=5555 $Y=615 $D=616
M3 vss 2 wlb<1> vss hvtnfet l=6e-08 w=2e-06 $X=5555 $Y=865 $D=616
M4 wlb<0> 3 vss vss hvtnfet l=6e-08 w=2e-06 $X=5555 $Y=1115 $D=616
M5 vss 3 wlb<0> vss hvtnfet l=6e-08 w=2e-06 $X=5555 $Y=1365 $D=616
M6 wlb<2> 4 vss vss hvtnfet l=6e-08 w=2e-06 $X=5555 $Y=1615 $D=616
M7 vss 4 wlb<2> vss hvtnfet l=6e-08 w=2e-06 $X=5555 $Y=1880 $D=616
M8 41 pxab<1> 2 vss hvtnfet l=6e-08 w=2e-06 $X=9205 $Y=615 $D=616
M9 vss 9 41 vss hvtnfet l=6e-08 w=2e-06 $X=9205 $Y=865 $D=616
M10 42 9 vss vss hvtnfet l=6e-08 w=2e-06 $X=9205 $Y=1115 $D=616
M11 42 pxab<0> 3 vss hvtnfet l=6e-08 w=2e-06 $X=9205 $Y=1365 $D=616
M12 43 9 vss vss hvtnfet l=6e-08 w=2e-06 $X=14845 $Y=100 $D=616
M13 1 pxab<3> 43 vss hvtnfet l=6e-08 w=2e-06 $X=14845 $Y=365 $D=616
M14 44 pxab<2> 4 vss hvtnfet l=6e-08 w=2e-06 $X=14845 $Y=1615 $D=616
M15 vss 9 44 vss hvtnfet l=6e-08 w=2e-06 $X=14845 $Y=1880 $D=616
M16 vss pxcb_n 9 vss hvtnfet l=6e-08 w=1e-06 $X=18165 $Y=615 $D=616
M17 9 pxbb_n vss vss hvtnfet l=6e-08 w=1e-06 $X=18165 $Y=865 $D=616
M18 vss pxbb_n 9 vss hvtnfet l=6e-08 w=1e-06 $X=18165 $Y=1115 $D=616
M19 9 pxcb_n vss vss hvtnfet l=6e-08 w=1e-06 $X=18165 $Y=1365 $D=616
M20 vss pxca_n 14 vss hvtnfet l=6e-08 w=1e-06 $X=24395 $Y=615 $D=616
M21 14 pxba_n vss vss hvtnfet l=6e-08 w=1e-06 $X=24395 $Y=865 $D=616
M22 vss pxba_n 14 vss hvtnfet l=6e-08 w=1e-06 $X=24395 $Y=1115 $D=616
M23 14 pxca_n vss vss hvtnfet l=6e-08 w=1e-06 $X=24395 $Y=1365 $D=616
M24 45 14 vss vss hvtnfet l=6e-08 w=2e-06 $X=26715 $Y=100 $D=616
M25 19 pxaa<3> 45 vss hvtnfet l=6e-08 w=2e-06 $X=26715 $Y=365 $D=616
M26 46 pxaa<2> 22 vss hvtnfet l=6e-08 w=2e-06 $X=26715 $Y=1615 $D=616
M27 vss 14 46 vss hvtnfet l=6e-08 w=2e-06 $X=26715 $Y=1880 $D=616
M28 47 pxaa<1> 20 vss hvtnfet l=6e-08 w=2e-06 $X=32355 $Y=615 $D=616
M29 vss 14 47 vss hvtnfet l=6e-08 w=2e-06 $X=32355 $Y=865 $D=616
M30 48 14 vss vss hvtnfet l=6e-08 w=2e-06 $X=32355 $Y=1115 $D=616
M31 48 pxaa<0> 21 vss hvtnfet l=6e-08 w=2e-06 $X=32355 $Y=1365 $D=616
M32 wla<3> 19 vss vss hvtnfet l=6e-08 w=2e-06 $X=36005 $Y=100 $D=616
M33 vss 19 wla<3> vss hvtnfet l=6e-08 w=2e-06 $X=36005 $Y=365 $D=616
M34 wla<1> 20 vss vss hvtnfet l=6e-08 w=2e-06 $X=36005 $Y=615 $D=616
M35 vss 20 wla<1> vss hvtnfet l=6e-08 w=2e-06 $X=36005 $Y=865 $D=616
M36 wla<0> 21 vss vss hvtnfet l=6e-08 w=2e-06 $X=36005 $Y=1115 $D=616
M37 vss 21 wla<0> vss hvtnfet l=6e-08 w=2e-06 $X=36005 $Y=1365 $D=616
M38 wla<2> 22 vss vss hvtnfet l=6e-08 w=2e-06 $X=36005 $Y=1615 $D=616
M39 vss 22 wla<2> vss hvtnfet l=6e-08 w=2e-06 $X=36005 $Y=1880 $D=616
M40 wlb<3> 1 vdd vdd hvtpfet l=6e-08 w=5e-06 $X=235 $Y=100 $D=636
M41 vdd 1 wlb<3> vdd hvtpfet l=6e-08 w=5e-06 $X=235 $Y=365 $D=636
M42 wlb<1> 2 vdd vdd hvtpfet l=6e-08 w=5e-06 $X=235 $Y=615 $D=636
M43 vdd 2 wlb<1> vdd hvtpfet l=6e-08 w=5e-06 $X=235 $Y=865 $D=636
M44 wlb<0> 3 vdd vdd hvtpfet l=6e-08 w=5e-06 $X=235 $Y=1115 $D=636
M45 vdd 3 wlb<0> vdd hvtpfet l=6e-08 w=5e-06 $X=235 $Y=1365 $D=636
M46 wlb<2> 4 vdd vdd hvtpfet l=6e-08 w=5e-06 $X=235 $Y=1615 $D=636
M47 vdd 4 wlb<2> vdd hvtpfet l=6e-08 w=5e-06 $X=235 $Y=1880 $D=636
M48 1 9 vdd vdd hvtpfet l=6e-08 w=2e-06 $X=11525 $Y=100 $D=636
M49 vdd pxab<3> 1 vdd hvtpfet l=6e-08 w=2e-06 $X=11525 $Y=365 $D=636
M50 2 pxab<1> vdd vdd hvtpfet l=6e-08 w=2e-06 $X=11525 $Y=615 $D=636
M51 vdd 9 2 vdd hvtpfet l=6e-08 w=2e-06 $X=11525 $Y=865 $D=636
M52 3 9 vdd vdd hvtpfet l=6e-08 w=2e-06 $X=11525 $Y=1115 $D=636
M53 vdd pxab<0> 3 vdd hvtpfet l=6e-08 w=2e-06 $X=11525 $Y=1365 $D=636
M54 4 pxab<2> vdd vdd hvtpfet l=6e-08 w=2e-06 $X=11525 $Y=1615 $D=636
M55 vdd 9 4 vdd hvtpfet l=6e-08 w=2e-06 $X=11525 $Y=1880 $D=636
M56 29 pxcb_n 9 vdd hvtpfet l=6e-08 w=2e-06 $X=19485 $Y=615 $D=636
M57 vdd pxbb_n 29 vdd hvtpfet l=6e-08 w=2e-06 $X=19485 $Y=865 $D=636
M58 29 pxbb_n vdd vdd hvtpfet l=6e-08 w=2e-06 $X=19485 $Y=1115 $D=636
M59 29 pxcb_n 9 vdd hvtpfet l=6e-08 w=2e-06 $X=19485 $Y=1365 $D=636
M60 30 pxca_n 14 vdd hvtpfet l=6e-08 w=2e-06 $X=22075 $Y=615 $D=636
M61 vdd pxba_n 30 vdd hvtpfet l=6e-08 w=2e-06 $X=22075 $Y=865 $D=636
M62 30 pxba_n vdd vdd hvtpfet l=6e-08 w=2e-06 $X=22075 $Y=1115 $D=636
M63 30 pxca_n 14 vdd hvtpfet l=6e-08 w=2e-06 $X=22075 $Y=1365 $D=636
M64 19 14 vdd vdd hvtpfet l=6e-08 w=2e-06 $X=30035 $Y=100 $D=636
M65 vdd pxaa<3> 19 vdd hvtpfet l=6e-08 w=2e-06 $X=30035 $Y=365 $D=636
M66 20 pxaa<1> vdd vdd hvtpfet l=6e-08 w=2e-06 $X=30035 $Y=615 $D=636
M67 vdd 14 20 vdd hvtpfet l=6e-08 w=2e-06 $X=30035 $Y=865 $D=636
M68 21 14 vdd vdd hvtpfet l=6e-08 w=2e-06 $X=30035 $Y=1115 $D=636
M69 vdd pxaa<0> 21 vdd hvtpfet l=6e-08 w=2e-06 $X=30035 $Y=1365 $D=636
M70 22 pxaa<2> vdd vdd hvtpfet l=6e-08 w=2e-06 $X=30035 $Y=1615 $D=636
M71 vdd 14 22 vdd hvtpfet l=6e-08 w=2e-06 $X=30035 $Y=1880 $D=636
M72 wla<3> 19 vdd vdd hvtpfet l=6e-08 w=5e-06 $X=38325 $Y=100 $D=636
M73 vdd 19 wla<3> vdd hvtpfet l=6e-08 w=5e-06 $X=38325 $Y=365 $D=636
M74 wla<1> 20 vdd vdd hvtpfet l=6e-08 w=5e-06 $X=38325 $Y=615 $D=636
M75 vdd 20 wla<1> vdd hvtpfet l=6e-08 w=5e-06 $X=38325 $Y=865 $D=636
M76 wla<0> 21 vdd vdd hvtpfet l=6e-08 w=5e-06 $X=38325 $Y=1115 $D=636
M77 vdd 21 wla<0> vdd hvtpfet l=6e-08 w=5e-06 $X=38325 $Y=1365 $D=636
M78 wla<2> 22 vdd vdd hvtpfet l=6e-08 w=5e-06 $X=38325 $Y=1615 $D=636
M79 vdd 22 wla<2> vdd hvtpfet l=6e-08 w=5e-06 $X=38325 $Y=1880 $D=636
.ends

************************************************************************
* Library Name: XMC55_DPS
* Cell Name:    xmc55_dps_xdec1_dummy_in
************************************************************************
.SUBCKT xmc55_dps_xdec1_dummy_in vdd vss
** N=606 EP=2 IP=0 FDC=8
M0 3 vdd vss vss hvtnfet l=6e-08 w=2e-06 $X=5555 $Y=100 $D=616
M1 4 vdd vss vss hvtnfet l=6e-08 w=2e-06 $X=14845 $Y=100 $D=616
M2 5 vdd vss vss hvtnfet l=6e-08 w=2e-06 $X=26715 $Y=100 $D=616
M3 6 vdd vss vss hvtnfet l=6e-08 w=2e-06 $X=36005 $Y=100 $D=616
M4 3 vdd vdd vdd hvtpfet l=6e-08 w=5e-06 $X=235 $Y=100 $D=636
M5 vdd vdd 4 vdd hvtpfet l=6e-08 w=2e-06 $X=11525 $Y=100 $D=636
M6 vdd vdd 5 vdd hvtpfet l=6e-08 w=2e-06 $X=30035 $Y=100 $D=636
M7 6 vdd vdd vdd hvtpfet l=6e-08 w=5e-06 $X=38325 $Y=100 $D=636
.ends

************************************************************************
* Library Name: XMC55_DPS
* Cell Name:    xmc55_dps_xdec1_dummy
************************************************************************
.SUBCKT xmc55_dps_xdec1_dummy vdd vss
** N=622 EP=2 IP=0 FDC=16
M0 3 vdd vss vss hvtnfet l=6e-08 w=2e-06 $X=5555 $Y=100 $D=616
M1 vss vdd 4 vss hvtnfet l=6e-08 w=2e-06 $X=5555 $Y=1160 $D=616
M2 5 vdd vss vss hvtnfet l=6e-08 w=2e-06 $X=14845 $Y=100 $D=616
M3 vss vdd 6 vss hvtnfet l=6e-08 w=2e-06 $X=14845 $Y=1160 $D=616
M4 7 vdd vss vss hvtnfet l=6e-08 w=2e-06 $X=26715 $Y=100 $D=616
M5 vss vdd 8 vss hvtnfet l=6e-08 w=2e-06 $X=26715 $Y=1160 $D=616
M6 9 vdd vss vss hvtnfet l=6e-08 w=2e-06 $X=36005 $Y=100 $D=616
M7 vss vdd 10 vss hvtnfet l=6e-08 w=2e-06 $X=36005 $Y=1160 $D=616
M8 3 vdd vdd vdd hvtpfet l=6e-08 w=5e-06 $X=235 $Y=100 $D=636
M9 vdd vdd 4 vdd hvtpfet l=6e-08 w=5e-06 $X=235 $Y=1160 $D=636
M10 vdd vdd 5 vdd hvtpfet l=6e-08 w=2e-06 $X=11525 $Y=100 $D=636
M11 vdd vdd 6 vdd hvtpfet l=6e-08 w=2e-06 $X=11525 $Y=1160 $D=636
M12 vdd vdd 7 vdd hvtpfet l=6e-08 w=2e-06 $X=30035 $Y=100 $D=636
M13 vdd vdd 8 vdd hvtpfet l=6e-08 w=2e-06 $X=30035 $Y=1160 $D=636
M14 9 vdd vdd vdd hvtpfet l=6e-08 w=5e-06 $X=38325 $Y=100 $D=636
M15 vdd vdd 10 vdd hvtpfet l=6e-08 w=5e-06 $X=38325 $Y=1160 $D=636
.ends

************************************************************************
* Library Name: XMC55_DPS
* Cell Name:    xmc55_dps_xdec1_dummy_out
************************************************************************
.SUBCKT xmc55_dps_xdec1_dummy_out vdd vss
** N=778 EP=2 IP=0 FDC=8
M0 2 vdd vss vss hvtnfet l=6e-08 w=2e-06 $X=5555 $Y=100 $D=616
M1 4 vdd vss vss hvtnfet l=6e-08 w=2e-06 $X=14845 $Y=100 $D=616
M2 5 vdd vss vss hvtnfet l=6e-08 w=2e-06 $X=26715 $Y=100 $D=616
M3 6 vdd vss vss hvtnfet l=6e-08 w=2e-06 $X=36005 $Y=100 $D=616
M4 2 vdd vdd vdd hvtpfet l=6e-08 w=5e-06 $X=235 $Y=100 $D=636
M5 vdd vdd 4 vdd hvtpfet l=6e-08 w=2e-06 $X=11525 $Y=100 $D=636
M6 vdd vdd 5 vdd hvtpfet l=6e-08 w=2e-06 $X=30035 $Y=100 $D=636
M7 6 vdd vdd vdd hvtpfet l=6e-08 w=5e-06 $X=38325 $Y=100 $D=636
.ends

************************************************************************
* Library Name: XMC55_DPS
* Cell Name:    CH974LP_dummy_rowx2
************************************************************************
.SUBCKT CH974LP_dummy_rowx2 blb blb_n gnd node wlb<1> wlb<0>
** N=55 EP=7 IP=0 FDC=6
M0 8 node gnd gnd srpddnfet l=6e-08 w=3.15e-07 $X=345 $Y=90 $D=778
M1 gnd node 9 gnd srpddnfet l=6e-08 w=3.15e-07 $X=345 $Y=870 $D=778
M2 blb wlb<0> node gnd srpgdnfet l=7.5e-08 w=1.05e-07 $X=130 $Y=345 $D=780
M3 blb wlb<1> node gnd srpgdnfet l=7.5e-08 w=1.05e-07 $X=130 $Y=600 $D=780
M4 blb_n wlb<0> 8 gnd srpgdnfet l=7.5e-08 w=1.05e-07 $X=430 $Y=345 $D=780
M5 9 wlb<1> blb_n gnd srpgdnfet l=7.5e-08 w=1.05e-07 $X=430 $Y=600 $D=780
.ends

************************************************************************
* Library Name: XMC55_DPS
* Cell Name:    CH974LP_bitcell_2x2
************************************************************************
.SUBCKT CH974LP_bitcell_2x2 bla<1> bla<0> bla_n<1> bla_n<0> blb<1> blb<0> 
+ blb_n<1> blb_n<0> gnd vdd wla<1> wla<0> wlb<1> wlb<0>
** N=185 EP=14 IP=0 FDC=32
M0 vdd 7 5 vdd srpudpfet l=7e-08 w=9e-08 $X=810 $Y=90 $D=776
M1 vdd 8 6 vdd srpudpfet l=7e-08 w=9e-08 $X=810 $Y=860 $D=776
M2 vdd 5 7 vdd srpudpfet l=7e-08 w=9e-08 $X=1010 $Y=350 $D=776
M3 vdd 6 8 vdd srpudpfet l=7e-08 w=9e-08 $X=1010 $Y=600 $D=776
M4 vdd 17 15 vdd srpudpfet l=7e-08 w=9e-08 $X=2720 $Y=350 $D=776
M5 vdd 18 16 vdd srpudpfet l=7e-08 w=9e-08 $X=2720 $Y=600 $D=776
M6 vdd 15 17 vdd srpudpfet l=7e-08 w=9e-08 $X=2920 $Y=90 $D=776
M7 vdd 16 18 vdd srpudpfet l=7e-08 w=9e-08 $X=2920 $Y=860 $D=776
M8 gnd 7 5 gnd srpddnfet l=6e-08 w=3.15e-07 $X=345 $Y=90 $D=778
M9 gnd 8 6 gnd srpddnfet l=6e-08 w=3.15e-07 $X=345 $Y=870 $D=778
M10 gnd 5 7 gnd srpddnfet l=6e-08 w=3.15e-07 $X=1250 $Y=360 $D=778
M11 gnd 6 8 gnd srpddnfet l=6e-08 w=3.15e-07 $X=1250 $Y=600 $D=778
M12 gnd 17 15 gnd srpddnfet l=6e-08 w=3.15e-07 $X=2255 $Y=360 $D=778
M13 gnd 18 16 gnd srpddnfet l=6e-08 w=3.15e-07 $X=2255 $Y=600 $D=778
M14 gnd 15 17 gnd srpddnfet l=6e-08 w=3.15e-07 $X=3160 $Y=90 $D=778
M15 gnd 16 18 gnd srpddnfet l=6e-08 w=3.15e-07 $X=3160 $Y=870 $D=778
M16 blb_n<1> wlb<0> 7 gnd srpgdnfet l=7.5e-08 w=1.05e-07 $X=130 $Y=345 $D=780
M17 blb_n<1> wlb<1> 8 gnd srpgdnfet l=7.5e-08 w=1.05e-07 $X=130 $Y=600 $D=780
M18 blb<1> wlb<0> 5 gnd srpgdnfet l=7.5e-08 w=1.05e-07 $X=430 $Y=345 $D=780
M19 6 wlb<1> blb<1> gnd srpgdnfet l=7.5e-08 w=1.05e-07 $X=430 $Y=600 $D=780
M20 7 wla<0> bla_n<1> gnd srpgdnfet l=7.5e-08 w=1.05e-07 $X=1375 $Y=90 $D=780
M21 bla_n<1> wla<1> 8 gnd srpgdnfet l=7.5e-08 w=1.05e-07 $X=1375 $Y=855 $D=780
M22 bla<1> wla<0> 5 gnd srpgdnfet l=7.5e-08 w=1.05e-07 $X=1675 $Y=90 $D=780
M23 bla<1> wla<1> 6 gnd srpgdnfet l=7.5e-08 w=1.05e-07 $X=1675 $Y=855 $D=780
M24 bla<0> wla<0> 17 gnd srpgdnfet l=7.5e-08 w=1.05e-07 $X=2040 $Y=90 $D=780
M25 bla<0> wla<1> 18 gnd srpgdnfet l=7.5e-08 w=1.05e-07 $X=2040 $Y=855 $D=780
M26 15 wla<0> bla_n<0> gnd srpgdnfet l=7.5e-08 w=1.05e-07 $X=2340 $Y=90 $D=780
M27 bla_n<0> wla<1> 16 gnd srpgdnfet l=7.5e-08 w=1.05e-07 $X=2340 $Y=855 $D=780
M28 blb<0> wlb<0> 17 gnd srpgdnfet l=7.5e-08 w=1.05e-07 $X=3285 $Y=345 $D=780
M29 18 wlb<1> blb<0> gnd srpgdnfet l=7.5e-08 w=1.05e-07 $X=3285 $Y=600 $D=780
M30 blb_n<0> wlb<0> 15 gnd srpgdnfet l=7.5e-08 w=1.05e-07 $X=3585 $Y=345 $D=780
M31 blb_n<0> wlb<1> 16 gnd srpgdnfet l=7.5e-08 w=1.05e-07 $X=3585 $Y=600 $D=780
.ends

************************************************************************

************************************************************************
* Cell Name:    dpram16x4096_AR_DUMMY_ROWX256
* View Name:    schematic
************************************************************************
.SUBCKT dpram16x4096_AR_DUMMY_ROWX256
+ BLB BLB_N GND NODE WLB<255> WLB<254> WLB<253> WLB<252> WLB<251> 
+ WLB<250> WLB<249> WLB<248> WLB<247> WLB<246> WLB<245> WLB<244> WLB<243> WLB<242> 
+ WLB<241> WLB<240> WLB<239> WLB<238> WLB<237> WLB<236> WLB<235> WLB<234> WLB<233> 
+ WLB<232> WLB<231> WLB<230> WLB<229> WLB<228> WLB<227> WLB<226> WLB<225> WLB<224> 
+ WLB<223> WLB<222> WLB<221> WLB<220> WLB<219> WLB<218> WLB<217> WLB<216> WLB<215> 
+ WLB<214> WLB<213> WLB<212> WLB<211> WLB<210> WLB<209> WLB<208> WLB<207> WLB<206> 
+ WLB<205> WLB<204> WLB<203> WLB<202> WLB<201> WLB<200> WLB<199> WLB<198> WLB<197> 
+ WLB<196> WLB<195> WLB<194> WLB<193> WLB<192> WLB<191> WLB<190> WLB<189> WLB<188> 
+ WLB<187> WLB<186> WLB<185> WLB<184> WLB<183> WLB<182> WLB<181> WLB<180> WLB<179> 
+ WLB<178> WLB<177> WLB<176> WLB<175> WLB<174> WLB<173> WLB<172> WLB<171> WLB<170> 
+ WLB<169> WLB<168> WLB<167> WLB<166> WLB<165> WLB<164> WLB<163> WLB<162> WLB<161> 
+ WLB<160> WLB<159> WLB<158> WLB<157> WLB<156> WLB<155> WLB<154> WLB<153> WLB<152> 
+ WLB<151> WLB<150> WLB<149> WLB<148> WLB<147> WLB<146> WLB<145> WLB<144> WLB<143> 
+ WLB<142> WLB<141> WLB<140> WLB<139> WLB<138> WLB<137> WLB<136> WLB<135> WLB<134> 
+ WLB<133> WLB<132> WLB<131> WLB<130> WLB<129> WLB<128> WLB<127> WLB<126> WLB<125> 
+ WLB<124> WLB<123> WLB<122> WLB<121> WLB<120> WLB<119> WLB<118> WLB<117> WLB<116> 
+ WLB<115> WLB<114> WLB<113> WLB<112> WLB<111> WLB<110> WLB<109> WLB<108> WLB<107> 
+ WLB<106> WLB<105> WLB<104> WLB<103> WLB<102> WLB<101> WLB<100> WLB<99> WLB<98> 
+ WLB<97> WLB<96> WLB<95> WLB<94> WLB<93> WLB<92> WLB<91> WLB<90> WLB<89> 
+ WLB<88> WLB<87> WLB<86> WLB<85> WLB<84> WLB<83> WLB<82> WLB<81> WLB<80> 
+ WLB<79> WLB<78> WLB<77> WLB<76> WLB<75> WLB<74> WLB<73> WLB<72> WLB<71> 
+ WLB<70> WLB<69> WLB<68> WLB<67> WLB<66> WLB<65> WLB<64> WLB<63> WLB<62> 
+ WLB<61> WLB<60> WLB<59> WLB<58> WLB<57> WLB<56> WLB<55> WLB<54> WLB<53> 
+ WLB<52> WLB<51> WLB<50> WLB<49> WLB<48> WLB<47> WLB<46> WLB<45> WLB<44> 
+ WLB<43> WLB<42> WLB<41> WLB<40> WLB<39> WLB<38> WLB<37> WLB<36> WLB<35> 
+ WLB<34> WLB<33> WLB<32> WLB<31> WLB<30> WLB<29> WLB<28> WLB<27> WLB<26> 
+ WLB<25> WLB<24> WLB<23> WLB<22> WLB<21> WLB<20> WLB<19> WLB<18> WLB<17> 
+ WLB<16> WLB<15> WLB<14> WLB<13> WLB<12> WLB<11> WLB<10> WLB<9> WLB<8> 
+ WLB<7> WLB<6> WLB<5> WLB<4> WLB<3> WLB<2> WLB<1> WLB<0> 
XBITCELLS<127>
+ BLB BLB_N GND NODE WLB<255> WLB<254>  / CH974LP_dummy_rowx2
XBITCELLS<126>
+ BLB BLB_N GND NODE WLB<253> WLB<252>  / CH974LP_dummy_rowx2
XBITCELLS<125>
+ BLB BLB_N GND NODE WLB<251> WLB<250>  / CH974LP_dummy_rowx2
XBITCELLS<124>
+ BLB BLB_N GND NODE WLB<249> WLB<248>  / CH974LP_dummy_rowx2
XBITCELLS<123>
+ BLB BLB_N GND NODE WLB<247> WLB<246>  / CH974LP_dummy_rowx2
XBITCELLS<122>
+ BLB BLB_N GND NODE WLB<245> WLB<244>  / CH974LP_dummy_rowx2
XBITCELLS<121>
+ BLB BLB_N GND NODE WLB<243> WLB<242>  / CH974LP_dummy_rowx2
XBITCELLS<120>
+ BLB BLB_N GND NODE WLB<241> WLB<240>  / CH974LP_dummy_rowx2
XBITCELLS<119>
+ BLB BLB_N GND NODE WLB<239> WLB<238>  / CH974LP_dummy_rowx2
XBITCELLS<118>
+ BLB BLB_N GND NODE WLB<237> WLB<236>  / CH974LP_dummy_rowx2
XBITCELLS<117>
+ BLB BLB_N GND NODE WLB<235> WLB<234>  / CH974LP_dummy_rowx2
XBITCELLS<116>
+ BLB BLB_N GND NODE WLB<233> WLB<232>  / CH974LP_dummy_rowx2
XBITCELLS<115>
+ BLB BLB_N GND NODE WLB<231> WLB<230>  / CH974LP_dummy_rowx2
XBITCELLS<114>
+ BLB BLB_N GND NODE WLB<229> WLB<228>  / CH974LP_dummy_rowx2
XBITCELLS<113>
+ BLB BLB_N GND NODE WLB<227> WLB<226>  / CH974LP_dummy_rowx2
XBITCELLS<112>
+ BLB BLB_N GND NODE WLB<225> WLB<224>  / CH974LP_dummy_rowx2
XBITCELLS<111>
+ BLB BLB_N GND NODE WLB<223> WLB<222>  / CH974LP_dummy_rowx2
XBITCELLS<110>
+ BLB BLB_N GND NODE WLB<221> WLB<220>  / CH974LP_dummy_rowx2
XBITCELLS<109>
+ BLB BLB_N GND NODE WLB<219> WLB<218>  / CH974LP_dummy_rowx2
XBITCELLS<108>
+ BLB BLB_N GND NODE WLB<217> WLB<216>  / CH974LP_dummy_rowx2
XBITCELLS<107>
+ BLB BLB_N GND NODE WLB<215> WLB<214>  / CH974LP_dummy_rowx2
XBITCELLS<106>
+ BLB BLB_N GND NODE WLB<213> WLB<212>  / CH974LP_dummy_rowx2
XBITCELLS<105>
+ BLB BLB_N GND NODE WLB<211> WLB<210>  / CH974LP_dummy_rowx2
XBITCELLS<104>
+ BLB BLB_N GND NODE WLB<209> WLB<208>  / CH974LP_dummy_rowx2
XBITCELLS<103>
+ BLB BLB_N GND NODE WLB<207> WLB<206>  / CH974LP_dummy_rowx2
XBITCELLS<102>
+ BLB BLB_N GND NODE WLB<205> WLB<204>  / CH974LP_dummy_rowx2
XBITCELLS<101>
+ BLB BLB_N GND NODE WLB<203> WLB<202>  / CH974LP_dummy_rowx2
XBITCELLS<100>
+ BLB BLB_N GND NODE WLB<201> WLB<200>  / CH974LP_dummy_rowx2
XBITCELLS<99>
+ BLB BLB_N GND NODE WLB<199> WLB<198>  / CH974LP_dummy_rowx2
XBITCELLS<98>
+ BLB BLB_N GND NODE WLB<197> WLB<196>  / CH974LP_dummy_rowx2
XBITCELLS<97>
+ BLB BLB_N GND NODE WLB<195> WLB<194>  / CH974LP_dummy_rowx2
XBITCELLS<96>
+ BLB BLB_N GND NODE WLB<193> WLB<192>  / CH974LP_dummy_rowx2
XBITCELLS<95>
+ BLB BLB_N GND NODE WLB<191> WLB<190>  / CH974LP_dummy_rowx2
XBITCELLS<94>
+ BLB BLB_N GND NODE WLB<189> WLB<188>  / CH974LP_dummy_rowx2
XBITCELLS<93>
+ BLB BLB_N GND NODE WLB<187> WLB<186>  / CH974LP_dummy_rowx2
XBITCELLS<92>
+ BLB BLB_N GND NODE WLB<185> WLB<184>  / CH974LP_dummy_rowx2
XBITCELLS<91>
+ BLB BLB_N GND NODE WLB<183> WLB<182>  / CH974LP_dummy_rowx2
XBITCELLS<90>
+ BLB BLB_N GND NODE WLB<181> WLB<180>  / CH974LP_dummy_rowx2
XBITCELLS<89>
+ BLB BLB_N GND NODE WLB<179> WLB<178>  / CH974LP_dummy_rowx2
XBITCELLS<88>
+ BLB BLB_N GND NODE WLB<177> WLB<176>  / CH974LP_dummy_rowx2
XBITCELLS<87>
+ BLB BLB_N GND NODE WLB<175> WLB<174>  / CH974LP_dummy_rowx2
XBITCELLS<86>
+ BLB BLB_N GND NODE WLB<173> WLB<172>  / CH974LP_dummy_rowx2
XBITCELLS<85>
+ BLB BLB_N GND NODE WLB<171> WLB<170>  / CH974LP_dummy_rowx2
XBITCELLS<84>
+ BLB BLB_N GND NODE WLB<169> WLB<168>  / CH974LP_dummy_rowx2
XBITCELLS<83>
+ BLB BLB_N GND NODE WLB<167> WLB<166>  / CH974LP_dummy_rowx2
XBITCELLS<82>
+ BLB BLB_N GND NODE WLB<165> WLB<164>  / CH974LP_dummy_rowx2
XBITCELLS<81>
+ BLB BLB_N GND NODE WLB<163> WLB<162>  / CH974LP_dummy_rowx2
XBITCELLS<80>
+ BLB BLB_N GND NODE WLB<161> WLB<160>  / CH974LP_dummy_rowx2
XBITCELLS<79>
+ BLB BLB_N GND NODE WLB<159> WLB<158>  / CH974LP_dummy_rowx2
XBITCELLS<78>
+ BLB BLB_N GND NODE WLB<157> WLB<156>  / CH974LP_dummy_rowx2
XBITCELLS<77>
+ BLB BLB_N GND NODE WLB<155> WLB<154>  / CH974LP_dummy_rowx2
XBITCELLS<76>
+ BLB BLB_N GND NODE WLB<153> WLB<152>  / CH974LP_dummy_rowx2
XBITCELLS<75>
+ BLB BLB_N GND NODE WLB<151> WLB<150>  / CH974LP_dummy_rowx2
XBITCELLS<74>
+ BLB BLB_N GND NODE WLB<149> WLB<148>  / CH974LP_dummy_rowx2
XBITCELLS<73>
+ BLB BLB_N GND NODE WLB<147> WLB<146>  / CH974LP_dummy_rowx2
XBITCELLS<72>
+ BLB BLB_N GND NODE WLB<145> WLB<144>  / CH974LP_dummy_rowx2
XBITCELLS<71>
+ BLB BLB_N GND NODE WLB<143> WLB<142>  / CH974LP_dummy_rowx2
XBITCELLS<70>
+ BLB BLB_N GND NODE WLB<141> WLB<140>  / CH974LP_dummy_rowx2
XBITCELLS<69>
+ BLB BLB_N GND NODE WLB<139> WLB<138>  / CH974LP_dummy_rowx2
XBITCELLS<68>
+ BLB BLB_N GND NODE WLB<137> WLB<136>  / CH974LP_dummy_rowx2
XBITCELLS<67>
+ BLB BLB_N GND NODE WLB<135> WLB<134>  / CH974LP_dummy_rowx2
XBITCELLS<66>
+ BLB BLB_N GND NODE WLB<133> WLB<132>  / CH974LP_dummy_rowx2
XBITCELLS<65>
+ BLB BLB_N GND NODE WLB<131> WLB<130>  / CH974LP_dummy_rowx2
XBITCELLS<64>
+ BLB BLB_N GND NODE WLB<129> WLB<128>  / CH974LP_dummy_rowx2
XBITCELLS<63>
+ BLB BLB_N GND NODE WLB<127> WLB<126>  / CH974LP_dummy_rowx2
XBITCELLS<62>
+ BLB BLB_N GND NODE WLB<125> WLB<124>  / CH974LP_dummy_rowx2
XBITCELLS<61>
+ BLB BLB_N GND NODE WLB<123> WLB<122>  / CH974LP_dummy_rowx2
XBITCELLS<60>
+ BLB BLB_N GND NODE WLB<121> WLB<120>  / CH974LP_dummy_rowx2
XBITCELLS<59>
+ BLB BLB_N GND NODE WLB<119> WLB<118>  / CH974LP_dummy_rowx2
XBITCELLS<58>
+ BLB BLB_N GND NODE WLB<117> WLB<116>  / CH974LP_dummy_rowx2
XBITCELLS<57>
+ BLB BLB_N GND NODE WLB<115> WLB<114>  / CH974LP_dummy_rowx2
XBITCELLS<56>
+ BLB BLB_N GND NODE WLB<113> WLB<112>  / CH974LP_dummy_rowx2
XBITCELLS<55>
+ BLB BLB_N GND NODE WLB<111> WLB<110>  / CH974LP_dummy_rowx2
XBITCELLS<54>
+ BLB BLB_N GND NODE WLB<109> WLB<108>  / CH974LP_dummy_rowx2
XBITCELLS<53>
+ BLB BLB_N GND NODE WLB<107> WLB<106>  / CH974LP_dummy_rowx2
XBITCELLS<52>
+ BLB BLB_N GND NODE WLB<105> WLB<104>  / CH974LP_dummy_rowx2
XBITCELLS<51>
+ BLB BLB_N GND NODE WLB<103> WLB<102>  / CH974LP_dummy_rowx2
XBITCELLS<50>
+ BLB BLB_N GND NODE WLB<101> WLB<100>  / CH974LP_dummy_rowx2
XBITCELLS<49>
+ BLB BLB_N GND NODE WLB<99> WLB<98>  / CH974LP_dummy_rowx2
XBITCELLS<48>
+ BLB BLB_N GND NODE WLB<97> WLB<96>  / CH974LP_dummy_rowx2
XBITCELLS<47>
+ BLB BLB_N GND NODE WLB<95> WLB<94>  / CH974LP_dummy_rowx2
XBITCELLS<46>
+ BLB BLB_N GND NODE WLB<93> WLB<92>  / CH974LP_dummy_rowx2
XBITCELLS<45>
+ BLB BLB_N GND NODE WLB<91> WLB<90>  / CH974LP_dummy_rowx2
XBITCELLS<44>
+ BLB BLB_N GND NODE WLB<89> WLB<88>  / CH974LP_dummy_rowx2
XBITCELLS<43>
+ BLB BLB_N GND NODE WLB<87> WLB<86>  / CH974LP_dummy_rowx2
XBITCELLS<42>
+ BLB BLB_N GND NODE WLB<85> WLB<84>  / CH974LP_dummy_rowx2
XBITCELLS<41>
+ BLB BLB_N GND NODE WLB<83> WLB<82>  / CH974LP_dummy_rowx2
XBITCELLS<40>
+ BLB BLB_N GND NODE WLB<81> WLB<80>  / CH974LP_dummy_rowx2
XBITCELLS<39>
+ BLB BLB_N GND NODE WLB<79> WLB<78>  / CH974LP_dummy_rowx2
XBITCELLS<38>
+ BLB BLB_N GND NODE WLB<77> WLB<76>  / CH974LP_dummy_rowx2
XBITCELLS<37>
+ BLB BLB_N GND NODE WLB<75> WLB<74>  / CH974LP_dummy_rowx2
XBITCELLS<36>
+ BLB BLB_N GND NODE WLB<73> WLB<72>  / CH974LP_dummy_rowx2
XBITCELLS<35>
+ BLB BLB_N GND NODE WLB<71> WLB<70>  / CH974LP_dummy_rowx2
XBITCELLS<34>
+ BLB BLB_N GND NODE WLB<69> WLB<68>  / CH974LP_dummy_rowx2
XBITCELLS<33>
+ BLB BLB_N GND NODE WLB<67> WLB<66>  / CH974LP_dummy_rowx2
XBITCELLS<32>
+ BLB BLB_N GND NODE WLB<65> WLB<64>  / CH974LP_dummy_rowx2
XBITCELLS<31>
+ BLB BLB_N GND NODE WLB<63> WLB<62>  / CH974LP_dummy_rowx2
XBITCELLS<30>
+ BLB BLB_N GND NODE WLB<61> WLB<60>  / CH974LP_dummy_rowx2
XBITCELLS<29>
+ BLB BLB_N GND NODE WLB<59> WLB<58>  / CH974LP_dummy_rowx2
XBITCELLS<28>
+ BLB BLB_N GND NODE WLB<57> WLB<56>  / CH974LP_dummy_rowx2
XBITCELLS<27>
+ BLB BLB_N GND NODE WLB<55> WLB<54>  / CH974LP_dummy_rowx2
XBITCELLS<26>
+ BLB BLB_N GND NODE WLB<53> WLB<52>  / CH974LP_dummy_rowx2
XBITCELLS<25>
+ BLB BLB_N GND NODE WLB<51> WLB<50>  / CH974LP_dummy_rowx2
XBITCELLS<24>
+ BLB BLB_N GND NODE WLB<49> WLB<48>  / CH974LP_dummy_rowx2
XBITCELLS<23>
+ BLB BLB_N GND NODE WLB<47> WLB<46>  / CH974LP_dummy_rowx2
XBITCELLS<22>
+ BLB BLB_N GND NODE WLB<45> WLB<44>  / CH974LP_dummy_rowx2
XBITCELLS<21>
+ BLB BLB_N GND NODE WLB<43> WLB<42>  / CH974LP_dummy_rowx2
XBITCELLS<20>
+ BLB BLB_N GND NODE WLB<41> WLB<40>  / CH974LP_dummy_rowx2
XBITCELLS<19>
+ BLB BLB_N GND NODE WLB<39> WLB<38>  / CH974LP_dummy_rowx2
XBITCELLS<18>
+ BLB BLB_N GND NODE WLB<37> WLB<36>  / CH974LP_dummy_rowx2
XBITCELLS<17>
+ BLB BLB_N GND NODE WLB<35> WLB<34>  / CH974LP_dummy_rowx2
XBITCELLS<16>
+ BLB BLB_N GND NODE WLB<33> WLB<32>  / CH974LP_dummy_rowx2
XBITCELLS<15>
+ BLB BLB_N GND NODE WLB<31> WLB<30>  / CH974LP_dummy_rowx2
XBITCELLS<14>
+ BLB BLB_N GND NODE WLB<29> WLB<28>  / CH974LP_dummy_rowx2
XBITCELLS<13>
+ BLB BLB_N GND NODE WLB<27> WLB<26>  / CH974LP_dummy_rowx2
XBITCELLS<12>
+ BLB BLB_N GND NODE WLB<25> WLB<24>  / CH974LP_dummy_rowx2
XBITCELLS<11>
+ BLB BLB_N GND NODE WLB<23> WLB<22>  / CH974LP_dummy_rowx2
XBITCELLS<10>
+ BLB BLB_N GND NODE WLB<21> WLB<20>  / CH974LP_dummy_rowx2
XBITCELLS<9>
+ BLB BLB_N GND NODE WLB<19> WLB<18>  / CH974LP_dummy_rowx2
XBITCELLS<8>
+ BLB BLB_N GND NODE WLB<17> WLB<16>  / CH974LP_dummy_rowx2
XBITCELLS<7>
+ BLB BLB_N GND NODE WLB<15> WLB<14>  / CH974LP_dummy_rowx2
XBITCELLS<6>
+ BLB BLB_N GND NODE WLB<13> WLB<12>  / CH974LP_dummy_rowx2
XBITCELLS<5>
+ BLB BLB_N GND NODE WLB<11> WLB<10>  / CH974LP_dummy_rowx2
XBITCELLS<4>
+ BLB BLB_N GND NODE WLB<9> WLB<8>  / CH974LP_dummy_rowx2
XBITCELLS<3>
+ BLB BLB_N GND NODE WLB<7> WLB<6>  / CH974LP_dummy_rowx2
XBITCELLS<2>
+ BLB BLB_N GND NODE WLB<5> WLB<4>  / CH974LP_dummy_rowx2
XBITCELLS<1>
+ BLB BLB_N GND NODE WLB<3> WLB<2>  / CH974LP_dummy_rowx2
XBITCELLS<0>
+ BLB BLB_N GND NODE WLB<1> WLB<0>  / CH974LP_dummy_rowx2
.ENDS

************************************************************************
* Cell Name:    dpram16x4096_COL2X8_EDGE_ROWX256
* View Name:    schematic
************************************************************************
.SUBCKT dpram16x4096_COL2X8_EDGE_ROWX256
+ B_WLB<255> B_WLB<254> B_WLB<253> B_WLB<252> B_WLB<251> B_WLB<250> B_WLB<249> B_WLB<248> B_WLB<247> 
+ B_WLB<246> B_WLB<245> B_WLB<244> B_WLB<243> B_WLB<242> B_WLB<241> B_WLB<240> B_WLB<239> B_WLB<238> 
+ B_WLB<237> B_WLB<236> B_WLB<235> B_WLB<234> B_WLB<233> B_WLB<232> B_WLB<231> B_WLB<230> B_WLB<229> 
+ B_WLB<228> B_WLB<227> B_WLB<226> B_WLB<225> B_WLB<224> B_WLB<223> B_WLB<222> B_WLB<221> B_WLB<220> 
+ B_WLB<219> B_WLB<218> B_WLB<217> B_WLB<216> B_WLB<215> B_WLB<214> B_WLB<213> B_WLB<212> B_WLB<211> 
+ B_WLB<210> B_WLB<209> B_WLB<208> B_WLB<207> B_WLB<206> B_WLB<205> B_WLB<204> B_WLB<203> B_WLB<202> 
+ B_WLB<201> B_WLB<200> B_WLB<199> B_WLB<198> B_WLB<197> B_WLB<196> B_WLB<195> B_WLB<194> B_WLB<193> 
+ B_WLB<192> B_WLB<191> B_WLB<190> B_WLB<189> B_WLB<188> B_WLB<187> B_WLB<186> B_WLB<185> B_WLB<184> 
+ B_WLB<183> B_WLB<182> B_WLB<181> B_WLB<180> B_WLB<179> B_WLB<178> B_WLB<177> B_WLB<176> B_WLB<175> 
+ B_WLB<174> B_WLB<173> B_WLB<172> B_WLB<171> B_WLB<170> B_WLB<169> B_WLB<168> B_WLB<167> B_WLB<166> 
+ B_WLB<165> B_WLB<164> B_WLB<163> B_WLB<162> B_WLB<161> B_WLB<160> B_WLB<159> B_WLB<158> B_WLB<157> 
+ B_WLB<156> B_WLB<155> B_WLB<154> B_WLB<153> B_WLB<152> B_WLB<151> B_WLB<150> B_WLB<149> B_WLB<148> 
+ B_WLB<147> B_WLB<146> B_WLB<145> B_WLB<144> B_WLB<143> B_WLB<142> B_WLB<141> B_WLB<140> B_WLB<139> 
+ B_WLB<138> B_WLB<137> B_WLB<136> B_WLB<135> B_WLB<134> B_WLB<133> B_WLB<132> B_WLB<131> B_WLB<130> 
+ B_WLB<129> B_WLB<128> B_WLB<127> B_WLB<126> B_WLB<125> B_WLB<124> B_WLB<123> B_WLB<122> B_WLB<121> 
+ B_WLB<120> B_WLB<119> B_WLB<118> B_WLB<117> B_WLB<116> B_WLB<115> B_WLB<114> B_WLB<113> B_WLB<112> 
+ B_WLB<111> B_WLB<110> B_WLB<109> B_WLB<108> B_WLB<107> B_WLB<106> B_WLB<105> B_WLB<104> B_WLB<103> 
+ B_WLB<102> B_WLB<101> B_WLB<100> B_WLB<99> B_WLB<98> B_WLB<97> B_WLB<96> B_WLB<95> B_WLB<94> 
+ B_WLB<93> B_WLB<92> B_WLB<91> B_WLB<90> B_WLB<89> B_WLB<88> B_WLB<87> B_WLB<86> B_WLB<85> 
+ B_WLB<84> B_WLB<83> B_WLB<82> B_WLB<81> B_WLB<80> B_WLB<79> B_WLB<78> B_WLB<77> B_WLB<76> 
+ B_WLB<75> B_WLB<74> B_WLB<73> B_WLB<72> B_WLB<71> B_WLB<70> B_WLB<69> B_WLB<68> B_WLB<67> 
+ B_WLB<66> B_WLB<65> B_WLB<64> B_WLB<63> B_WLB<62> B_WLB<61> B_WLB<60> B_WLB<59> B_WLB<58> 
+ B_WLB<57> B_WLB<56> B_WLB<55> B_WLB<54> B_WLB<53> B_WLB<52> B_WLB<51> B_WLB<50> B_WLB<49> 
+ B_WLB<48> B_WLB<47> B_WLB<46> B_WLB<45> B_WLB<44> B_WLB<43> B_WLB<42> B_WLB<41> B_WLB<40> 
+ B_WLB<39> B_WLB<38> B_WLB<37> B_WLB<36> B_WLB<35> B_WLB<34> B_WLB<33> B_WLB<32> B_WLB<31> 
+ B_WLB<30> B_WLB<29> B_WLB<28> B_WLB<27> B_WLB<26> B_WLB<25> B_WLB<24> B_WLB<23> B_WLB<22> 
+ B_WLB<21> B_WLB<20> B_WLB<19> B_WLB<18> B_WLB<17> B_WLB<16> B_WLB<15> B_WLB<14> B_WLB<13> 
+ B_WLB<12> B_WLB<11> B_WLB<10> B_WLB<9> B_WLB<8> B_WLB<7> B_WLB<6> B_WLB<5> B_WLB<4> 
+ B_WLB<3> B_WLB<2> B_WLB<1> B_WLB<0> T_WLB<255> T_WLB<254> T_WLB<253> T_WLB<252> T_WLB<251> 
+ T_WLB<250> T_WLB<249> T_WLB<248> T_WLB<247> T_WLB<246> T_WLB<245> T_WLB<244> T_WLB<243> T_WLB<242> 
+ T_WLB<241> T_WLB<240> T_WLB<239> T_WLB<238> T_WLB<237> T_WLB<236> T_WLB<235> T_WLB<234> T_WLB<233> 
+ T_WLB<232> T_WLB<231> T_WLB<230> T_WLB<229> T_WLB<228> T_WLB<227> T_WLB<226> T_WLB<225> T_WLB<224> 
+ T_WLB<223> T_WLB<222> T_WLB<221> T_WLB<220> T_WLB<219> T_WLB<218> T_WLB<217> T_WLB<216> T_WLB<215> 
+ T_WLB<214> T_WLB<213> T_WLB<212> T_WLB<211> T_WLB<210> T_WLB<209> T_WLB<208> T_WLB<207> T_WLB<206> 
+ T_WLB<205> T_WLB<204> T_WLB<203> T_WLB<202> T_WLB<201> T_WLB<200> T_WLB<199> T_WLB<198> T_WLB<197> 
+ T_WLB<196> T_WLB<195> T_WLB<194> T_WLB<193> T_WLB<192> T_WLB<191> T_WLB<190> T_WLB<189> T_WLB<188> 
+ T_WLB<187> T_WLB<186> T_WLB<185> T_WLB<184> T_WLB<183> T_WLB<182> T_WLB<181> T_WLB<180> T_WLB<179> 
+ T_WLB<178> T_WLB<177> T_WLB<176> T_WLB<175> T_WLB<174> T_WLB<173> T_WLB<172> T_WLB<171> T_WLB<170> 
+ T_WLB<169> T_WLB<168> T_WLB<167> T_WLB<166> T_WLB<165> T_WLB<164> T_WLB<163> T_WLB<162> T_WLB<161> 
+ T_WLB<160> T_WLB<159> T_WLB<158> T_WLB<157> T_WLB<156> T_WLB<155> T_WLB<154> T_WLB<153> T_WLB<152> 
+ T_WLB<151> T_WLB<150> T_WLB<149> T_WLB<148> T_WLB<147> T_WLB<146> T_WLB<145> T_WLB<144> T_WLB<143> 
+ T_WLB<142> T_WLB<141> T_WLB<140> T_WLB<139> T_WLB<138> T_WLB<137> T_WLB<136> T_WLB<135> T_WLB<134> 
+ T_WLB<133> T_WLB<132> T_WLB<131> T_WLB<130> T_WLB<129> T_WLB<128> T_WLB<127> T_WLB<126> T_WLB<125> 
+ T_WLB<124> T_WLB<123> T_WLB<122> T_WLB<121> T_WLB<120> T_WLB<119> T_WLB<118> T_WLB<117> T_WLB<116> 
+ T_WLB<115> T_WLB<114> T_WLB<113> T_WLB<112> T_WLB<111> T_WLB<110> T_WLB<109> T_WLB<108> T_WLB<107> 
+ T_WLB<106> T_WLB<105> T_WLB<104> T_WLB<103> T_WLB<102> T_WLB<101> T_WLB<100> T_WLB<99> T_WLB<98> 
+ T_WLB<97> T_WLB<96> T_WLB<95> T_WLB<94> T_WLB<93> T_WLB<92> T_WLB<91> T_WLB<90> T_WLB<89> 
+ T_WLB<88> T_WLB<87> T_WLB<86> T_WLB<85> T_WLB<84> T_WLB<83> T_WLB<82> T_WLB<81> T_WLB<80> 
+ T_WLB<79> T_WLB<78> T_WLB<77> T_WLB<76> T_WLB<75> T_WLB<74> T_WLB<73> T_WLB<72> T_WLB<71> 
+ T_WLB<70> T_WLB<69> T_WLB<68> T_WLB<67> T_WLB<66> T_WLB<65> T_WLB<64> T_WLB<63> T_WLB<62> 
+ T_WLB<61> T_WLB<60> T_WLB<59> T_WLB<58> T_WLB<57> T_WLB<56> T_WLB<55> T_WLB<54> T_WLB<53> 
+ T_WLB<52> T_WLB<51> T_WLB<50> T_WLB<49> T_WLB<48> T_WLB<47> T_WLB<46> T_WLB<45> T_WLB<44> 
+ T_WLB<43> T_WLB<42> T_WLB<41> T_WLB<40> T_WLB<39> T_WLB<38> T_WLB<37> T_WLB<36> T_WLB<35> 
+ T_WLB<34> T_WLB<33> T_WLB<32> T_WLB<31> T_WLB<30> T_WLB<29> T_WLB<28> T_WLB<27> T_WLB<26> 
+ T_WLB<25> T_WLB<24> T_WLB<23> T_WLB<22> T_WLB<21> T_WLB<20> T_WLB<19> T_WLB<18> T_WLB<17> 
+ T_WLB<16> T_WLB<15> T_WLB<14> T_WLB<13> T_WLB<12> T_WLB<11> T_WLB<10> T_WLB<9> T_WLB<8> 
+ T_WLB<7> T_WLB<6> T_WLB<5> T_WLB<4> T_WLB<3> T_WLB<2> T_WLB<1> T_WLB<0> TIE_LOW 
+ VDD VSS 
XCOL
+ NET14 VDD VSS  / xmc55_dps_localc8io_edge
XAR_TOP
+ VSS VSS VSS VSS T_WLB<255> T_WLB<254> T_WLB<253> T_WLB<252> T_WLB<251> 
+ T_WLB<250> T_WLB<249> T_WLB<248> T_WLB<247> T_WLB<246> T_WLB<245> T_WLB<244> T_WLB<243> T_WLB<242> 
+ T_WLB<241> T_WLB<240> T_WLB<239> T_WLB<238> T_WLB<237> T_WLB<236> T_WLB<235> T_WLB<234> T_WLB<233> 
+ T_WLB<232> T_WLB<231> T_WLB<230> T_WLB<229> T_WLB<228> T_WLB<227> T_WLB<226> T_WLB<225> T_WLB<224> 
+ T_WLB<223> T_WLB<222> T_WLB<221> T_WLB<220> T_WLB<219> T_WLB<218> T_WLB<217> T_WLB<216> T_WLB<215> 
+ T_WLB<214> T_WLB<213> T_WLB<212> T_WLB<211> T_WLB<210> T_WLB<209> T_WLB<208> T_WLB<207> T_WLB<206> 
+ T_WLB<205> T_WLB<204> T_WLB<203> T_WLB<202> T_WLB<201> T_WLB<200> T_WLB<199> T_WLB<198> T_WLB<197> 
+ T_WLB<196> T_WLB<195> T_WLB<194> T_WLB<193> T_WLB<192> T_WLB<191> T_WLB<190> T_WLB<189> T_WLB<188> 
+ T_WLB<187> T_WLB<186> T_WLB<185> T_WLB<184> T_WLB<183> T_WLB<182> T_WLB<181> T_WLB<180> T_WLB<179> 
+ T_WLB<178> T_WLB<177> T_WLB<176> T_WLB<175> T_WLB<174> T_WLB<173> T_WLB<172> T_WLB<171> T_WLB<170> 
+ T_WLB<169> T_WLB<168> T_WLB<167> T_WLB<166> T_WLB<165> T_WLB<164> T_WLB<163> T_WLB<162> T_WLB<161> 
+ T_WLB<160> T_WLB<159> T_WLB<158> T_WLB<157> T_WLB<156> T_WLB<155> T_WLB<154> T_WLB<153> T_WLB<152> 
+ T_WLB<151> T_WLB<150> T_WLB<149> T_WLB<148> T_WLB<147> T_WLB<146> T_WLB<145> T_WLB<144> T_WLB<143> 
+ T_WLB<142> T_WLB<141> T_WLB<140> T_WLB<139> T_WLB<138> T_WLB<137> T_WLB<136> T_WLB<135> T_WLB<134> 
+ T_WLB<133> T_WLB<132> T_WLB<131> T_WLB<130> T_WLB<129> T_WLB<128> T_WLB<127> T_WLB<126> T_WLB<125> 
+ T_WLB<124> T_WLB<123> T_WLB<122> T_WLB<121> T_WLB<120> T_WLB<119> T_WLB<118> T_WLB<117> T_WLB<116> 
+ T_WLB<115> T_WLB<114> T_WLB<113> T_WLB<112> T_WLB<111> T_WLB<110> T_WLB<109> T_WLB<108> T_WLB<107> 
+ T_WLB<106> T_WLB<105> T_WLB<104> T_WLB<103> T_WLB<102> T_WLB<101> T_WLB<100> T_WLB<99> T_WLB<98> 
+ T_WLB<97> T_WLB<96> T_WLB<95> T_WLB<94> T_WLB<93> T_WLB<92> T_WLB<91> T_WLB<90> T_WLB<89> 
+ T_WLB<88> T_WLB<87> T_WLB<86> T_WLB<85> T_WLB<84> T_WLB<83> T_WLB<82> T_WLB<81> T_WLB<80> 
+ T_WLB<79> T_WLB<78> T_WLB<77> T_WLB<76> T_WLB<75> T_WLB<74> T_WLB<73> T_WLB<72> T_WLB<71> 
+ T_WLB<70> T_WLB<69> T_WLB<68> T_WLB<67> T_WLB<66> T_WLB<65> T_WLB<64> T_WLB<63> T_WLB<62> 
+ T_WLB<61> T_WLB<60> T_WLB<59> T_WLB<58> T_WLB<57> T_WLB<56> T_WLB<55> T_WLB<54> T_WLB<53> 
+ T_WLB<52> T_WLB<51> T_WLB<50> T_WLB<49> T_WLB<48> T_WLB<47> T_WLB<46> T_WLB<45> T_WLB<44> 
+ T_WLB<43> T_WLB<42> T_WLB<41> T_WLB<40> T_WLB<39> T_WLB<38> T_WLB<37> T_WLB<36> T_WLB<35> 
+ T_WLB<34> T_WLB<33> T_WLB<32> T_WLB<31> T_WLB<30> T_WLB<29> T_WLB<28> T_WLB<27> T_WLB<26> 
+ T_WLB<25> T_WLB<24> T_WLB<23> T_WLB<22> T_WLB<21> T_WLB<20> T_WLB<19> T_WLB<18> T_WLB<17> 
+ T_WLB<16> T_WLB<15> T_WLB<14> T_WLB<13> T_WLB<12> T_WLB<11> T_WLB<10> T_WLB<9> T_WLB<8> 
+ T_WLB<7> T_WLB<6> T_WLB<5> T_WLB<4> T_WLB<3> T_WLB<2> T_WLB<1> T_WLB<0>  / dpram16x4096_AR_DUMMY_ROWX256
XAR_BOT
+ VSS VSS VSS VSS B_WLB<255> B_WLB<254> B_WLB<253> B_WLB<252> B_WLB<251> 
+ B_WLB<250> B_WLB<249> B_WLB<248> B_WLB<247> B_WLB<246> B_WLB<245> B_WLB<244> B_WLB<243> B_WLB<242> 
+ B_WLB<241> B_WLB<240> B_WLB<239> B_WLB<238> B_WLB<237> B_WLB<236> B_WLB<235> B_WLB<234> B_WLB<233> 
+ B_WLB<232> B_WLB<231> B_WLB<230> B_WLB<229> B_WLB<228> B_WLB<227> B_WLB<226> B_WLB<225> B_WLB<224> 
+ B_WLB<223> B_WLB<222> B_WLB<221> B_WLB<220> B_WLB<219> B_WLB<218> B_WLB<217> B_WLB<216> B_WLB<215> 
+ B_WLB<214> B_WLB<213> B_WLB<212> B_WLB<211> B_WLB<210> B_WLB<209> B_WLB<208> B_WLB<207> B_WLB<206> 
+ B_WLB<205> B_WLB<204> B_WLB<203> B_WLB<202> B_WLB<201> B_WLB<200> B_WLB<199> B_WLB<198> B_WLB<197> 
+ B_WLB<196> B_WLB<195> B_WLB<194> B_WLB<193> B_WLB<192> B_WLB<191> B_WLB<190> B_WLB<189> B_WLB<188> 
+ B_WLB<187> B_WLB<186> B_WLB<185> B_WLB<184> B_WLB<183> B_WLB<182> B_WLB<181> B_WLB<180> B_WLB<179> 
+ B_WLB<178> B_WLB<177> B_WLB<176> B_WLB<175> B_WLB<174> B_WLB<173> B_WLB<172> B_WLB<171> B_WLB<170> 
+ B_WLB<169> B_WLB<168> B_WLB<167> B_WLB<166> B_WLB<165> B_WLB<164> B_WLB<163> B_WLB<162> B_WLB<161> 
+ B_WLB<160> B_WLB<159> B_WLB<158> B_WLB<157> B_WLB<156> B_WLB<155> B_WLB<154> B_WLB<153> B_WLB<152> 
+ B_WLB<151> B_WLB<150> B_WLB<149> B_WLB<148> B_WLB<147> B_WLB<146> B_WLB<145> B_WLB<144> B_WLB<143> 
+ B_WLB<142> B_WLB<141> B_WLB<140> B_WLB<139> B_WLB<138> B_WLB<137> B_WLB<136> B_WLB<135> B_WLB<134> 
+ B_WLB<133> B_WLB<132> B_WLB<131> B_WLB<130> B_WLB<129> B_WLB<128> B_WLB<127> B_WLB<126> B_WLB<125> 
+ B_WLB<124> B_WLB<123> B_WLB<122> B_WLB<121> B_WLB<120> B_WLB<119> B_WLB<118> B_WLB<117> B_WLB<116> 
+ B_WLB<115> B_WLB<114> B_WLB<113> B_WLB<112> B_WLB<111> B_WLB<110> B_WLB<109> B_WLB<108> B_WLB<107> 
+ B_WLB<106> B_WLB<105> B_WLB<104> B_WLB<103> B_WLB<102> B_WLB<101> B_WLB<100> B_WLB<99> B_WLB<98> 
+ B_WLB<97> B_WLB<96> B_WLB<95> B_WLB<94> B_WLB<93> B_WLB<92> B_WLB<91> B_WLB<90> B_WLB<89> 
+ B_WLB<88> B_WLB<87> B_WLB<86> B_WLB<85> B_WLB<84> B_WLB<83> B_WLB<82> B_WLB<81> B_WLB<80> 
+ B_WLB<79> B_WLB<78> B_WLB<77> B_WLB<76> B_WLB<75> B_WLB<74> B_WLB<73> B_WLB<72> B_WLB<71> 
+ B_WLB<70> B_WLB<69> B_WLB<68> B_WLB<67> B_WLB<66> B_WLB<65> B_WLB<64> B_WLB<63> B_WLB<62> 
+ B_WLB<61> B_WLB<60> B_WLB<59> B_WLB<58> B_WLB<57> B_WLB<56> B_WLB<55> B_WLB<54> B_WLB<53> 
+ B_WLB<52> B_WLB<51> B_WLB<50> B_WLB<49> B_WLB<48> B_WLB<47> B_WLB<46> B_WLB<45> B_WLB<44> 
+ B_WLB<43> B_WLB<42> B_WLB<41> B_WLB<40> B_WLB<39> B_WLB<38> B_WLB<37> B_WLB<36> B_WLB<35> 
+ B_WLB<34> B_WLB<33> B_WLB<32> B_WLB<31> B_WLB<30> B_WLB<29> B_WLB<28> B_WLB<27> B_WLB<26> 
+ B_WLB<25> B_WLB<24> B_WLB<23> B_WLB<22> B_WLB<21> B_WLB<20> B_WLB<19> B_WLB<18> B_WLB<17> 
+ B_WLB<16> B_WLB<15> B_WLB<14> B_WLB<13> B_WLB<12> B_WLB<11> B_WLB<10> B_WLB<9> B_WLB<8> 
+ B_WLB<7> B_WLB<6> B_WLB<5> B_WLB<4> B_WLB<3> B_WLB<2> B_WLB<1> B_WLB<0>  / dpram16x4096_AR_DUMMY_ROWX256
XBUF0
+ TIE_LOW VDD VSS  / xmc55_dps_collar_edge
.ENDS

************************************************************************
* Cell Name:    dpram16x4096_COL2X8_DUM_ROWX256
* View Name:    schematic
************************************************************************
.SUBCKT dpram16x4096_COL2X8_DUM_ROWX256
+ B_WLB<255> B_WLB<254> B_WLB<253> B_WLB<252> B_WLB<251> B_WLB<250> B_WLB<249> B_WLB<248> B_WLB<247> 
+ B_WLB<246> B_WLB<245> B_WLB<244> B_WLB<243> B_WLB<242> B_WLB<241> B_WLB<240> B_WLB<239> B_WLB<238> 
+ B_WLB<237> B_WLB<236> B_WLB<235> B_WLB<234> B_WLB<233> B_WLB<232> B_WLB<231> B_WLB<230> B_WLB<229> 
+ B_WLB<228> B_WLB<227> B_WLB<226> B_WLB<225> B_WLB<224> B_WLB<223> B_WLB<222> B_WLB<221> B_WLB<220> 
+ B_WLB<219> B_WLB<218> B_WLB<217> B_WLB<216> B_WLB<215> B_WLB<214> B_WLB<213> B_WLB<212> B_WLB<211> 
+ B_WLB<210> B_WLB<209> B_WLB<208> B_WLB<207> B_WLB<206> B_WLB<205> B_WLB<204> B_WLB<203> B_WLB<202> 
+ B_WLB<201> B_WLB<200> B_WLB<199> B_WLB<198> B_WLB<197> B_WLB<196> B_WLB<195> B_WLB<194> B_WLB<193> 
+ B_WLB<192> B_WLB<191> B_WLB<190> B_WLB<189> B_WLB<188> B_WLB<187> B_WLB<186> B_WLB<185> B_WLB<184> 
+ B_WLB<183> B_WLB<182> B_WLB<181> B_WLB<180> B_WLB<179> B_WLB<178> B_WLB<177> B_WLB<176> B_WLB<175> 
+ B_WLB<174> B_WLB<173> B_WLB<172> B_WLB<171> B_WLB<170> B_WLB<169> B_WLB<168> B_WLB<167> B_WLB<166> 
+ B_WLB<165> B_WLB<164> B_WLB<163> B_WLB<162> B_WLB<161> B_WLB<160> B_WLB<159> B_WLB<158> B_WLB<157> 
+ B_WLB<156> B_WLB<155> B_WLB<154> B_WLB<153> B_WLB<152> B_WLB<151> B_WLB<150> B_WLB<149> B_WLB<148> 
+ B_WLB<147> B_WLB<146> B_WLB<145> B_WLB<144> B_WLB<143> B_WLB<142> B_WLB<141> B_WLB<140> B_WLB<139> 
+ B_WLB<138> B_WLB<137> B_WLB<136> B_WLB<135> B_WLB<134> B_WLB<133> B_WLB<132> B_WLB<131> B_WLB<130> 
+ B_WLB<129> B_WLB<128> B_WLB<127> B_WLB<126> B_WLB<125> B_WLB<124> B_WLB<123> B_WLB<122> B_WLB<121> 
+ B_WLB<120> B_WLB<119> B_WLB<118> B_WLB<117> B_WLB<116> B_WLB<115> B_WLB<114> B_WLB<113> B_WLB<112> 
+ B_WLB<111> B_WLB<110> B_WLB<109> B_WLB<108> B_WLB<107> B_WLB<106> B_WLB<105> B_WLB<104> B_WLB<103> 
+ B_WLB<102> B_WLB<101> B_WLB<100> B_WLB<99> B_WLB<98> B_WLB<97> B_WLB<96> B_WLB<95> B_WLB<94> 
+ B_WLB<93> B_WLB<92> B_WLB<91> B_WLB<90> B_WLB<89> B_WLB<88> B_WLB<87> B_WLB<86> B_WLB<85> 
+ B_WLB<84> B_WLB<83> B_WLB<82> B_WLB<81> B_WLB<80> B_WLB<79> B_WLB<78> B_WLB<77> B_WLB<76> 
+ B_WLB<75> B_WLB<74> B_WLB<73> B_WLB<72> B_WLB<71> B_WLB<70> B_WLB<69> B_WLB<68> B_WLB<67> 
+ B_WLB<66> B_WLB<65> B_WLB<64> B_WLB<63> B_WLB<62> B_WLB<61> B_WLB<60> B_WLB<59> B_WLB<58> 
+ B_WLB<57> B_WLB<56> B_WLB<55> B_WLB<54> B_WLB<53> B_WLB<52> B_WLB<51> B_WLB<50> B_WLB<49> 
+ B_WLB<48> B_WLB<47> B_WLB<46> B_WLB<45> B_WLB<44> B_WLB<43> B_WLB<42> B_WLB<41> B_WLB<40> 
+ B_WLB<39> B_WLB<38> B_WLB<37> B_WLB<36> B_WLB<35> B_WLB<34> B_WLB<33> B_WLB<32> B_WLB<31> 
+ B_WLB<30> B_WLB<29> B_WLB<28> B_WLB<27> B_WLB<26> B_WLB<25> B_WLB<24> B_WLB<23> B_WLB<22> 
+ B_WLB<21> B_WLB<20> B_WLB<19> B_WLB<18> B_WLB<17> B_WLB<16> B_WLB<15> B_WLB<14> B_WLB<13> 
+ B_WLB<12> B_WLB<11> B_WLB<10> B_WLB<9> B_WLB<8> B_WLB<7> B_WLB<6> B_WLB<5> B_WLB<4> 
+ B_WLB<3> B_WLB<2> B_WLB<1> B_WLB<0> DBL_PD_N<3> DBL_PD_N<2> DBL_PD_N<1> DBL_PD_N<0> DWL<1> 
+ DWL<0> STCLK T_WLB<255> T_WLB<254> T_WLB<253> T_WLB<252> T_WLB<251> T_WLB<250> T_WLB<249> 
+ T_WLB<248> T_WLB<247> T_WLB<246> T_WLB<245> T_WLB<244> T_WLB<243> T_WLB<242> T_WLB<241> T_WLB<240> 
+ T_WLB<239> T_WLB<238> T_WLB<237> T_WLB<236> T_WLB<235> T_WLB<234> T_WLB<233> T_WLB<232> T_WLB<231> 
+ T_WLB<230> T_WLB<229> T_WLB<228> T_WLB<227> T_WLB<226> T_WLB<225> T_WLB<224> T_WLB<223> T_WLB<222> 
+ T_WLB<221> T_WLB<220> T_WLB<219> T_WLB<218> T_WLB<217> T_WLB<216> T_WLB<215> T_WLB<214> T_WLB<213> 
+ T_WLB<212> T_WLB<211> T_WLB<210> T_WLB<209> T_WLB<208> T_WLB<207> T_WLB<206> T_WLB<205> T_WLB<204> 
+ T_WLB<203> T_WLB<202> T_WLB<201> T_WLB<200> T_WLB<199> T_WLB<198> T_WLB<197> T_WLB<196> T_WLB<195> 
+ T_WLB<194> T_WLB<193> T_WLB<192> T_WLB<191> T_WLB<190> T_WLB<189> T_WLB<188> T_WLB<187> T_WLB<186> 
+ T_WLB<185> T_WLB<184> T_WLB<183> T_WLB<182> T_WLB<181> T_WLB<180> T_WLB<179> T_WLB<178> T_WLB<177> 
+ T_WLB<176> T_WLB<175> T_WLB<174> T_WLB<173> T_WLB<172> T_WLB<171> T_WLB<170> T_WLB<169> T_WLB<168> 
+ T_WLB<167> T_WLB<166> T_WLB<165> T_WLB<164> T_WLB<163> T_WLB<162> T_WLB<161> T_WLB<160> T_WLB<159> 
+ T_WLB<158> T_WLB<157> T_WLB<156> T_WLB<155> T_WLB<154> T_WLB<153> T_WLB<152> T_WLB<151> T_WLB<150> 
+ T_WLB<149> T_WLB<148> T_WLB<147> T_WLB<146> T_WLB<145> T_WLB<144> T_WLB<143> T_WLB<142> T_WLB<141> 
+ T_WLB<140> T_WLB<139> T_WLB<138> T_WLB<137> T_WLB<136> T_WLB<135> T_WLB<134> T_WLB<133> T_WLB<132> 
+ T_WLB<131> T_WLB<130> T_WLB<129> T_WLB<128> T_WLB<127> T_WLB<126> T_WLB<125> T_WLB<124> T_WLB<123> 
+ T_WLB<122> T_WLB<121> T_WLB<120> T_WLB<119> T_WLB<118> T_WLB<117> T_WLB<116> T_WLB<115> T_WLB<114> 
+ T_WLB<113> T_WLB<112> T_WLB<111> T_WLB<110> T_WLB<109> T_WLB<108> T_WLB<107> T_WLB<106> T_WLB<105> 
+ T_WLB<104> T_WLB<103> T_WLB<102> T_WLB<101> T_WLB<100> T_WLB<99> T_WLB<98> T_WLB<97> T_WLB<96> 
+ T_WLB<95> T_WLB<94> T_WLB<93> T_WLB<92> T_WLB<91> T_WLB<90> T_WLB<89> T_WLB<88> T_WLB<87> 
+ T_WLB<86> T_WLB<85> T_WLB<84> T_WLB<83> T_WLB<82> T_WLB<81> T_WLB<80> T_WLB<79> T_WLB<78> 
+ T_WLB<77> T_WLB<76> T_WLB<75> T_WLB<74> T_WLB<73> T_WLB<72> T_WLB<71> T_WLB<70> T_WLB<69> 
+ T_WLB<68> T_WLB<67> T_WLB<66> T_WLB<65> T_WLB<64> T_WLB<63> T_WLB<62> T_WLB<61> T_WLB<60> 
+ T_WLB<59> T_WLB<58> T_WLB<57> T_WLB<56> T_WLB<55> T_WLB<54> T_WLB<53> T_WLB<52> T_WLB<51> 
+ T_WLB<50> T_WLB<49> T_WLB<48> T_WLB<47> T_WLB<46> T_WLB<45> T_WLB<44> T_WLB<43> T_WLB<42> 
+ T_WLB<41> T_WLB<40> T_WLB<39> T_WLB<38> T_WLB<37> T_WLB<36> T_WLB<35> T_WLB<34> T_WLB<33> 
+ T_WLB<32> T_WLB<31> T_WLB<30> T_WLB<29> T_WLB<28> T_WLB<27> T_WLB<26> T_WLB<25> T_WLB<24> 
+ T_WLB<23> T_WLB<22> T_WLB<21> T_WLB<20> T_WLB<19> T_WLB<18> T_WLB<17> T_WLB<16> T_WLB<15> 
+ T_WLB<14> T_WLB<13> T_WLB<12> T_WLB<11> T_WLB<10> T_WLB<9> T_WLB<8> T_WLB<7> T_WLB<6> 
+ T_WLB<5> T_WLB<4> T_WLB<3> T_WLB<2> T_WLB<1> T_WLB<0> VDD VSS 
XCOL
+ B_DBL DWL<1> B_TIE_LOW DBL_PD_N<3> DBL_PD_N<2> DBL_PD_N<1> DBL_PD_N<0> STCLK T_DBL 
+ DWL<0> T_TIE_LOW VDD VSS  / xmc55_dps_localc8io_dummy
XAR_TOP
+ VSS T_DBL VSS T_TIE_LOW T_WLB<255> T_WLB<254> T_WLB<253> T_WLB<252> T_WLB<251> 
+ T_WLB<250> T_WLB<249> T_WLB<248> T_WLB<247> T_WLB<246> T_WLB<245> T_WLB<244> T_WLB<243> T_WLB<242> 
+ T_WLB<241> T_WLB<240> T_WLB<239> T_WLB<238> T_WLB<237> T_WLB<236> T_WLB<235> T_WLB<234> T_WLB<233> 
+ T_WLB<232> T_WLB<231> T_WLB<230> T_WLB<229> T_WLB<228> T_WLB<227> T_WLB<226> T_WLB<225> T_WLB<224> 
+ T_WLB<223> T_WLB<222> T_WLB<221> T_WLB<220> T_WLB<219> T_WLB<218> T_WLB<217> T_WLB<216> T_WLB<215> 
+ T_WLB<214> T_WLB<213> T_WLB<212> T_WLB<211> T_WLB<210> T_WLB<209> T_WLB<208> T_WLB<207> T_WLB<206> 
+ T_WLB<205> T_WLB<204> T_WLB<203> T_WLB<202> T_WLB<201> T_WLB<200> T_WLB<199> T_WLB<198> T_WLB<197> 
+ T_WLB<196> T_WLB<195> T_WLB<194> T_WLB<193> T_WLB<192> T_WLB<191> T_WLB<190> T_WLB<189> T_WLB<188> 
+ T_WLB<187> T_WLB<186> T_WLB<185> T_WLB<184> T_WLB<183> T_WLB<182> T_WLB<181> T_WLB<180> T_WLB<179> 
+ T_WLB<178> T_WLB<177> T_WLB<176> T_WLB<175> T_WLB<174> T_WLB<173> T_WLB<172> T_WLB<171> T_WLB<170> 
+ T_WLB<169> T_WLB<168> T_WLB<167> T_WLB<166> T_WLB<165> T_WLB<164> T_WLB<163> T_WLB<162> T_WLB<161> 
+ T_WLB<160> T_WLB<159> T_WLB<158> T_WLB<157> T_WLB<156> T_WLB<155> T_WLB<154> T_WLB<153> T_WLB<152> 
+ T_WLB<151> T_WLB<150> T_WLB<149> T_WLB<148> T_WLB<147> T_WLB<146> T_WLB<145> T_WLB<144> T_WLB<143> 
+ T_WLB<142> T_WLB<141> T_WLB<140> T_WLB<139> T_WLB<138> T_WLB<137> T_WLB<136> T_WLB<135> T_WLB<134> 
+ T_WLB<133> T_WLB<132> T_WLB<131> T_WLB<130> T_WLB<129> T_WLB<128> T_WLB<127> T_WLB<126> T_WLB<125> 
+ T_WLB<124> T_WLB<123> T_WLB<122> T_WLB<121> T_WLB<120> T_WLB<119> T_WLB<118> T_WLB<117> T_WLB<116> 
+ T_WLB<115> T_WLB<114> T_WLB<113> T_WLB<112> T_WLB<111> T_WLB<110> T_WLB<109> T_WLB<108> T_WLB<107> 
+ T_WLB<106> T_WLB<105> T_WLB<104> T_WLB<103> T_WLB<102> T_WLB<101> T_WLB<100> T_WLB<99> T_WLB<98> 
+ T_WLB<97> T_WLB<96> T_WLB<95> T_WLB<94> T_WLB<93> T_WLB<92> T_WLB<91> T_WLB<90> T_WLB<89> 
+ T_WLB<88> T_WLB<87> T_WLB<86> T_WLB<85> T_WLB<84> T_WLB<83> T_WLB<82> T_WLB<81> T_WLB<80> 
+ T_WLB<79> T_WLB<78> T_WLB<77> T_WLB<76> T_WLB<75> T_WLB<74> T_WLB<73> T_WLB<72> T_WLB<71> 
+ T_WLB<70> T_WLB<69> T_WLB<68> T_WLB<67> T_WLB<66> T_WLB<65> T_WLB<64> T_WLB<63> T_WLB<62> 
+ T_WLB<61> T_WLB<60> T_WLB<59> T_WLB<58> T_WLB<57> T_WLB<56> T_WLB<55> T_WLB<54> T_WLB<53> 
+ T_WLB<52> T_WLB<51> T_WLB<50> T_WLB<49> T_WLB<48> T_WLB<47> T_WLB<46> T_WLB<45> T_WLB<44> 
+ T_WLB<43> T_WLB<42> T_WLB<41> T_WLB<40> T_WLB<39> T_WLB<38> T_WLB<37> T_WLB<36> T_WLB<35> 
+ T_WLB<34> T_WLB<33> T_WLB<32> T_WLB<31> T_WLB<30> T_WLB<29> T_WLB<28> T_WLB<27> T_WLB<26> 
+ T_WLB<25> T_WLB<24> T_WLB<23> T_WLB<22> T_WLB<21> T_WLB<20> T_WLB<19> T_WLB<18> T_WLB<17> 
+ T_WLB<16> T_WLB<15> T_WLB<14> T_WLB<13> T_WLB<12> T_WLB<11> T_WLB<10> T_WLB<9> T_WLB<8> 
+ T_WLB<7> T_WLB<6> T_WLB<5> T_WLB<4> T_WLB<3> T_WLB<2> T_WLB<1> T_WLB<0>  / dpram16x4096_AR_DUMMY_ROWX256
XAR_BOT
+ VSS B_DBL VSS B_TIE_LOW B_WLB<255> B_WLB<254> B_WLB<253> B_WLB<252> B_WLB<251> 
+ B_WLB<250> B_WLB<249> B_WLB<248> B_WLB<247> B_WLB<246> B_WLB<245> B_WLB<244> B_WLB<243> B_WLB<242> 
+ B_WLB<241> B_WLB<240> B_WLB<239> B_WLB<238> B_WLB<237> B_WLB<236> B_WLB<235> B_WLB<234> B_WLB<233> 
+ B_WLB<232> B_WLB<231> B_WLB<230> B_WLB<229> B_WLB<228> B_WLB<227> B_WLB<226> B_WLB<225> B_WLB<224> 
+ B_WLB<223> B_WLB<222> B_WLB<221> B_WLB<220> B_WLB<219> B_WLB<218> B_WLB<217> B_WLB<216> B_WLB<215> 
+ B_WLB<214> B_WLB<213> B_WLB<212> B_WLB<211> B_WLB<210> B_WLB<209> B_WLB<208> B_WLB<207> B_WLB<206> 
+ B_WLB<205> B_WLB<204> B_WLB<203> B_WLB<202> B_WLB<201> B_WLB<200> B_WLB<199> B_WLB<198> B_WLB<197> 
+ B_WLB<196> B_WLB<195> B_WLB<194> B_WLB<193> B_WLB<192> B_WLB<191> B_WLB<190> B_WLB<189> B_WLB<188> 
+ B_WLB<187> B_WLB<186> B_WLB<185> B_WLB<184> B_WLB<183> B_WLB<182> B_WLB<181> B_WLB<180> B_WLB<179> 
+ B_WLB<178> B_WLB<177> B_WLB<176> B_WLB<175> B_WLB<174> B_WLB<173> B_WLB<172> B_WLB<171> B_WLB<170> 
+ B_WLB<169> B_WLB<168> B_WLB<167> B_WLB<166> B_WLB<165> B_WLB<164> B_WLB<163> B_WLB<162> B_WLB<161> 
+ B_WLB<160> B_WLB<159> B_WLB<158> B_WLB<157> B_WLB<156> B_WLB<155> B_WLB<154> B_WLB<153> B_WLB<152> 
+ B_WLB<151> B_WLB<150> B_WLB<149> B_WLB<148> B_WLB<147> B_WLB<146> B_WLB<145> B_WLB<144> B_WLB<143> 
+ B_WLB<142> B_WLB<141> B_WLB<140> B_WLB<139> B_WLB<138> B_WLB<137> B_WLB<136> B_WLB<135> B_WLB<134> 
+ B_WLB<133> B_WLB<132> B_WLB<131> B_WLB<130> B_WLB<129> B_WLB<128> B_WLB<127> B_WLB<126> B_WLB<125> 
+ B_WLB<124> B_WLB<123> B_WLB<122> B_WLB<121> B_WLB<120> B_WLB<119> B_WLB<118> B_WLB<117> B_WLB<116> 
+ B_WLB<115> B_WLB<114> B_WLB<113> B_WLB<112> B_WLB<111> B_WLB<110> B_WLB<109> B_WLB<108> B_WLB<107> 
+ B_WLB<106> B_WLB<105> B_WLB<104> B_WLB<103> B_WLB<102> B_WLB<101> B_WLB<100> B_WLB<99> B_WLB<98> 
+ B_WLB<97> B_WLB<96> B_WLB<95> B_WLB<94> B_WLB<93> B_WLB<92> B_WLB<91> B_WLB<90> B_WLB<89> 
+ B_WLB<88> B_WLB<87> B_WLB<86> B_WLB<85> B_WLB<84> B_WLB<83> B_WLB<82> B_WLB<81> B_WLB<80> 
+ B_WLB<79> B_WLB<78> B_WLB<77> B_WLB<76> B_WLB<75> B_WLB<74> B_WLB<73> B_WLB<72> B_WLB<71> 
+ B_WLB<70> B_WLB<69> B_WLB<68> B_WLB<67> B_WLB<66> B_WLB<65> B_WLB<64> B_WLB<63> B_WLB<62> 
+ B_WLB<61> B_WLB<60> B_WLB<59> B_WLB<58> B_WLB<57> B_WLB<56> B_WLB<55> B_WLB<54> B_WLB<53> 
+ B_WLB<52> B_WLB<51> B_WLB<50> B_WLB<49> B_WLB<48> B_WLB<47> B_WLB<46> B_WLB<45> B_WLB<44> 
+ B_WLB<43> B_WLB<42> B_WLB<41> B_WLB<40> B_WLB<39> B_WLB<38> B_WLB<37> B_WLB<36> B_WLB<35> 
+ B_WLB<34> B_WLB<33> B_WLB<32> B_WLB<31> B_WLB<30> B_WLB<29> B_WLB<28> B_WLB<27> B_WLB<26> 
+ B_WLB<25> B_WLB<24> B_WLB<23> B_WLB<22> B_WLB<21> B_WLB<20> B_WLB<19> B_WLB<18> B_WLB<17> 
+ B_WLB<16> B_WLB<15> B_WLB<14> B_WLB<13> B_WLB<12> B_WLB<11> B_WLB<10> B_WLB<9> B_WLB<8> 
+ B_WLB<7> B_WLB<6> B_WLB<5> B_WLB<4> B_WLB<3> B_WLB<2> B_WLB<1> B_WLB<0>  / dpram16x4096_AR_DUMMY_ROWX256
.ENDS

************************************************************************
* Cell Name:    dpram16x4096_AR_COLX8_ROWX256
* View Name:    schematic
************************************************************************
.SUBCKT dpram16x4096_AR_COLX8_ROWX256
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<255> WLA<254> WLA<253> WLA<252> WLA<251> WLA<250> WLA<249> WLA<248> 
+ WLA<247> WLA<246> WLA<245> WLA<244> WLA<243> WLA<242> WLA<241> WLA<240> WLA<239> 
+ WLA<238> WLA<237> WLA<236> WLA<235> WLA<234> WLA<233> WLA<232> WLA<231> WLA<230> 
+ WLA<229> WLA<228> WLA<227> WLA<226> WLA<225> WLA<224> WLA<223> WLA<222> WLA<221> 
+ WLA<220> WLA<219> WLA<218> WLA<217> WLA<216> WLA<215> WLA<214> WLA<213> WLA<212> 
+ WLA<211> WLA<210> WLA<209> WLA<208> WLA<207> WLA<206> WLA<205> WLA<204> WLA<203> 
+ WLA<202> WLA<201> WLA<200> WLA<199> WLA<198> WLA<197> WLA<196> WLA<195> WLA<194> 
+ WLA<193> WLA<192> WLA<191> WLA<190> WLA<189> WLA<188> WLA<187> WLA<186> WLA<185> 
+ WLA<184> WLA<183> WLA<182> WLA<181> WLA<180> WLA<179> WLA<178> WLA<177> WLA<176> 
+ WLA<175> WLA<174> WLA<173> WLA<172> WLA<171> WLA<170> WLA<169> WLA<168> WLA<167> 
+ WLA<166> WLA<165> WLA<164> WLA<163> WLA<162> WLA<161> WLA<160> WLA<159> WLA<158> 
+ WLA<157> WLA<156> WLA<155> WLA<154> WLA<153> WLA<152> WLA<151> WLA<150> WLA<149> 
+ WLA<148> WLA<147> WLA<146> WLA<145> WLA<144> WLA<143> WLA<142> WLA<141> WLA<140> 
+ WLA<139> WLA<138> WLA<137> WLA<136> WLA<135> WLA<134> WLA<133> WLA<132> WLA<131> 
+ WLA<130> WLA<129> WLA<128> WLA<127> WLA<126> WLA<125> WLA<124> WLA<123> WLA<122> 
+ WLA<121> WLA<120> WLA<119> WLA<118> WLA<117> WLA<116> WLA<115> WLA<114> WLA<113> 
+ WLA<112> WLA<111> WLA<110> WLA<109> WLA<108> WLA<107> WLA<106> WLA<105> WLA<104> 
+ WLA<103> WLA<102> WLA<101> WLA<100> WLA<99> WLA<98> WLA<97> WLA<96> WLA<95> 
+ WLA<94> WLA<93> WLA<92> WLA<91> WLA<90> WLA<89> WLA<88> WLA<87> WLA<86> 
+ WLA<85> WLA<84> WLA<83> WLA<82> WLA<81> WLA<80> WLA<79> WLA<78> WLA<77> 
+ WLA<76> WLA<75> WLA<74> WLA<73> WLA<72> WLA<71> WLA<70> WLA<69> WLA<68> 
+ WLA<67> WLA<66> WLA<65> WLA<64> WLA<63> WLA<62> WLA<61> WLA<60> WLA<59> 
+ WLA<58> WLA<57> WLA<56> WLA<55> WLA<54> WLA<53> WLA<52> WLA<51> WLA<50> 
+ WLA<49> WLA<48> WLA<47> WLA<46> WLA<45> WLA<44> WLA<43> WLA<42> WLA<41> 
+ WLA<40> WLA<39> WLA<38> WLA<37> WLA<36> WLA<35> WLA<34> WLA<33> WLA<32> 
+ WLA<31> WLA<30> WLA<29> WLA<28> WLA<27> WLA<26> WLA<25> WLA<24> WLA<23> 
+ WLA<22> WLA<21> WLA<20> WLA<19> WLA<18> WLA<17> WLA<16> WLA<15> WLA<14> 
+ WLA<13> WLA<12> WLA<11> WLA<10> WLA<9> WLA<8> WLA<7> WLA<6> WLA<5> 
+ WLA<4> WLA<3> WLA<2> WLA<1> WLA<0> WLB<255> WLB<254> WLB<253> WLB<252> 
+ WLB<251> WLB<250> WLB<249> WLB<248> WLB<247> WLB<246> WLB<245> WLB<244> WLB<243> 
+ WLB<242> WLB<241> WLB<240> WLB<239> WLB<238> WLB<237> WLB<236> WLB<235> WLB<234> 
+ WLB<233> WLB<232> WLB<231> WLB<230> WLB<229> WLB<228> WLB<227> WLB<226> WLB<225> 
+ WLB<224> WLB<223> WLB<222> WLB<221> WLB<220> WLB<219> WLB<218> WLB<217> WLB<216> 
+ WLB<215> WLB<214> WLB<213> WLB<212> WLB<211> WLB<210> WLB<209> WLB<208> WLB<207> 
+ WLB<206> WLB<205> WLB<204> WLB<203> WLB<202> WLB<201> WLB<200> WLB<199> WLB<198> 
+ WLB<197> WLB<196> WLB<195> WLB<194> WLB<193> WLB<192> WLB<191> WLB<190> WLB<189> 
+ WLB<188> WLB<187> WLB<186> WLB<185> WLB<184> WLB<183> WLB<182> WLB<181> WLB<180> 
+ WLB<179> WLB<178> WLB<177> WLB<176> WLB<175> WLB<174> WLB<173> WLB<172> WLB<171> 
+ WLB<170> WLB<169> WLB<168> WLB<167> WLB<166> WLB<165> WLB<164> WLB<163> WLB<162> 
+ WLB<161> WLB<160> WLB<159> WLB<158> WLB<157> WLB<156> WLB<155> WLB<154> WLB<153> 
+ WLB<152> WLB<151> WLB<150> WLB<149> WLB<148> WLB<147> WLB<146> WLB<145> WLB<144> 
+ WLB<143> WLB<142> WLB<141> WLB<140> WLB<139> WLB<138> WLB<137> WLB<136> WLB<135> 
+ WLB<134> WLB<133> WLB<132> WLB<131> WLB<130> WLB<129> WLB<128> WLB<127> WLB<126> 
+ WLB<125> WLB<124> WLB<123> WLB<122> WLB<121> WLB<120> WLB<119> WLB<118> WLB<117> 
+ WLB<116> WLB<115> WLB<114> WLB<113> WLB<112> WLB<111> WLB<110> WLB<109> WLB<108> 
+ WLB<107> WLB<106> WLB<105> WLB<104> WLB<103> WLB<102> WLB<101> WLB<100> WLB<99> 
+ WLB<98> WLB<97> WLB<96> WLB<95> WLB<94> WLB<93> WLB<92> WLB<91> WLB<90> 
+ WLB<89> WLB<88> WLB<87> WLB<86> WLB<85> WLB<84> WLB<83> WLB<82> WLB<81> 
+ WLB<80> WLB<79> WLB<78> WLB<77> WLB<76> WLB<75> WLB<74> WLB<73> WLB<72> 
+ WLB<71> WLB<70> WLB<69> WLB<68> WLB<67> WLB<66> WLB<65> WLB<64> WLB<63> 
+ WLB<62> WLB<61> WLB<60> WLB<59> WLB<58> WLB<57> WLB<56> WLB<55> WLB<54> 
+ WLB<53> WLB<52> WLB<51> WLB<50> WLB<49> WLB<48> WLB<47> WLB<46> WLB<45> 
+ WLB<44> WLB<43> WLB<42> WLB<41> WLB<40> WLB<39> WLB<38> WLB<37> WLB<36> 
+ WLB<35> WLB<34> WLB<33> WLB<32> WLB<31> WLB<30> WLB<29> WLB<28> WLB<27> 
+ WLB<26> WLB<25> WLB<24> WLB<23> WLB<22> WLB<21> WLB<20> WLB<19> WLB<18> 
+ WLB<17> WLB<16> WLB<15> WLB<14> WLB<13> WLB<12> WLB<11> WLB<10> WLB<9> 
+ WLB<8> WLB<7> WLB<6> WLB<5> WLB<4> WLB<3> WLB<2> WLB<1> WLB<0> 
+ 
XBITCELLS<127>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<255> WLA<254> WLB<255> WLB<254>  / CH974LP_bitcell_2x2
XBITCELLS<126>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<253> WLA<252> WLB<253> WLB<252>  / CH974LP_bitcell_2x2
XBITCELLS<125>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<251> WLA<250> WLB<251> WLB<250>  / CH974LP_bitcell_2x2
XBITCELLS<124>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<249> WLA<248> WLB<249> WLB<248>  / CH974LP_bitcell_2x2
XBITCELLS<123>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<247> WLA<246> WLB<247> WLB<246>  / CH974LP_bitcell_2x2
XBITCELLS<122>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<245> WLA<244> WLB<245> WLB<244>  / CH974LP_bitcell_2x2
XBITCELLS<121>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<243> WLA<242> WLB<243> WLB<242>  / CH974LP_bitcell_2x2
XBITCELLS<120>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<241> WLA<240> WLB<241> WLB<240>  / CH974LP_bitcell_2x2
XBITCELLS<119>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<239> WLA<238> WLB<239> WLB<238>  / CH974LP_bitcell_2x2
XBITCELLS<118>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<237> WLA<236> WLB<237> WLB<236>  / CH974LP_bitcell_2x2
XBITCELLS<117>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<235> WLA<234> WLB<235> WLB<234>  / CH974LP_bitcell_2x2
XBITCELLS<116>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<233> WLA<232> WLB<233> WLB<232>  / CH974LP_bitcell_2x2
XBITCELLS<115>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<231> WLA<230> WLB<231> WLB<230>  / CH974LP_bitcell_2x2
XBITCELLS<114>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<229> WLA<228> WLB<229> WLB<228>  / CH974LP_bitcell_2x2
XBITCELLS<113>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<227> WLA<226> WLB<227> WLB<226>  / CH974LP_bitcell_2x2
XBITCELLS<112>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<225> WLA<224> WLB<225> WLB<224>  / CH974LP_bitcell_2x2
XBITCELLS<111>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<223> WLA<222> WLB<223> WLB<222>  / CH974LP_bitcell_2x2
XBITCELLS<110>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<221> WLA<220> WLB<221> WLB<220>  / CH974LP_bitcell_2x2
XBITCELLS<109>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<219> WLA<218> WLB<219> WLB<218>  / CH974LP_bitcell_2x2
XBITCELLS<108>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<217> WLA<216> WLB<217> WLB<216>  / CH974LP_bitcell_2x2
XBITCELLS<107>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<215> WLA<214> WLB<215> WLB<214>  / CH974LP_bitcell_2x2
XBITCELLS<106>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<213> WLA<212> WLB<213> WLB<212>  / CH974LP_bitcell_2x2
XBITCELLS<105>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<211> WLA<210> WLB<211> WLB<210>  / CH974LP_bitcell_2x2
XBITCELLS<104>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<209> WLA<208> WLB<209> WLB<208>  / CH974LP_bitcell_2x2
XBITCELLS<103>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<207> WLA<206> WLB<207> WLB<206>  / CH974LP_bitcell_2x2
XBITCELLS<102>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<205> WLA<204> WLB<205> WLB<204>  / CH974LP_bitcell_2x2
XBITCELLS<101>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<203> WLA<202> WLB<203> WLB<202>  / CH974LP_bitcell_2x2
XBITCELLS<100>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<201> WLA<200> WLB<201> WLB<200>  / CH974LP_bitcell_2x2
XBITCELLS<99>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<199> WLA<198> WLB<199> WLB<198>  / CH974LP_bitcell_2x2
XBITCELLS<98>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<197> WLA<196> WLB<197> WLB<196>  / CH974LP_bitcell_2x2
XBITCELLS<97>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<195> WLA<194> WLB<195> WLB<194>  / CH974LP_bitcell_2x2
XBITCELLS<96>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<193> WLA<192> WLB<193> WLB<192>  / CH974LP_bitcell_2x2
XBITCELLS<95>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<191> WLA<190> WLB<191> WLB<190>  / CH974LP_bitcell_2x2
XBITCELLS<94>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<189> WLA<188> WLB<189> WLB<188>  / CH974LP_bitcell_2x2
XBITCELLS<93>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<187> WLA<186> WLB<187> WLB<186>  / CH974LP_bitcell_2x2
XBITCELLS<92>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<185> WLA<184> WLB<185> WLB<184>  / CH974LP_bitcell_2x2
XBITCELLS<91>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<183> WLA<182> WLB<183> WLB<182>  / CH974LP_bitcell_2x2
XBITCELLS<90>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<181> WLA<180> WLB<181> WLB<180>  / CH974LP_bitcell_2x2
XBITCELLS<89>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<179> WLA<178> WLB<179> WLB<178>  / CH974LP_bitcell_2x2
XBITCELLS<88>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<177> WLA<176> WLB<177> WLB<176>  / CH974LP_bitcell_2x2
XBITCELLS<87>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<175> WLA<174> WLB<175> WLB<174>  / CH974LP_bitcell_2x2
XBITCELLS<86>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<173> WLA<172> WLB<173> WLB<172>  / CH974LP_bitcell_2x2
XBITCELLS<85>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<171> WLA<170> WLB<171> WLB<170>  / CH974LP_bitcell_2x2
XBITCELLS<84>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<169> WLA<168> WLB<169> WLB<168>  / CH974LP_bitcell_2x2
XBITCELLS<83>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<167> WLA<166> WLB<167> WLB<166>  / CH974LP_bitcell_2x2
XBITCELLS<82>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<165> WLA<164> WLB<165> WLB<164>  / CH974LP_bitcell_2x2
XBITCELLS<81>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<163> WLA<162> WLB<163> WLB<162>  / CH974LP_bitcell_2x2
XBITCELLS<80>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<161> WLA<160> WLB<161> WLB<160>  / CH974LP_bitcell_2x2
XBITCELLS<79>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<159> WLA<158> WLB<159> WLB<158>  / CH974LP_bitcell_2x2
XBITCELLS<78>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<157> WLA<156> WLB<157> WLB<156>  / CH974LP_bitcell_2x2
XBITCELLS<77>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<155> WLA<154> WLB<155> WLB<154>  / CH974LP_bitcell_2x2
XBITCELLS<76>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<153> WLA<152> WLB<153> WLB<152>  / CH974LP_bitcell_2x2
XBITCELLS<75>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<151> WLA<150> WLB<151> WLB<150>  / CH974LP_bitcell_2x2
XBITCELLS<74>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<149> WLA<148> WLB<149> WLB<148>  / CH974LP_bitcell_2x2
XBITCELLS<73>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<147> WLA<146> WLB<147> WLB<146>  / CH974LP_bitcell_2x2
XBITCELLS<72>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<145> WLA<144> WLB<145> WLB<144>  / CH974LP_bitcell_2x2
XBITCELLS<71>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<143> WLA<142> WLB<143> WLB<142>  / CH974LP_bitcell_2x2
XBITCELLS<70>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<141> WLA<140> WLB<141> WLB<140>  / CH974LP_bitcell_2x2
XBITCELLS<69>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<139> WLA<138> WLB<139> WLB<138>  / CH974LP_bitcell_2x2
XBITCELLS<68>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<137> WLA<136> WLB<137> WLB<136>  / CH974LP_bitcell_2x2
XBITCELLS<67>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<135> WLA<134> WLB<135> WLB<134>  / CH974LP_bitcell_2x2
XBITCELLS<66>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<133> WLA<132> WLB<133> WLB<132>  / CH974LP_bitcell_2x2
XBITCELLS<65>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<131> WLA<130> WLB<131> WLB<130>  / CH974LP_bitcell_2x2
XBITCELLS<64>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<129> WLA<128> WLB<129> WLB<128>  / CH974LP_bitcell_2x2
XBITCELLS<63>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<127> WLA<126> WLB<127> WLB<126>  / CH974LP_bitcell_2x2
XBITCELLS<62>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<125> WLA<124> WLB<125> WLB<124>  / CH974LP_bitcell_2x2
XBITCELLS<61>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<123> WLA<122> WLB<123> WLB<122>  / CH974LP_bitcell_2x2
XBITCELLS<60>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<121> WLA<120> WLB<121> WLB<120>  / CH974LP_bitcell_2x2
XBITCELLS<59>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<119> WLA<118> WLB<119> WLB<118>  / CH974LP_bitcell_2x2
XBITCELLS<58>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<117> WLA<116> WLB<117> WLB<116>  / CH974LP_bitcell_2x2
XBITCELLS<57>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<115> WLA<114> WLB<115> WLB<114>  / CH974LP_bitcell_2x2
XBITCELLS<56>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<113> WLA<112> WLB<113> WLB<112>  / CH974LP_bitcell_2x2
XBITCELLS<55>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<111> WLA<110> WLB<111> WLB<110>  / CH974LP_bitcell_2x2
XBITCELLS<54>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<109> WLA<108> WLB<109> WLB<108>  / CH974LP_bitcell_2x2
XBITCELLS<53>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<107> WLA<106> WLB<107> WLB<106>  / CH974LP_bitcell_2x2
XBITCELLS<52>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<105> WLA<104> WLB<105> WLB<104>  / CH974LP_bitcell_2x2
XBITCELLS<51>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<103> WLA<102> WLB<103> WLB<102>  / CH974LP_bitcell_2x2
XBITCELLS<50>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<101> WLA<100> WLB<101> WLB<100>  / CH974LP_bitcell_2x2
XBITCELLS<49>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<99> WLA<98> WLB<99> WLB<98>  / CH974LP_bitcell_2x2
XBITCELLS<48>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<97> WLA<96> WLB<97> WLB<96>  / CH974LP_bitcell_2x2
XBITCELLS<47>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<95> WLA<94> WLB<95> WLB<94>  / CH974LP_bitcell_2x2
XBITCELLS<46>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<93> WLA<92> WLB<93> WLB<92>  / CH974LP_bitcell_2x2
XBITCELLS<45>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<91> WLA<90> WLB<91> WLB<90>  / CH974LP_bitcell_2x2
XBITCELLS<44>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<89> WLA<88> WLB<89> WLB<88>  / CH974LP_bitcell_2x2
XBITCELLS<43>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<87> WLA<86> WLB<87> WLB<86>  / CH974LP_bitcell_2x2
XBITCELLS<42>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<85> WLA<84> WLB<85> WLB<84>  / CH974LP_bitcell_2x2
XBITCELLS<41>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<83> WLA<82> WLB<83> WLB<82>  / CH974LP_bitcell_2x2
XBITCELLS<40>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<81> WLA<80> WLB<81> WLB<80>  / CH974LP_bitcell_2x2
XBITCELLS<39>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<79> WLA<78> WLB<79> WLB<78>  / CH974LP_bitcell_2x2
XBITCELLS<38>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<77> WLA<76> WLB<77> WLB<76>  / CH974LP_bitcell_2x2
XBITCELLS<37>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<75> WLA<74> WLB<75> WLB<74>  / CH974LP_bitcell_2x2
XBITCELLS<36>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<73> WLA<72> WLB<73> WLB<72>  / CH974LP_bitcell_2x2
XBITCELLS<35>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<71> WLA<70> WLB<71> WLB<70>  / CH974LP_bitcell_2x2
XBITCELLS<34>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<69> WLA<68> WLB<69> WLB<68>  / CH974LP_bitcell_2x2
XBITCELLS<33>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<67> WLA<66> WLB<67> WLB<66>  / CH974LP_bitcell_2x2
XBITCELLS<32>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<65> WLA<64> WLB<65> WLB<64>  / CH974LP_bitcell_2x2
XBITCELLS<31>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<63> WLA<62> WLB<63> WLB<62>  / CH974LP_bitcell_2x2
XBITCELLS<30>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<61> WLA<60> WLB<61> WLB<60>  / CH974LP_bitcell_2x2
XBITCELLS<29>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<59> WLA<58> WLB<59> WLB<58>  / CH974LP_bitcell_2x2
XBITCELLS<28>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<57> WLA<56> WLB<57> WLB<56>  / CH974LP_bitcell_2x2
XBITCELLS<27>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<55> WLA<54> WLB<55> WLB<54>  / CH974LP_bitcell_2x2
XBITCELLS<26>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<53> WLA<52> WLB<53> WLB<52>  / CH974LP_bitcell_2x2
XBITCELLS<25>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<51> WLA<50> WLB<51> WLB<50>  / CH974LP_bitcell_2x2
XBITCELLS<24>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<49> WLA<48> WLB<49> WLB<48>  / CH974LP_bitcell_2x2
XBITCELLS<23>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<47> WLA<46> WLB<47> WLB<46>  / CH974LP_bitcell_2x2
XBITCELLS<22>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<45> WLA<44> WLB<45> WLB<44>  / CH974LP_bitcell_2x2
XBITCELLS<21>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<43> WLA<42> WLB<43> WLB<42>  / CH974LP_bitcell_2x2
XBITCELLS<20>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<41> WLA<40> WLB<41> WLB<40>  / CH974LP_bitcell_2x2
XBITCELLS<19>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<39> WLA<38> WLB<39> WLB<38>  / CH974LP_bitcell_2x2
XBITCELLS<18>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<37> WLA<36> WLB<37> WLB<36>  / CH974LP_bitcell_2x2
XBITCELLS<17>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<35> WLA<34> WLB<35> WLB<34>  / CH974LP_bitcell_2x2
XBITCELLS<16>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<33> WLA<32> WLB<33> WLB<32>  / CH974LP_bitcell_2x2
XBITCELLS<15>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<31> WLA<30> WLB<31> WLB<30>  / CH974LP_bitcell_2x2
XBITCELLS<14>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<29> WLA<28> WLB<29> WLB<28>  / CH974LP_bitcell_2x2
XBITCELLS<13>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<27> WLA<26> WLB<27> WLB<26>  / CH974LP_bitcell_2x2
XBITCELLS<12>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<25> WLA<24> WLB<25> WLB<24>  / CH974LP_bitcell_2x2
XBITCELLS<11>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<23> WLA<22> WLB<23> WLB<22>  / CH974LP_bitcell_2x2
XBITCELLS<10>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<21> WLA<20> WLB<21> WLB<20>  / CH974LP_bitcell_2x2
XBITCELLS<9>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<19> WLA<18> WLB<19> WLB<18>  / CH974LP_bitcell_2x2
XBITCELLS<8>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<17> WLA<16> WLB<17> WLB<16>  / CH974LP_bitcell_2x2
XBITCELLS<7>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<15> WLA<14> WLB<15> WLB<14>  / CH974LP_bitcell_2x2
XBITCELLS<6>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<13> WLA<12> WLB<13> WLB<12>  / CH974LP_bitcell_2x2
XBITCELLS<5>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<11> WLA<10> WLB<11> WLB<10>  / CH974LP_bitcell_2x2
XBITCELLS<4>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<9> WLA<8> WLB<9> WLB<8>  / CH974LP_bitcell_2x2
XBITCELLS<3>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<7> WLA<6> WLB<7> WLB<6>  / CH974LP_bitcell_2x2
XBITCELLS<2>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<5> WLA<4> WLB<5> WLB<4>  / CH974LP_bitcell_2x2
XBITCELLS<1>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<3> WLA<2> WLB<3> WLB<2>  / CH974LP_bitcell_2x2
XBITCELLS<0>
+ BLA<1> BLA<0> BLA_N<1> BLA_N<0> BLB<1> BLB<0> BLB_N<1> BLB_N<0> GND 
+ VDD WLA<1> WLA<0> WLB<1> WLB<0>  / CH974LP_bitcell_2x2
.ENDS

************************************************************************
* Cell Name:    dpram16x4096_SingleCOL2X8_ROWX256
* View Name:    schematic
************************************************************************
.SUBCKT dpram16x4096_SingleCOL2X8_ROWX256
+ B_CA<3> B_CA<2> B_CA<1> B_CA<0> B_CB<3> B_CB<2> B_CB<1> B_CB<0> B_MA<3> 
+ B_MA<2> B_MA<1> B_MA<0> B_MB<3> B_MB<2> B_MB<1> B_MB<0> B_TM_PREA_N B_TM_PREB_N 
+ B_WLA<255> B_WLA<254> B_WLA<253> B_WLA<252> B_WLA<251> B_WLA<250> B_WLA<249> B_WLA<248> B_WLA<247> 
+ B_WLA<246> B_WLA<245> B_WLA<244> B_WLA<243> B_WLA<242> B_WLA<241> B_WLA<240> B_WLA<239> B_WLA<238> 
+ B_WLA<237> B_WLA<236> B_WLA<235> B_WLA<234> B_WLA<233> B_WLA<232> B_WLA<231> B_WLA<230> B_WLA<229> 
+ B_WLA<228> B_WLA<227> B_WLA<226> B_WLA<225> B_WLA<224> B_WLA<223> B_WLA<222> B_WLA<221> B_WLA<220> 
+ B_WLA<219> B_WLA<218> B_WLA<217> B_WLA<216> B_WLA<215> B_WLA<214> B_WLA<213> B_WLA<212> B_WLA<211> 
+ B_WLA<210> B_WLA<209> B_WLA<208> B_WLA<207> B_WLA<206> B_WLA<205> B_WLA<204> B_WLA<203> B_WLA<202> 
+ B_WLA<201> B_WLA<200> B_WLA<199> B_WLA<198> B_WLA<197> B_WLA<196> B_WLA<195> B_WLA<194> B_WLA<193> 
+ B_WLA<192> B_WLA<191> B_WLA<190> B_WLA<189> B_WLA<188> B_WLA<187> B_WLA<186> B_WLA<185> B_WLA<184> 
+ B_WLA<183> B_WLA<182> B_WLA<181> B_WLA<180> B_WLA<179> B_WLA<178> B_WLA<177> B_WLA<176> B_WLA<175> 
+ B_WLA<174> B_WLA<173> B_WLA<172> B_WLA<171> B_WLA<170> B_WLA<169> B_WLA<168> B_WLA<167> B_WLA<166> 
+ B_WLA<165> B_WLA<164> B_WLA<163> B_WLA<162> B_WLA<161> B_WLA<160> B_WLA<159> B_WLA<158> B_WLA<157> 
+ B_WLA<156> B_WLA<155> B_WLA<154> B_WLA<153> B_WLA<152> B_WLA<151> B_WLA<150> B_WLA<149> B_WLA<148> 
+ B_WLA<147> B_WLA<146> B_WLA<145> B_WLA<144> B_WLA<143> B_WLA<142> B_WLA<141> B_WLA<140> B_WLA<139> 
+ B_WLA<138> B_WLA<137> B_WLA<136> B_WLA<135> B_WLA<134> B_WLA<133> B_WLA<132> B_WLA<131> B_WLA<130> 
+ B_WLA<129> B_WLA<128> B_WLA<127> B_WLA<126> B_WLA<125> B_WLA<124> B_WLA<123> B_WLA<122> B_WLA<121> 
+ B_WLA<120> B_WLA<119> B_WLA<118> B_WLA<117> B_WLA<116> B_WLA<115> B_WLA<114> B_WLA<113> B_WLA<112> 
+ B_WLA<111> B_WLA<110> B_WLA<109> B_WLA<108> B_WLA<107> B_WLA<106> B_WLA<105> B_WLA<104> B_WLA<103> 
+ B_WLA<102> B_WLA<101> B_WLA<100> B_WLA<99> B_WLA<98> B_WLA<97> B_WLA<96> B_WLA<95> B_WLA<94> 
+ B_WLA<93> B_WLA<92> B_WLA<91> B_WLA<90> B_WLA<89> B_WLA<88> B_WLA<87> B_WLA<86> B_WLA<85> 
+ B_WLA<84> B_WLA<83> B_WLA<82> B_WLA<81> B_WLA<80> B_WLA<79> B_WLA<78> B_WLA<77> B_WLA<76> 
+ B_WLA<75> B_WLA<74> B_WLA<73> B_WLA<72> B_WLA<71> B_WLA<70> B_WLA<69> B_WLA<68> B_WLA<67> 
+ B_WLA<66> B_WLA<65> B_WLA<64> B_WLA<63> B_WLA<62> B_WLA<61> B_WLA<60> B_WLA<59> B_WLA<58> 
+ B_WLA<57> B_WLA<56> B_WLA<55> B_WLA<54> B_WLA<53> B_WLA<52> B_WLA<51> B_WLA<50> B_WLA<49> 
+ B_WLA<48> B_WLA<47> B_WLA<46> B_WLA<45> B_WLA<44> B_WLA<43> B_WLA<42> B_WLA<41> B_WLA<40> 
+ B_WLA<39> B_WLA<38> B_WLA<37> B_WLA<36> B_WLA<35> B_WLA<34> B_WLA<33> B_WLA<32> B_WLA<31> 
+ B_WLA<30> B_WLA<29> B_WLA<28> B_WLA<27> B_WLA<26> B_WLA<25> B_WLA<24> B_WLA<23> B_WLA<22> 
+ B_WLA<21> B_WLA<20> B_WLA<19> B_WLA<18> B_WLA<17> B_WLA<16> B_WLA<15> B_WLA<14> B_WLA<13> 
+ B_WLA<12> B_WLA<11> B_WLA<10> B_WLA<9> B_WLA<8> B_WLA<7> B_WLA<6> B_WLA<5> B_WLA<4> 
+ B_WLA<3> B_WLA<2> B_WLA<1> B_WLA<0> B_WLB<255> B_WLB<254> B_WLB<253> B_WLB<252> B_WLB<251> 
+ B_WLB<250> B_WLB<249> B_WLB<248> B_WLB<247> B_WLB<246> B_WLB<245> B_WLB<244> B_WLB<243> B_WLB<242> 
+ B_WLB<241> B_WLB<240> B_WLB<239> B_WLB<238> B_WLB<237> B_WLB<236> B_WLB<235> B_WLB<234> B_WLB<233> 
+ B_WLB<232> B_WLB<231> B_WLB<230> B_WLB<229> B_WLB<228> B_WLB<227> B_WLB<226> B_WLB<225> B_WLB<224> 
+ B_WLB<223> B_WLB<222> B_WLB<221> B_WLB<220> B_WLB<219> B_WLB<218> B_WLB<217> B_WLB<216> B_WLB<215> 
+ B_WLB<214> B_WLB<213> B_WLB<212> B_WLB<211> B_WLB<210> B_WLB<209> B_WLB<208> B_WLB<207> B_WLB<206> 
+ B_WLB<205> B_WLB<204> B_WLB<203> B_WLB<202> B_WLB<201> B_WLB<200> B_WLB<199> B_WLB<198> B_WLB<197> 
+ B_WLB<196> B_WLB<195> B_WLB<194> B_WLB<193> B_WLB<192> B_WLB<191> B_WLB<190> B_WLB<189> B_WLB<188> 
+ B_WLB<187> B_WLB<186> B_WLB<185> B_WLB<184> B_WLB<183> B_WLB<182> B_WLB<181> B_WLB<180> B_WLB<179> 
+ B_WLB<178> B_WLB<177> B_WLB<176> B_WLB<175> B_WLB<174> B_WLB<173> B_WLB<172> B_WLB<171> B_WLB<170> 
+ B_WLB<169> B_WLB<168> B_WLB<167> B_WLB<166> B_WLB<165> B_WLB<164> B_WLB<163> B_WLB<162> B_WLB<161> 
+ B_WLB<160> B_WLB<159> B_WLB<158> B_WLB<157> B_WLB<156> B_WLB<155> B_WLB<154> B_WLB<153> B_WLB<152> 
+ B_WLB<151> B_WLB<150> B_WLB<149> B_WLB<148> B_WLB<147> B_WLB<146> B_WLB<145> B_WLB<144> B_WLB<143> 
+ B_WLB<142> B_WLB<141> B_WLB<140> B_WLB<139> B_WLB<138> B_WLB<137> B_WLB<136> B_WLB<135> B_WLB<134> 
+ B_WLB<133> B_WLB<132> B_WLB<131> B_WLB<130> B_WLB<129> B_WLB<128> B_WLB<127> B_WLB<126> B_WLB<125> 
+ B_WLB<124> B_WLB<123> B_WLB<122> B_WLB<121> B_WLB<120> B_WLB<119> B_WLB<118> B_WLB<117> B_WLB<116> 
+ B_WLB<115> B_WLB<114> B_WLB<113> B_WLB<112> B_WLB<111> B_WLB<110> B_WLB<109> B_WLB<108> B_WLB<107> 
+ B_WLB<106> B_WLB<105> B_WLB<104> B_WLB<103> B_WLB<102> B_WLB<101> B_WLB<100> B_WLB<99> B_WLB<98> 
+ B_WLB<97> B_WLB<96> B_WLB<95> B_WLB<94> B_WLB<93> B_WLB<92> B_WLB<91> B_WLB<90> B_WLB<89> 
+ B_WLB<88> B_WLB<87> B_WLB<86> B_WLB<85> B_WLB<84> B_WLB<83> B_WLB<82> B_WLB<81> B_WLB<80> 
+ B_WLB<79> B_WLB<78> B_WLB<77> B_WLB<76> B_WLB<75> B_WLB<74> B_WLB<73> B_WLB<72> B_WLB<71> 
+ B_WLB<70> B_WLB<69> B_WLB<68> B_WLB<67> B_WLB<66> B_WLB<65> B_WLB<64> B_WLB<63> B_WLB<62> 
+ B_WLB<61> B_WLB<60> B_WLB<59> B_WLB<58> B_WLB<57> B_WLB<56> B_WLB<55> B_WLB<54> B_WLB<53> 
+ B_WLB<52> B_WLB<51> B_WLB<50> B_WLB<49> B_WLB<48> B_WLB<47> B_WLB<46> B_WLB<45> B_WLB<44> 
+ B_WLB<43> B_WLB<42> B_WLB<41> B_WLB<40> B_WLB<39> B_WLB<38> B_WLB<37> B_WLB<36> B_WLB<35> 
+ B_WLB<34> B_WLB<33> B_WLB<32> B_WLB<31> B_WLB<30> B_WLB<29> B_WLB<28> B_WLB<27> B_WLB<26> 
+ B_WLB<25> B_WLB<24> B_WLB<23> B_WLB<22> B_WLB<21> B_WLB<20> B_WLB<19> B_WLB<18> B_WLB<17> 
+ B_WLB<16> B_WLB<15> B_WLB<14> B_WLB<13> B_WLB<12> B_WLB<11> B_WLB<10> B_WLB<9> B_WLB<8> 
+ B_WLB<7> B_WLB<6> B_WLB<5> B_WLB<4> B_WLB<3> B_WLB<2> B_WLB<1> B_WLB<0> BWENA<1> 
+ BWENA<0> BWENB<1> BWENB<0> CLK_DQA CLK_DQA_N CLK_DQB CLK_DQB_N DA<1> DA<0> 
+ DB<1> DB<0> DDQA DDQA_N DDQB DDQB_N LWEA LWEB QA<1> 
+ QA<0> QB<1> QB<0> SA_PREA_N SA_PREB_N SAEA_N SAEB_N T_CA<3> T_CA<2> 
+ T_CA<1> T_CA<0> T_CB<3> T_CB<2> T_CB<1> T_CB<0> T_MA<3> T_MA<2> T_MA<1> 
+ T_MA<0> T_MB<3> T_MB<2> T_MB<1> T_MB<0> T_TM_PREA_N T_TM_PREB_N T_WLA<255> T_WLA<254> 
+ T_WLA<253> T_WLA<252> T_WLA<251> T_WLA<250> T_WLA<249> T_WLA<248> T_WLA<247> T_WLA<246> T_WLA<245> 
+ T_WLA<244> T_WLA<243> T_WLA<242> T_WLA<241> T_WLA<240> T_WLA<239> T_WLA<238> T_WLA<237> T_WLA<236> 
+ T_WLA<235> T_WLA<234> T_WLA<233> T_WLA<232> T_WLA<231> T_WLA<230> T_WLA<229> T_WLA<228> T_WLA<227> 
+ T_WLA<226> T_WLA<225> T_WLA<224> T_WLA<223> T_WLA<222> T_WLA<221> T_WLA<220> T_WLA<219> T_WLA<218> 
+ T_WLA<217> T_WLA<216> T_WLA<215> T_WLA<214> T_WLA<213> T_WLA<212> T_WLA<211> T_WLA<210> T_WLA<209> 
+ T_WLA<208> T_WLA<207> T_WLA<206> T_WLA<205> T_WLA<204> T_WLA<203> T_WLA<202> T_WLA<201> T_WLA<200> 
+ T_WLA<199> T_WLA<198> T_WLA<197> T_WLA<196> T_WLA<195> T_WLA<194> T_WLA<193> T_WLA<192> T_WLA<191> 
+ T_WLA<190> T_WLA<189> T_WLA<188> T_WLA<187> T_WLA<186> T_WLA<185> T_WLA<184> T_WLA<183> T_WLA<182> 
+ T_WLA<181> T_WLA<180> T_WLA<179> T_WLA<178> T_WLA<177> T_WLA<176> T_WLA<175> T_WLA<174> T_WLA<173> 
+ T_WLA<172> T_WLA<171> T_WLA<170> T_WLA<169> T_WLA<168> T_WLA<167> T_WLA<166> T_WLA<165> T_WLA<164> 
+ T_WLA<163> T_WLA<162> T_WLA<161> T_WLA<160> T_WLA<159> T_WLA<158> T_WLA<157> T_WLA<156> T_WLA<155> 
+ T_WLA<154> T_WLA<153> T_WLA<152> T_WLA<151> T_WLA<150> T_WLA<149> T_WLA<148> T_WLA<147> T_WLA<146> 
+ T_WLA<145> T_WLA<144> T_WLA<143> T_WLA<142> T_WLA<141> T_WLA<140> T_WLA<139> T_WLA<138> T_WLA<137> 
+ T_WLA<136> T_WLA<135> T_WLA<134> T_WLA<133> T_WLA<132> T_WLA<131> T_WLA<130> T_WLA<129> T_WLA<128> 
+ T_WLA<127> T_WLA<126> T_WLA<125> T_WLA<124> T_WLA<123> T_WLA<122> T_WLA<121> T_WLA<120> T_WLA<119> 
+ T_WLA<118> T_WLA<117> T_WLA<116> T_WLA<115> T_WLA<114> T_WLA<113> T_WLA<112> T_WLA<111> T_WLA<110> 
+ T_WLA<109> T_WLA<108> T_WLA<107> T_WLA<106> T_WLA<105> T_WLA<104> T_WLA<103> T_WLA<102> T_WLA<101> 
+ T_WLA<100> T_WLA<99> T_WLA<98> T_WLA<97> T_WLA<96> T_WLA<95> T_WLA<94> T_WLA<93> T_WLA<92> 
+ T_WLA<91> T_WLA<90> T_WLA<89> T_WLA<88> T_WLA<87> T_WLA<86> T_WLA<85> T_WLA<84> T_WLA<83> 
+ T_WLA<82> T_WLA<81> T_WLA<80> T_WLA<79> T_WLA<78> T_WLA<77> T_WLA<76> T_WLA<75> T_WLA<74> 
+ T_WLA<73> T_WLA<72> T_WLA<71> T_WLA<70> T_WLA<69> T_WLA<68> T_WLA<67> T_WLA<66> T_WLA<65> 
+ T_WLA<64> T_WLA<63> T_WLA<62> T_WLA<61> T_WLA<60> T_WLA<59> T_WLA<58> T_WLA<57> T_WLA<56> 
+ T_WLA<55> T_WLA<54> T_WLA<53> T_WLA<52> T_WLA<51> T_WLA<50> T_WLA<49> T_WLA<48> T_WLA<47> 
+ T_WLA<46> T_WLA<45> T_WLA<44> T_WLA<43> T_WLA<42> T_WLA<41> T_WLA<40> T_WLA<39> T_WLA<38> 
+ T_WLA<37> T_WLA<36> T_WLA<35> T_WLA<34> T_WLA<33> T_WLA<32> T_WLA<31> T_WLA<30> T_WLA<29> 
+ T_WLA<28> T_WLA<27> T_WLA<26> T_WLA<25> T_WLA<24> T_WLA<23> T_WLA<22> T_WLA<21> T_WLA<20> 
+ T_WLA<19> T_WLA<18> T_WLA<17> T_WLA<16> T_WLA<15> T_WLA<14> T_WLA<13> T_WLA<12> T_WLA<11> 
+ T_WLA<10> T_WLA<9> T_WLA<8> T_WLA<7> T_WLA<6> T_WLA<5> T_WLA<4> T_WLA<3> T_WLA<2> 
+ T_WLA<1> T_WLA<0> T_WLB<255> T_WLB<254> T_WLB<253> T_WLB<252> T_WLB<251> T_WLB<250> T_WLB<249> 
+ T_WLB<248> T_WLB<247> T_WLB<246> T_WLB<245> T_WLB<244> T_WLB<243> T_WLB<242> T_WLB<241> T_WLB<240> 
+ T_WLB<239> T_WLB<238> T_WLB<237> T_WLB<236> T_WLB<235> T_WLB<234> T_WLB<233> T_WLB<232> T_WLB<231> 
+ T_WLB<230> T_WLB<229> T_WLB<228> T_WLB<227> T_WLB<226> T_WLB<225> T_WLB<224> T_WLB<223> T_WLB<222> 
+ T_WLB<221> T_WLB<220> T_WLB<219> T_WLB<218> T_WLB<217> T_WLB<216> T_WLB<215> T_WLB<214> T_WLB<213> 
+ T_WLB<212> T_WLB<211> T_WLB<210> T_WLB<209> T_WLB<208> T_WLB<207> T_WLB<206> T_WLB<205> T_WLB<204> 
+ T_WLB<203> T_WLB<202> T_WLB<201> T_WLB<200> T_WLB<199> T_WLB<198> T_WLB<197> T_WLB<196> T_WLB<195> 
+ T_WLB<194> T_WLB<193> T_WLB<192> T_WLB<191> T_WLB<190> T_WLB<189> T_WLB<188> T_WLB<187> T_WLB<186> 
+ T_WLB<185> T_WLB<184> T_WLB<183> T_WLB<182> T_WLB<181> T_WLB<180> T_WLB<179> T_WLB<178> T_WLB<177> 
+ T_WLB<176> T_WLB<175> T_WLB<174> T_WLB<173> T_WLB<172> T_WLB<171> T_WLB<170> T_WLB<169> T_WLB<168> 
+ T_WLB<167> T_WLB<166> T_WLB<165> T_WLB<164> T_WLB<163> T_WLB<162> T_WLB<161> T_WLB<160> T_WLB<159> 
+ T_WLB<158> T_WLB<157> T_WLB<156> T_WLB<155> T_WLB<154> T_WLB<153> T_WLB<152> T_WLB<151> T_WLB<150> 
+ T_WLB<149> T_WLB<148> T_WLB<147> T_WLB<146> T_WLB<145> T_WLB<144> T_WLB<143> T_WLB<142> T_WLB<141> 
+ T_WLB<140> T_WLB<139> T_WLB<138> T_WLB<137> T_WLB<136> T_WLB<135> T_WLB<134> T_WLB<133> T_WLB<132> 
+ T_WLB<131> T_WLB<130> T_WLB<129> T_WLB<128> T_WLB<127> T_WLB<126> T_WLB<125> T_WLB<124> T_WLB<123> 
+ T_WLB<122> T_WLB<121> T_WLB<120> T_WLB<119> T_WLB<118> T_WLB<117> T_WLB<116> T_WLB<115> T_WLB<114> 
+ T_WLB<113> T_WLB<112> T_WLB<111> T_WLB<110> T_WLB<109> T_WLB<108> T_WLB<107> T_WLB<106> T_WLB<105> 
+ T_WLB<104> T_WLB<103> T_WLB<102> T_WLB<101> T_WLB<100> T_WLB<99> T_WLB<98> T_WLB<97> T_WLB<96> 
+ T_WLB<95> T_WLB<94> T_WLB<93> T_WLB<92> T_WLB<91> T_WLB<90> T_WLB<89> T_WLB<88> T_WLB<87> 
+ T_WLB<86> T_WLB<85> T_WLB<84> T_WLB<83> T_WLB<82> T_WLB<81> T_WLB<80> T_WLB<79> T_WLB<78> 
+ T_WLB<77> T_WLB<76> T_WLB<75> T_WLB<74> T_WLB<73> T_WLB<72> T_WLB<71> T_WLB<70> T_WLB<69> 
+ T_WLB<68> T_WLB<67> T_WLB<66> T_WLB<65> T_WLB<64> T_WLB<63> T_WLB<62> T_WLB<61> T_WLB<60> 
+ T_WLB<59> T_WLB<58> T_WLB<57> T_WLB<56> T_WLB<55> T_WLB<54> T_WLB<53> T_WLB<52> T_WLB<51> 
+ T_WLB<50> T_WLB<49> T_WLB<48> T_WLB<47> T_WLB<46> T_WLB<45> T_WLB<44> T_WLB<43> T_WLB<42> 
+ T_WLB<41> T_WLB<40> T_WLB<39> T_WLB<38> T_WLB<37> T_WLB<36> T_WLB<35> T_WLB<34> T_WLB<33> 
+ T_WLB<32> T_WLB<31> T_WLB<30> T_WLB<29> T_WLB<28> T_WLB<27> T_WLB<26> T_WLB<25> T_WLB<24> 
+ T_WLB<23> T_WLB<22> T_WLB<21> T_WLB<20> T_WLB<19> T_WLB<18> T_WLB<17> T_WLB<16> T_WLB<15> 
+ T_WLB<14> T_WLB<13> T_WLB<12> T_WLB<11> T_WLB<10> T_WLB<9> T_WLB<8> T_WLB<7> T_WLB<6> 
+ T_WLB<5> T_WLB<4> T_WLB<3> T_WLB<2> T_WLB<1> T_WLB<0> VDD VSS 
XCOL0
+ B_BLA<7> B_BLA<6> B_BLA<5> B_BLA<4> B_BLA<3> B_BLA<2> B_BLA<1> B_BLA<0> B_BLA_N<7> 
+ B_BLA_N<6> B_BLA_N<5> B_BLA_N<4> B_BLA_N<3> B_BLA_N<2> B_BLA_N<1> B_BLA_N<0> B_BLB<7> B_BLB<6> 
+ B_BLB<5> B_BLB<4> B_BLB<3> B_BLB<2> B_BLB<1> B_BLB<0> B_BLB_N<7> B_BLB_N<6> B_BLB_N<5> 
+ B_BLB_N<4> B_BLB_N<3> B_BLB_N<2> B_BLB_N<1> B_BLB_N<0> B_CA<3> B_CA<2> B_CA<1> B_CA<0> 
+ B_CB<3> B_CB<2> B_CB<1> B_CB<0> B_MA<3> B_MA<2> B_MA<1> B_MA<0> B_MB<3> 
+ B_MB<2> B_MB<1> B_MB<0> B_TM_PREA_N B_TM_PREB_N BWENA_INT<0> BWENB_INT<0> CLK_DQA CLK_DQA_N 
+ CLK_DQB CLK_DQB_N DA_INT<0> DB_INT<0> DDQA DDQA_N DDQB DDQB_N LWEA 
+ LWEB QA_INT<0> QB_INT<0> SA_PREA_N SA_PREB_N SAEA_N SAEB_N T_BLA<7> T_BLA<6> 
+ T_BLA<5> T_BLA<4> T_BLA<3> T_BLA<2> T_BLA<1> T_BLA<0> T_BLA_N<7> T_BLA_N<6> T_BLA_N<5> 
+ T_BLA_N<4> T_BLA_N<3> T_BLA_N<2> T_BLA_N<1> T_BLA_N<0> T_BLB<7> T_BLB<6> T_BLB<5> T_BLB<4> 
+ T_BLB<3> T_BLB<2> T_BLB<1> T_BLB<0> T_BLB_N<7> T_BLB_N<6> T_BLB_N<5> T_BLB_N<4> T_BLB_N<3> 
+ T_BLB_N<2> T_BLB_N<1> T_BLB_N<0> T_CA<3> T_CA<2> T_CA<1> T_CA<0> T_CB<3> T_CB<2> 
+ T_CB<1> T_CB<0> T_MA<3> T_MA<2> T_MA<1> T_MA<0> T_MB<3> T_MB<2> T_MB<1> 
+ T_MB<0> T_TM_PREA_N T_TM_PREB_N VDD VSS  / xmc55_dps_localc8io_bw
XCOL1
+ B_BLA<15> B_BLA<14> B_BLA<13> B_BLA<12> B_BLA<11> B_BLA<10> B_BLA<9> B_BLA<8> B_BLA_N<15> 
+ B_BLA_N<14> B_BLA_N<13> B_BLA_N<12> B_BLA_N<11> B_BLA_N<10> B_BLA_N<9> B_BLA_N<8> B_BLB<15> B_BLB<14> 
+ B_BLB<13> B_BLB<12> B_BLB<11> B_BLB<10> B_BLB<9> B_BLB<8> B_BLB_N<15> B_BLB_N<14> B_BLB_N<13> 
+ B_BLB_N<12> B_BLB_N<11> B_BLB_N<10> B_BLB_N<9> B_BLB_N<8> B_CA<3> B_CA<2> B_CA<1> B_CA<0> 
+ B_CB<3> B_CB<2> B_CB<1> B_CB<0> B_MA<3> B_MA<2> B_MA<1> B_MA<0> B_MB<3> 
+ B_MB<2> B_MB<1> B_MB<0> B_TM_PREA_N B_TM_PREB_N BWENA_INT<1> BWENB_INT<1> CLK_DQA CLK_DQA_N 
+ CLK_DQB CLK_DQB_N DA_INT<1> DB_INT<1> NET019 NET018 NET10 NET11 LWEA 
+ LWEB QA_INT<1> QB_INT<1> SA_PREA_N SA_PREB_N SAEA_N SAEB_N T_BLA<15> T_BLA<14> 
+ T_BLA<13> T_BLA<12> T_BLA<11> T_BLA<10> T_BLA<9> T_BLA<8> T_BLA_N<15> T_BLA_N<14> T_BLA_N<13> 
+ T_BLA_N<12> T_BLA_N<11> T_BLA_N<10> T_BLA_N<9> T_BLA_N<8> T_BLB<15> T_BLB<14> T_BLB<13> T_BLB<12> 
+ T_BLB<11> T_BLB<10> T_BLB<9> T_BLB<8> T_BLB_N<15> T_BLB_N<14> T_BLB_N<13> T_BLB_N<12> T_BLB_N<11> 
+ T_BLB_N<10> T_BLB_N<9> T_BLB_N<8> T_CA<3> T_CA<2> T_CA<1> T_CA<0> T_CB<3> T_CB<2> 
+ T_CB<1> T_CB<0> T_MA<3> T_MA<2> T_MA<1> T_MA<0> T_MB<3> T_MB<2> T_MB<1> 
+ T_MB<0> T_TM_PREA_N T_TM_PREB_N VDD VSS  / xmc55_dps_localc8io_bw
XAR_TOP<7>
+ T_BLA<15> T_BLA<14> T_BLA_N<15> T_BLA_N<14> T_BLB<15> T_BLB<14> T_BLB_N<15> T_BLB_N<14> VSS 
+ VDD T_WLA<255> T_WLA<254> T_WLA<253> T_WLA<252> T_WLA<251> T_WLA<250> T_WLA<249> T_WLA<248> 
+ T_WLA<247> T_WLA<246> T_WLA<245> T_WLA<244> T_WLA<243> T_WLA<242> T_WLA<241> T_WLA<240> T_WLA<239> 
+ T_WLA<238> T_WLA<237> T_WLA<236> T_WLA<235> T_WLA<234> T_WLA<233> T_WLA<232> T_WLA<231> T_WLA<230> 
+ T_WLA<229> T_WLA<228> T_WLA<227> T_WLA<226> T_WLA<225> T_WLA<224> T_WLA<223> T_WLA<222> T_WLA<221> 
+ T_WLA<220> T_WLA<219> T_WLA<218> T_WLA<217> T_WLA<216> T_WLA<215> T_WLA<214> T_WLA<213> T_WLA<212> 
+ T_WLA<211> T_WLA<210> T_WLA<209> T_WLA<208> T_WLA<207> T_WLA<206> T_WLA<205> T_WLA<204> T_WLA<203> 
+ T_WLA<202> T_WLA<201> T_WLA<200> T_WLA<199> T_WLA<198> T_WLA<197> T_WLA<196> T_WLA<195> T_WLA<194> 
+ T_WLA<193> T_WLA<192> T_WLA<191> T_WLA<190> T_WLA<189> T_WLA<188> T_WLA<187> T_WLA<186> T_WLA<185> 
+ T_WLA<184> T_WLA<183> T_WLA<182> T_WLA<181> T_WLA<180> T_WLA<179> T_WLA<178> T_WLA<177> T_WLA<176> 
+ T_WLA<175> T_WLA<174> T_WLA<173> T_WLA<172> T_WLA<171> T_WLA<170> T_WLA<169> T_WLA<168> T_WLA<167> 
+ T_WLA<166> T_WLA<165> T_WLA<164> T_WLA<163> T_WLA<162> T_WLA<161> T_WLA<160> T_WLA<159> T_WLA<158> 
+ T_WLA<157> T_WLA<156> T_WLA<155> T_WLA<154> T_WLA<153> T_WLA<152> T_WLA<151> T_WLA<150> T_WLA<149> 
+ T_WLA<148> T_WLA<147> T_WLA<146> T_WLA<145> T_WLA<144> T_WLA<143> T_WLA<142> T_WLA<141> T_WLA<140> 
+ T_WLA<139> T_WLA<138> T_WLA<137> T_WLA<136> T_WLA<135> T_WLA<134> T_WLA<133> T_WLA<132> T_WLA<131> 
+ T_WLA<130> T_WLA<129> T_WLA<128> T_WLA<127> T_WLA<126> T_WLA<125> T_WLA<124> T_WLA<123> T_WLA<122> 
+ T_WLA<121> T_WLA<120> T_WLA<119> T_WLA<118> T_WLA<117> T_WLA<116> T_WLA<115> T_WLA<114> T_WLA<113> 
+ T_WLA<112> T_WLA<111> T_WLA<110> T_WLA<109> T_WLA<108> T_WLA<107> T_WLA<106> T_WLA<105> T_WLA<104> 
+ T_WLA<103> T_WLA<102> T_WLA<101> T_WLA<100> T_WLA<99> T_WLA<98> T_WLA<97> T_WLA<96> T_WLA<95> 
+ T_WLA<94> T_WLA<93> T_WLA<92> T_WLA<91> T_WLA<90> T_WLA<89> T_WLA<88> T_WLA<87> T_WLA<86> 
+ T_WLA<85> T_WLA<84> T_WLA<83> T_WLA<82> T_WLA<81> T_WLA<80> T_WLA<79> T_WLA<78> T_WLA<77> 
+ T_WLA<76> T_WLA<75> T_WLA<74> T_WLA<73> T_WLA<72> T_WLA<71> T_WLA<70> T_WLA<69> T_WLA<68> 
+ T_WLA<67> T_WLA<66> T_WLA<65> T_WLA<64> T_WLA<63> T_WLA<62> T_WLA<61> T_WLA<60> T_WLA<59> 
+ T_WLA<58> T_WLA<57> T_WLA<56> T_WLA<55> T_WLA<54> T_WLA<53> T_WLA<52> T_WLA<51> T_WLA<50> 
+ T_WLA<49> T_WLA<48> T_WLA<47> T_WLA<46> T_WLA<45> T_WLA<44> T_WLA<43> T_WLA<42> T_WLA<41> 
+ T_WLA<40> T_WLA<39> T_WLA<38> T_WLA<37> T_WLA<36> T_WLA<35> T_WLA<34> T_WLA<33> T_WLA<32> 
+ T_WLA<31> T_WLA<30> T_WLA<29> T_WLA<28> T_WLA<27> T_WLA<26> T_WLA<25> T_WLA<24> T_WLA<23> 
+ T_WLA<22> T_WLA<21> T_WLA<20> T_WLA<19> T_WLA<18> T_WLA<17> T_WLA<16> T_WLA<15> T_WLA<14> 
+ T_WLA<13> T_WLA<12> T_WLA<11> T_WLA<10> T_WLA<9> T_WLA<8> T_WLA<7> T_WLA<6> T_WLA<5> 
+ T_WLA<4> T_WLA<3> T_WLA<2> T_WLA<1> T_WLA<0> T_WLB<255> T_WLB<254> T_WLB<253> T_WLB<252> 
+ T_WLB<251> T_WLB<250> T_WLB<249> T_WLB<248> T_WLB<247> T_WLB<246> T_WLB<245> T_WLB<244> T_WLB<243> 
+ T_WLB<242> T_WLB<241> T_WLB<240> T_WLB<239> T_WLB<238> T_WLB<237> T_WLB<236> T_WLB<235> T_WLB<234> 
+ T_WLB<233> T_WLB<232> T_WLB<231> T_WLB<230> T_WLB<229> T_WLB<228> T_WLB<227> T_WLB<226> T_WLB<225> 
+ T_WLB<224> T_WLB<223> T_WLB<222> T_WLB<221> T_WLB<220> T_WLB<219> T_WLB<218> T_WLB<217> T_WLB<216> 
+ T_WLB<215> T_WLB<214> T_WLB<213> T_WLB<212> T_WLB<211> T_WLB<210> T_WLB<209> T_WLB<208> T_WLB<207> 
+ T_WLB<206> T_WLB<205> T_WLB<204> T_WLB<203> T_WLB<202> T_WLB<201> T_WLB<200> T_WLB<199> T_WLB<198> 
+ T_WLB<197> T_WLB<196> T_WLB<195> T_WLB<194> T_WLB<193> T_WLB<192> T_WLB<191> T_WLB<190> T_WLB<189> 
+ T_WLB<188> T_WLB<187> T_WLB<186> T_WLB<185> T_WLB<184> T_WLB<183> T_WLB<182> T_WLB<181> T_WLB<180> 
+ T_WLB<179> T_WLB<178> T_WLB<177> T_WLB<176> T_WLB<175> T_WLB<174> T_WLB<173> T_WLB<172> T_WLB<171> 
+ T_WLB<170> T_WLB<169> T_WLB<168> T_WLB<167> T_WLB<166> T_WLB<165> T_WLB<164> T_WLB<163> T_WLB<162> 
+ T_WLB<161> T_WLB<160> T_WLB<159> T_WLB<158> T_WLB<157> T_WLB<156> T_WLB<155> T_WLB<154> T_WLB<153> 
+ T_WLB<152> T_WLB<151> T_WLB<150> T_WLB<149> T_WLB<148> T_WLB<147> T_WLB<146> T_WLB<145> T_WLB<144> 
+ T_WLB<143> T_WLB<142> T_WLB<141> T_WLB<140> T_WLB<139> T_WLB<138> T_WLB<137> T_WLB<136> T_WLB<135> 
+ T_WLB<134> T_WLB<133> T_WLB<132> T_WLB<131> T_WLB<130> T_WLB<129> T_WLB<128> T_WLB<127> T_WLB<126> 
+ T_WLB<125> T_WLB<124> T_WLB<123> T_WLB<122> T_WLB<121> T_WLB<120> T_WLB<119> T_WLB<118> T_WLB<117> 
+ T_WLB<116> T_WLB<115> T_WLB<114> T_WLB<113> T_WLB<112> T_WLB<111> T_WLB<110> T_WLB<109> T_WLB<108> 
+ T_WLB<107> T_WLB<106> T_WLB<105> T_WLB<104> T_WLB<103> T_WLB<102> T_WLB<101> T_WLB<100> T_WLB<99> 
+ T_WLB<98> T_WLB<97> T_WLB<96> T_WLB<95> T_WLB<94> T_WLB<93> T_WLB<92> T_WLB<91> T_WLB<90> 
+ T_WLB<89> T_WLB<88> T_WLB<87> T_WLB<86> T_WLB<85> T_WLB<84> T_WLB<83> T_WLB<82> T_WLB<81> 
+ T_WLB<80> T_WLB<79> T_WLB<78> T_WLB<77> T_WLB<76> T_WLB<75> T_WLB<74> T_WLB<73> T_WLB<72> 
+ T_WLB<71> T_WLB<70> T_WLB<69> T_WLB<68> T_WLB<67> T_WLB<66> T_WLB<65> T_WLB<64> T_WLB<63> 
+ T_WLB<62> T_WLB<61> T_WLB<60> T_WLB<59> T_WLB<58> T_WLB<57> T_WLB<56> T_WLB<55> T_WLB<54> 
+ T_WLB<53> T_WLB<52> T_WLB<51> T_WLB<50> T_WLB<49> T_WLB<48> T_WLB<47> T_WLB<46> T_WLB<45> 
+ T_WLB<44> T_WLB<43> T_WLB<42> T_WLB<41> T_WLB<40> T_WLB<39> T_WLB<38> T_WLB<37> T_WLB<36> 
+ T_WLB<35> T_WLB<34> T_WLB<33> T_WLB<32> T_WLB<31> T_WLB<30> T_WLB<29> T_WLB<28> T_WLB<27> 
+ T_WLB<26> T_WLB<25> T_WLB<24> T_WLB<23> T_WLB<22> T_WLB<21> T_WLB<20> T_WLB<19> T_WLB<18> 
+ T_WLB<17> T_WLB<16> T_WLB<15> T_WLB<14> T_WLB<13> T_WLB<12> T_WLB<11> T_WLB<10> T_WLB<9> 
+ T_WLB<8> T_WLB<7> T_WLB<6> T_WLB<5> T_WLB<4> T_WLB<3> T_WLB<2> T_WLB<1> T_WLB<0> 
+  / dpram16x4096_AR_COLX8_ROWX256
XAR_BOT<7>
+ B_BLA<15> B_BLA<14> B_BLA_N<15> B_BLA_N<14> B_BLB<15> B_BLB<14> B_BLB_N<15> B_BLB_N<14> VSS 
+ VDD B_WLA<255> B_WLA<254> B_WLA<253> B_WLA<252> B_WLA<251> B_WLA<250> B_WLA<249> B_WLA<248> 
+ B_WLA<247> B_WLA<246> B_WLA<245> B_WLA<244> B_WLA<243> B_WLA<242> B_WLA<241> B_WLA<240> B_WLA<239> 
+ B_WLA<238> B_WLA<237> B_WLA<236> B_WLA<235> B_WLA<234> B_WLA<233> B_WLA<232> B_WLA<231> B_WLA<230> 
+ B_WLA<229> B_WLA<228> B_WLA<227> B_WLA<226> B_WLA<225> B_WLA<224> B_WLA<223> B_WLA<222> B_WLA<221> 
+ B_WLA<220> B_WLA<219> B_WLA<218> B_WLA<217> B_WLA<216> B_WLA<215> B_WLA<214> B_WLA<213> B_WLA<212> 
+ B_WLA<211> B_WLA<210> B_WLA<209> B_WLA<208> B_WLA<207> B_WLA<206> B_WLA<205> B_WLA<204> B_WLA<203> 
+ B_WLA<202> B_WLA<201> B_WLA<200> B_WLA<199> B_WLA<198> B_WLA<197> B_WLA<196> B_WLA<195> B_WLA<194> 
+ B_WLA<193> B_WLA<192> B_WLA<191> B_WLA<190> B_WLA<189> B_WLA<188> B_WLA<187> B_WLA<186> B_WLA<185> 
+ B_WLA<184> B_WLA<183> B_WLA<182> B_WLA<181> B_WLA<180> B_WLA<179> B_WLA<178> B_WLA<177> B_WLA<176> 
+ B_WLA<175> B_WLA<174> B_WLA<173> B_WLA<172> B_WLA<171> B_WLA<170> B_WLA<169> B_WLA<168> B_WLA<167> 
+ B_WLA<166> B_WLA<165> B_WLA<164> B_WLA<163> B_WLA<162> B_WLA<161> B_WLA<160> B_WLA<159> B_WLA<158> 
+ B_WLA<157> B_WLA<156> B_WLA<155> B_WLA<154> B_WLA<153> B_WLA<152> B_WLA<151> B_WLA<150> B_WLA<149> 
+ B_WLA<148> B_WLA<147> B_WLA<146> B_WLA<145> B_WLA<144> B_WLA<143> B_WLA<142> B_WLA<141> B_WLA<140> 
+ B_WLA<139> B_WLA<138> B_WLA<137> B_WLA<136> B_WLA<135> B_WLA<134> B_WLA<133> B_WLA<132> B_WLA<131> 
+ B_WLA<130> B_WLA<129> B_WLA<128> B_WLA<127> B_WLA<126> B_WLA<125> B_WLA<124> B_WLA<123> B_WLA<122> 
+ B_WLA<121> B_WLA<120> B_WLA<119> B_WLA<118> B_WLA<117> B_WLA<116> B_WLA<115> B_WLA<114> B_WLA<113> 
+ B_WLA<112> B_WLA<111> B_WLA<110> B_WLA<109> B_WLA<108> B_WLA<107> B_WLA<106> B_WLA<105> B_WLA<104> 
+ B_WLA<103> B_WLA<102> B_WLA<101> B_WLA<100> B_WLA<99> B_WLA<98> B_WLA<97> B_WLA<96> B_WLA<95> 
+ B_WLA<94> B_WLA<93> B_WLA<92> B_WLA<91> B_WLA<90> B_WLA<89> B_WLA<88> B_WLA<87> B_WLA<86> 
+ B_WLA<85> B_WLA<84> B_WLA<83> B_WLA<82> B_WLA<81> B_WLA<80> B_WLA<79> B_WLA<78> B_WLA<77> 
+ B_WLA<76> B_WLA<75> B_WLA<74> B_WLA<73> B_WLA<72> B_WLA<71> B_WLA<70> B_WLA<69> B_WLA<68> 
+ B_WLA<67> B_WLA<66> B_WLA<65> B_WLA<64> B_WLA<63> B_WLA<62> B_WLA<61> B_WLA<60> B_WLA<59> 
+ B_WLA<58> B_WLA<57> B_WLA<56> B_WLA<55> B_WLA<54> B_WLA<53> B_WLA<52> B_WLA<51> B_WLA<50> 
+ B_WLA<49> B_WLA<48> B_WLA<47> B_WLA<46> B_WLA<45> B_WLA<44> B_WLA<43> B_WLA<42> B_WLA<41> 
+ B_WLA<40> B_WLA<39> B_WLA<38> B_WLA<37> B_WLA<36> B_WLA<35> B_WLA<34> B_WLA<33> B_WLA<32> 
+ B_WLA<31> B_WLA<30> B_WLA<29> B_WLA<28> B_WLA<27> B_WLA<26> B_WLA<25> B_WLA<24> B_WLA<23> 
+ B_WLA<22> B_WLA<21> B_WLA<20> B_WLA<19> B_WLA<18> B_WLA<17> B_WLA<16> B_WLA<15> B_WLA<14> 
+ B_WLA<13> B_WLA<12> B_WLA<11> B_WLA<10> B_WLA<9> B_WLA<8> B_WLA<7> B_WLA<6> B_WLA<5> 
+ B_WLA<4> B_WLA<3> B_WLA<2> B_WLA<1> B_WLA<0> B_WLB<255> B_WLB<254> B_WLB<253> B_WLB<252> 
+ B_WLB<251> B_WLB<250> B_WLB<249> B_WLB<248> B_WLB<247> B_WLB<246> B_WLB<245> B_WLB<244> B_WLB<243> 
+ B_WLB<242> B_WLB<241> B_WLB<240> B_WLB<239> B_WLB<238> B_WLB<237> B_WLB<236> B_WLB<235> B_WLB<234> 
+ B_WLB<233> B_WLB<232> B_WLB<231> B_WLB<230> B_WLB<229> B_WLB<228> B_WLB<227> B_WLB<226> B_WLB<225> 
+ B_WLB<224> B_WLB<223> B_WLB<222> B_WLB<221> B_WLB<220> B_WLB<219> B_WLB<218> B_WLB<217> B_WLB<216> 
+ B_WLB<215> B_WLB<214> B_WLB<213> B_WLB<212> B_WLB<211> B_WLB<210> B_WLB<209> B_WLB<208> B_WLB<207> 
+ B_WLB<206> B_WLB<205> B_WLB<204> B_WLB<203> B_WLB<202> B_WLB<201> B_WLB<200> B_WLB<199> B_WLB<198> 
+ B_WLB<197> B_WLB<196> B_WLB<195> B_WLB<194> B_WLB<193> B_WLB<192> B_WLB<191> B_WLB<190> B_WLB<189> 
+ B_WLB<188> B_WLB<187> B_WLB<186> B_WLB<185> B_WLB<184> B_WLB<183> B_WLB<182> B_WLB<181> B_WLB<180> 
+ B_WLB<179> B_WLB<178> B_WLB<177> B_WLB<176> B_WLB<175> B_WLB<174> B_WLB<173> B_WLB<172> B_WLB<171> 
+ B_WLB<170> B_WLB<169> B_WLB<168> B_WLB<167> B_WLB<166> B_WLB<165> B_WLB<164> B_WLB<163> B_WLB<162> 
+ B_WLB<161> B_WLB<160> B_WLB<159> B_WLB<158> B_WLB<157> B_WLB<156> B_WLB<155> B_WLB<154> B_WLB<153> 
+ B_WLB<152> B_WLB<151> B_WLB<150> B_WLB<149> B_WLB<148> B_WLB<147> B_WLB<146> B_WLB<145> B_WLB<144> 
+ B_WLB<143> B_WLB<142> B_WLB<141> B_WLB<140> B_WLB<139> B_WLB<138> B_WLB<137> B_WLB<136> B_WLB<135> 
+ B_WLB<134> B_WLB<133> B_WLB<132> B_WLB<131> B_WLB<130> B_WLB<129> B_WLB<128> B_WLB<127> B_WLB<126> 
+ B_WLB<125> B_WLB<124> B_WLB<123> B_WLB<122> B_WLB<121> B_WLB<120> B_WLB<119> B_WLB<118> B_WLB<117> 
+ B_WLB<116> B_WLB<115> B_WLB<114> B_WLB<113> B_WLB<112> B_WLB<111> B_WLB<110> B_WLB<109> B_WLB<108> 
+ B_WLB<107> B_WLB<106> B_WLB<105> B_WLB<104> B_WLB<103> B_WLB<102> B_WLB<101> B_WLB<100> B_WLB<99> 
+ B_WLB<98> B_WLB<97> B_WLB<96> B_WLB<95> B_WLB<94> B_WLB<93> B_WLB<92> B_WLB<91> B_WLB<90> 
+ B_WLB<89> B_WLB<88> B_WLB<87> B_WLB<86> B_WLB<85> B_WLB<84> B_WLB<83> B_WLB<82> B_WLB<81> 
+ B_WLB<80> B_WLB<79> B_WLB<78> B_WLB<77> B_WLB<76> B_WLB<75> B_WLB<74> B_WLB<73> B_WLB<72> 
+ B_WLB<71> B_WLB<70> B_WLB<69> B_WLB<68> B_WLB<67> B_WLB<66> B_WLB<65> B_WLB<64> B_WLB<63> 
+ B_WLB<62> B_WLB<61> B_WLB<60> B_WLB<59> B_WLB<58> B_WLB<57> B_WLB<56> B_WLB<55> B_WLB<54> 
+ B_WLB<53> B_WLB<52> B_WLB<51> B_WLB<50> B_WLB<49> B_WLB<48> B_WLB<47> B_WLB<46> B_WLB<45> 
+ B_WLB<44> B_WLB<43> B_WLB<42> B_WLB<41> B_WLB<40> B_WLB<39> B_WLB<38> B_WLB<37> B_WLB<36> 
+ B_WLB<35> B_WLB<34> B_WLB<33> B_WLB<32> B_WLB<31> B_WLB<30> B_WLB<29> B_WLB<28> B_WLB<27> 
+ B_WLB<26> B_WLB<25> B_WLB<24> B_WLB<23> B_WLB<22> B_WLB<21> B_WLB<20> B_WLB<19> B_WLB<18> 
+ B_WLB<17> B_WLB<16> B_WLB<15> B_WLB<14> B_WLB<13> B_WLB<12> B_WLB<11> B_WLB<10> B_WLB<9> 
+ B_WLB<8> B_WLB<7> B_WLB<6> B_WLB<5> B_WLB<4> B_WLB<3> B_WLB<2> B_WLB<1> B_WLB<0> 
+  / dpram16x4096_AR_COLX8_ROWX256
XAR_TOP<6>
+ T_BLA<13> T_BLA<12> T_BLA_N<13> T_BLA_N<12> T_BLB<13> T_BLB<12> T_BLB_N<13> T_BLB_N<12> VSS 
+ VDD T_WLA<255> T_WLA<254> T_WLA<253> T_WLA<252> T_WLA<251> T_WLA<250> T_WLA<249> T_WLA<248> 
+ T_WLA<247> T_WLA<246> T_WLA<245> T_WLA<244> T_WLA<243> T_WLA<242> T_WLA<241> T_WLA<240> T_WLA<239> 
+ T_WLA<238> T_WLA<237> T_WLA<236> T_WLA<235> T_WLA<234> T_WLA<233> T_WLA<232> T_WLA<231> T_WLA<230> 
+ T_WLA<229> T_WLA<228> T_WLA<227> T_WLA<226> T_WLA<225> T_WLA<224> T_WLA<223> T_WLA<222> T_WLA<221> 
+ T_WLA<220> T_WLA<219> T_WLA<218> T_WLA<217> T_WLA<216> T_WLA<215> T_WLA<214> T_WLA<213> T_WLA<212> 
+ T_WLA<211> T_WLA<210> T_WLA<209> T_WLA<208> T_WLA<207> T_WLA<206> T_WLA<205> T_WLA<204> T_WLA<203> 
+ T_WLA<202> T_WLA<201> T_WLA<200> T_WLA<199> T_WLA<198> T_WLA<197> T_WLA<196> T_WLA<195> T_WLA<194> 
+ T_WLA<193> T_WLA<192> T_WLA<191> T_WLA<190> T_WLA<189> T_WLA<188> T_WLA<187> T_WLA<186> T_WLA<185> 
+ T_WLA<184> T_WLA<183> T_WLA<182> T_WLA<181> T_WLA<180> T_WLA<179> T_WLA<178> T_WLA<177> T_WLA<176> 
+ T_WLA<175> T_WLA<174> T_WLA<173> T_WLA<172> T_WLA<171> T_WLA<170> T_WLA<169> T_WLA<168> T_WLA<167> 
+ T_WLA<166> T_WLA<165> T_WLA<164> T_WLA<163> T_WLA<162> T_WLA<161> T_WLA<160> T_WLA<159> T_WLA<158> 
+ T_WLA<157> T_WLA<156> T_WLA<155> T_WLA<154> T_WLA<153> T_WLA<152> T_WLA<151> T_WLA<150> T_WLA<149> 
+ T_WLA<148> T_WLA<147> T_WLA<146> T_WLA<145> T_WLA<144> T_WLA<143> T_WLA<142> T_WLA<141> T_WLA<140> 
+ T_WLA<139> T_WLA<138> T_WLA<137> T_WLA<136> T_WLA<135> T_WLA<134> T_WLA<133> T_WLA<132> T_WLA<131> 
+ T_WLA<130> T_WLA<129> T_WLA<128> T_WLA<127> T_WLA<126> T_WLA<125> T_WLA<124> T_WLA<123> T_WLA<122> 
+ T_WLA<121> T_WLA<120> T_WLA<119> T_WLA<118> T_WLA<117> T_WLA<116> T_WLA<115> T_WLA<114> T_WLA<113> 
+ T_WLA<112> T_WLA<111> T_WLA<110> T_WLA<109> T_WLA<108> T_WLA<107> T_WLA<106> T_WLA<105> T_WLA<104> 
+ T_WLA<103> T_WLA<102> T_WLA<101> T_WLA<100> T_WLA<99> T_WLA<98> T_WLA<97> T_WLA<96> T_WLA<95> 
+ T_WLA<94> T_WLA<93> T_WLA<92> T_WLA<91> T_WLA<90> T_WLA<89> T_WLA<88> T_WLA<87> T_WLA<86> 
+ T_WLA<85> T_WLA<84> T_WLA<83> T_WLA<82> T_WLA<81> T_WLA<80> T_WLA<79> T_WLA<78> T_WLA<77> 
+ T_WLA<76> T_WLA<75> T_WLA<74> T_WLA<73> T_WLA<72> T_WLA<71> T_WLA<70> T_WLA<69> T_WLA<68> 
+ T_WLA<67> T_WLA<66> T_WLA<65> T_WLA<64> T_WLA<63> T_WLA<62> T_WLA<61> T_WLA<60> T_WLA<59> 
+ T_WLA<58> T_WLA<57> T_WLA<56> T_WLA<55> T_WLA<54> T_WLA<53> T_WLA<52> T_WLA<51> T_WLA<50> 
+ T_WLA<49> T_WLA<48> T_WLA<47> T_WLA<46> T_WLA<45> T_WLA<44> T_WLA<43> T_WLA<42> T_WLA<41> 
+ T_WLA<40> T_WLA<39> T_WLA<38> T_WLA<37> T_WLA<36> T_WLA<35> T_WLA<34> T_WLA<33> T_WLA<32> 
+ T_WLA<31> T_WLA<30> T_WLA<29> T_WLA<28> T_WLA<27> T_WLA<26> T_WLA<25> T_WLA<24> T_WLA<23> 
+ T_WLA<22> T_WLA<21> T_WLA<20> T_WLA<19> T_WLA<18> T_WLA<17> T_WLA<16> T_WLA<15> T_WLA<14> 
+ T_WLA<13> T_WLA<12> T_WLA<11> T_WLA<10> T_WLA<9> T_WLA<8> T_WLA<7> T_WLA<6> T_WLA<5> 
+ T_WLA<4> T_WLA<3> T_WLA<2> T_WLA<1> T_WLA<0> T_WLB<255> T_WLB<254> T_WLB<253> T_WLB<252> 
+ T_WLB<251> T_WLB<250> T_WLB<249> T_WLB<248> T_WLB<247> T_WLB<246> T_WLB<245> T_WLB<244> T_WLB<243> 
+ T_WLB<242> T_WLB<241> T_WLB<240> T_WLB<239> T_WLB<238> T_WLB<237> T_WLB<236> T_WLB<235> T_WLB<234> 
+ T_WLB<233> T_WLB<232> T_WLB<231> T_WLB<230> T_WLB<229> T_WLB<228> T_WLB<227> T_WLB<226> T_WLB<225> 
+ T_WLB<224> T_WLB<223> T_WLB<222> T_WLB<221> T_WLB<220> T_WLB<219> T_WLB<218> T_WLB<217> T_WLB<216> 
+ T_WLB<215> T_WLB<214> T_WLB<213> T_WLB<212> T_WLB<211> T_WLB<210> T_WLB<209> T_WLB<208> T_WLB<207> 
+ T_WLB<206> T_WLB<205> T_WLB<204> T_WLB<203> T_WLB<202> T_WLB<201> T_WLB<200> T_WLB<199> T_WLB<198> 
+ T_WLB<197> T_WLB<196> T_WLB<195> T_WLB<194> T_WLB<193> T_WLB<192> T_WLB<191> T_WLB<190> T_WLB<189> 
+ T_WLB<188> T_WLB<187> T_WLB<186> T_WLB<185> T_WLB<184> T_WLB<183> T_WLB<182> T_WLB<181> T_WLB<180> 
+ T_WLB<179> T_WLB<178> T_WLB<177> T_WLB<176> T_WLB<175> T_WLB<174> T_WLB<173> T_WLB<172> T_WLB<171> 
+ T_WLB<170> T_WLB<169> T_WLB<168> T_WLB<167> T_WLB<166> T_WLB<165> T_WLB<164> T_WLB<163> T_WLB<162> 
+ T_WLB<161> T_WLB<160> T_WLB<159> T_WLB<158> T_WLB<157> T_WLB<156> T_WLB<155> T_WLB<154> T_WLB<153> 
+ T_WLB<152> T_WLB<151> T_WLB<150> T_WLB<149> T_WLB<148> T_WLB<147> T_WLB<146> T_WLB<145> T_WLB<144> 
+ T_WLB<143> T_WLB<142> T_WLB<141> T_WLB<140> T_WLB<139> T_WLB<138> T_WLB<137> T_WLB<136> T_WLB<135> 
+ T_WLB<134> T_WLB<133> T_WLB<132> T_WLB<131> T_WLB<130> T_WLB<129> T_WLB<128> T_WLB<127> T_WLB<126> 
+ T_WLB<125> T_WLB<124> T_WLB<123> T_WLB<122> T_WLB<121> T_WLB<120> T_WLB<119> T_WLB<118> T_WLB<117> 
+ T_WLB<116> T_WLB<115> T_WLB<114> T_WLB<113> T_WLB<112> T_WLB<111> T_WLB<110> T_WLB<109> T_WLB<108> 
+ T_WLB<107> T_WLB<106> T_WLB<105> T_WLB<104> T_WLB<103> T_WLB<102> T_WLB<101> T_WLB<100> T_WLB<99> 
+ T_WLB<98> T_WLB<97> T_WLB<96> T_WLB<95> T_WLB<94> T_WLB<93> T_WLB<92> T_WLB<91> T_WLB<90> 
+ T_WLB<89> T_WLB<88> T_WLB<87> T_WLB<86> T_WLB<85> T_WLB<84> T_WLB<83> T_WLB<82> T_WLB<81> 
+ T_WLB<80> T_WLB<79> T_WLB<78> T_WLB<77> T_WLB<76> T_WLB<75> T_WLB<74> T_WLB<73> T_WLB<72> 
+ T_WLB<71> T_WLB<70> T_WLB<69> T_WLB<68> T_WLB<67> T_WLB<66> T_WLB<65> T_WLB<64> T_WLB<63> 
+ T_WLB<62> T_WLB<61> T_WLB<60> T_WLB<59> T_WLB<58> T_WLB<57> T_WLB<56> T_WLB<55> T_WLB<54> 
+ T_WLB<53> T_WLB<52> T_WLB<51> T_WLB<50> T_WLB<49> T_WLB<48> T_WLB<47> T_WLB<46> T_WLB<45> 
+ T_WLB<44> T_WLB<43> T_WLB<42> T_WLB<41> T_WLB<40> T_WLB<39> T_WLB<38> T_WLB<37> T_WLB<36> 
+ T_WLB<35> T_WLB<34> T_WLB<33> T_WLB<32> T_WLB<31> T_WLB<30> T_WLB<29> T_WLB<28> T_WLB<27> 
+ T_WLB<26> T_WLB<25> T_WLB<24> T_WLB<23> T_WLB<22> T_WLB<21> T_WLB<20> T_WLB<19> T_WLB<18> 
+ T_WLB<17> T_WLB<16> T_WLB<15> T_WLB<14> T_WLB<13> T_WLB<12> T_WLB<11> T_WLB<10> T_WLB<9> 
+ T_WLB<8> T_WLB<7> T_WLB<6> T_WLB<5> T_WLB<4> T_WLB<3> T_WLB<2> T_WLB<1> T_WLB<0> 
+  / dpram16x4096_AR_COLX8_ROWX256
XAR_BOT<6>
+ B_BLA<13> B_BLA<12> B_BLA_N<13> B_BLA_N<12> B_BLB<13> B_BLB<12> B_BLB_N<13> B_BLB_N<12> VSS 
+ VDD B_WLA<255> B_WLA<254> B_WLA<253> B_WLA<252> B_WLA<251> B_WLA<250> B_WLA<249> B_WLA<248> 
+ B_WLA<247> B_WLA<246> B_WLA<245> B_WLA<244> B_WLA<243> B_WLA<242> B_WLA<241> B_WLA<240> B_WLA<239> 
+ B_WLA<238> B_WLA<237> B_WLA<236> B_WLA<235> B_WLA<234> B_WLA<233> B_WLA<232> B_WLA<231> B_WLA<230> 
+ B_WLA<229> B_WLA<228> B_WLA<227> B_WLA<226> B_WLA<225> B_WLA<224> B_WLA<223> B_WLA<222> B_WLA<221> 
+ B_WLA<220> B_WLA<219> B_WLA<218> B_WLA<217> B_WLA<216> B_WLA<215> B_WLA<214> B_WLA<213> B_WLA<212> 
+ B_WLA<211> B_WLA<210> B_WLA<209> B_WLA<208> B_WLA<207> B_WLA<206> B_WLA<205> B_WLA<204> B_WLA<203> 
+ B_WLA<202> B_WLA<201> B_WLA<200> B_WLA<199> B_WLA<198> B_WLA<197> B_WLA<196> B_WLA<195> B_WLA<194> 
+ B_WLA<193> B_WLA<192> B_WLA<191> B_WLA<190> B_WLA<189> B_WLA<188> B_WLA<187> B_WLA<186> B_WLA<185> 
+ B_WLA<184> B_WLA<183> B_WLA<182> B_WLA<181> B_WLA<180> B_WLA<179> B_WLA<178> B_WLA<177> B_WLA<176> 
+ B_WLA<175> B_WLA<174> B_WLA<173> B_WLA<172> B_WLA<171> B_WLA<170> B_WLA<169> B_WLA<168> B_WLA<167> 
+ B_WLA<166> B_WLA<165> B_WLA<164> B_WLA<163> B_WLA<162> B_WLA<161> B_WLA<160> B_WLA<159> B_WLA<158> 
+ B_WLA<157> B_WLA<156> B_WLA<155> B_WLA<154> B_WLA<153> B_WLA<152> B_WLA<151> B_WLA<150> B_WLA<149> 
+ B_WLA<148> B_WLA<147> B_WLA<146> B_WLA<145> B_WLA<144> B_WLA<143> B_WLA<142> B_WLA<141> B_WLA<140> 
+ B_WLA<139> B_WLA<138> B_WLA<137> B_WLA<136> B_WLA<135> B_WLA<134> B_WLA<133> B_WLA<132> B_WLA<131> 
+ B_WLA<130> B_WLA<129> B_WLA<128> B_WLA<127> B_WLA<126> B_WLA<125> B_WLA<124> B_WLA<123> B_WLA<122> 
+ B_WLA<121> B_WLA<120> B_WLA<119> B_WLA<118> B_WLA<117> B_WLA<116> B_WLA<115> B_WLA<114> B_WLA<113> 
+ B_WLA<112> B_WLA<111> B_WLA<110> B_WLA<109> B_WLA<108> B_WLA<107> B_WLA<106> B_WLA<105> B_WLA<104> 
+ B_WLA<103> B_WLA<102> B_WLA<101> B_WLA<100> B_WLA<99> B_WLA<98> B_WLA<97> B_WLA<96> B_WLA<95> 
+ B_WLA<94> B_WLA<93> B_WLA<92> B_WLA<91> B_WLA<90> B_WLA<89> B_WLA<88> B_WLA<87> B_WLA<86> 
+ B_WLA<85> B_WLA<84> B_WLA<83> B_WLA<82> B_WLA<81> B_WLA<80> B_WLA<79> B_WLA<78> B_WLA<77> 
+ B_WLA<76> B_WLA<75> B_WLA<74> B_WLA<73> B_WLA<72> B_WLA<71> B_WLA<70> B_WLA<69> B_WLA<68> 
+ B_WLA<67> B_WLA<66> B_WLA<65> B_WLA<64> B_WLA<63> B_WLA<62> B_WLA<61> B_WLA<60> B_WLA<59> 
+ B_WLA<58> B_WLA<57> B_WLA<56> B_WLA<55> B_WLA<54> B_WLA<53> B_WLA<52> B_WLA<51> B_WLA<50> 
+ B_WLA<49> B_WLA<48> B_WLA<47> B_WLA<46> B_WLA<45> B_WLA<44> B_WLA<43> B_WLA<42> B_WLA<41> 
+ B_WLA<40> B_WLA<39> B_WLA<38> B_WLA<37> B_WLA<36> B_WLA<35> B_WLA<34> B_WLA<33> B_WLA<32> 
+ B_WLA<31> B_WLA<30> B_WLA<29> B_WLA<28> B_WLA<27> B_WLA<26> B_WLA<25> B_WLA<24> B_WLA<23> 
+ B_WLA<22> B_WLA<21> B_WLA<20> B_WLA<19> B_WLA<18> B_WLA<17> B_WLA<16> B_WLA<15> B_WLA<14> 
+ B_WLA<13> B_WLA<12> B_WLA<11> B_WLA<10> B_WLA<9> B_WLA<8> B_WLA<7> B_WLA<6> B_WLA<5> 
+ B_WLA<4> B_WLA<3> B_WLA<2> B_WLA<1> B_WLA<0> B_WLB<255> B_WLB<254> B_WLB<253> B_WLB<252> 
+ B_WLB<251> B_WLB<250> B_WLB<249> B_WLB<248> B_WLB<247> B_WLB<246> B_WLB<245> B_WLB<244> B_WLB<243> 
+ B_WLB<242> B_WLB<241> B_WLB<240> B_WLB<239> B_WLB<238> B_WLB<237> B_WLB<236> B_WLB<235> B_WLB<234> 
+ B_WLB<233> B_WLB<232> B_WLB<231> B_WLB<230> B_WLB<229> B_WLB<228> B_WLB<227> B_WLB<226> B_WLB<225> 
+ B_WLB<224> B_WLB<223> B_WLB<222> B_WLB<221> B_WLB<220> B_WLB<219> B_WLB<218> B_WLB<217> B_WLB<216> 
+ B_WLB<215> B_WLB<214> B_WLB<213> B_WLB<212> B_WLB<211> B_WLB<210> B_WLB<209> B_WLB<208> B_WLB<207> 
+ B_WLB<206> B_WLB<205> B_WLB<204> B_WLB<203> B_WLB<202> B_WLB<201> B_WLB<200> B_WLB<199> B_WLB<198> 
+ B_WLB<197> B_WLB<196> B_WLB<195> B_WLB<194> B_WLB<193> B_WLB<192> B_WLB<191> B_WLB<190> B_WLB<189> 
+ B_WLB<188> B_WLB<187> B_WLB<186> B_WLB<185> B_WLB<184> B_WLB<183> B_WLB<182> B_WLB<181> B_WLB<180> 
+ B_WLB<179> B_WLB<178> B_WLB<177> B_WLB<176> B_WLB<175> B_WLB<174> B_WLB<173> B_WLB<172> B_WLB<171> 
+ B_WLB<170> B_WLB<169> B_WLB<168> B_WLB<167> B_WLB<166> B_WLB<165> B_WLB<164> B_WLB<163> B_WLB<162> 
+ B_WLB<161> B_WLB<160> B_WLB<159> B_WLB<158> B_WLB<157> B_WLB<156> B_WLB<155> B_WLB<154> B_WLB<153> 
+ B_WLB<152> B_WLB<151> B_WLB<150> B_WLB<149> B_WLB<148> B_WLB<147> B_WLB<146> B_WLB<145> B_WLB<144> 
+ B_WLB<143> B_WLB<142> B_WLB<141> B_WLB<140> B_WLB<139> B_WLB<138> B_WLB<137> B_WLB<136> B_WLB<135> 
+ B_WLB<134> B_WLB<133> B_WLB<132> B_WLB<131> B_WLB<130> B_WLB<129> B_WLB<128> B_WLB<127> B_WLB<126> 
+ B_WLB<125> B_WLB<124> B_WLB<123> B_WLB<122> B_WLB<121> B_WLB<120> B_WLB<119> B_WLB<118> B_WLB<117> 
+ B_WLB<116> B_WLB<115> B_WLB<114> B_WLB<113> B_WLB<112> B_WLB<111> B_WLB<110> B_WLB<109> B_WLB<108> 
+ B_WLB<107> B_WLB<106> B_WLB<105> B_WLB<104> B_WLB<103> B_WLB<102> B_WLB<101> B_WLB<100> B_WLB<99> 
+ B_WLB<98> B_WLB<97> B_WLB<96> B_WLB<95> B_WLB<94> B_WLB<93> B_WLB<92> B_WLB<91> B_WLB<90> 
+ B_WLB<89> B_WLB<88> B_WLB<87> B_WLB<86> B_WLB<85> B_WLB<84> B_WLB<83> B_WLB<82> B_WLB<81> 
+ B_WLB<80> B_WLB<79> B_WLB<78> B_WLB<77> B_WLB<76> B_WLB<75> B_WLB<74> B_WLB<73> B_WLB<72> 
+ B_WLB<71> B_WLB<70> B_WLB<69> B_WLB<68> B_WLB<67> B_WLB<66> B_WLB<65> B_WLB<64> B_WLB<63> 
+ B_WLB<62> B_WLB<61> B_WLB<60> B_WLB<59> B_WLB<58> B_WLB<57> B_WLB<56> B_WLB<55> B_WLB<54> 
+ B_WLB<53> B_WLB<52> B_WLB<51> B_WLB<50> B_WLB<49> B_WLB<48> B_WLB<47> B_WLB<46> B_WLB<45> 
+ B_WLB<44> B_WLB<43> B_WLB<42> B_WLB<41> B_WLB<40> B_WLB<39> B_WLB<38> B_WLB<37> B_WLB<36> 
+ B_WLB<35> B_WLB<34> B_WLB<33> B_WLB<32> B_WLB<31> B_WLB<30> B_WLB<29> B_WLB<28> B_WLB<27> 
+ B_WLB<26> B_WLB<25> B_WLB<24> B_WLB<23> B_WLB<22> B_WLB<21> B_WLB<20> B_WLB<19> B_WLB<18> 
+ B_WLB<17> B_WLB<16> B_WLB<15> B_WLB<14> B_WLB<13> B_WLB<12> B_WLB<11> B_WLB<10> B_WLB<9> 
+ B_WLB<8> B_WLB<7> B_WLB<6> B_WLB<5> B_WLB<4> B_WLB<3> B_WLB<2> B_WLB<1> B_WLB<0> 
+  / dpram16x4096_AR_COLX8_ROWX256
XAR_TOP<5>
+ T_BLA<11> T_BLA<10> T_BLA_N<11> T_BLA_N<10> T_BLB<11> T_BLB<10> T_BLB_N<11> T_BLB_N<10> VSS 
+ VDD T_WLA<255> T_WLA<254> T_WLA<253> T_WLA<252> T_WLA<251> T_WLA<250> T_WLA<249> T_WLA<248> 
+ T_WLA<247> T_WLA<246> T_WLA<245> T_WLA<244> T_WLA<243> T_WLA<242> T_WLA<241> T_WLA<240> T_WLA<239> 
+ T_WLA<238> T_WLA<237> T_WLA<236> T_WLA<235> T_WLA<234> T_WLA<233> T_WLA<232> T_WLA<231> T_WLA<230> 
+ T_WLA<229> T_WLA<228> T_WLA<227> T_WLA<226> T_WLA<225> T_WLA<224> T_WLA<223> T_WLA<222> T_WLA<221> 
+ T_WLA<220> T_WLA<219> T_WLA<218> T_WLA<217> T_WLA<216> T_WLA<215> T_WLA<214> T_WLA<213> T_WLA<212> 
+ T_WLA<211> T_WLA<210> T_WLA<209> T_WLA<208> T_WLA<207> T_WLA<206> T_WLA<205> T_WLA<204> T_WLA<203> 
+ T_WLA<202> T_WLA<201> T_WLA<200> T_WLA<199> T_WLA<198> T_WLA<197> T_WLA<196> T_WLA<195> T_WLA<194> 
+ T_WLA<193> T_WLA<192> T_WLA<191> T_WLA<190> T_WLA<189> T_WLA<188> T_WLA<187> T_WLA<186> T_WLA<185> 
+ T_WLA<184> T_WLA<183> T_WLA<182> T_WLA<181> T_WLA<180> T_WLA<179> T_WLA<178> T_WLA<177> T_WLA<176> 
+ T_WLA<175> T_WLA<174> T_WLA<173> T_WLA<172> T_WLA<171> T_WLA<170> T_WLA<169> T_WLA<168> T_WLA<167> 
+ T_WLA<166> T_WLA<165> T_WLA<164> T_WLA<163> T_WLA<162> T_WLA<161> T_WLA<160> T_WLA<159> T_WLA<158> 
+ T_WLA<157> T_WLA<156> T_WLA<155> T_WLA<154> T_WLA<153> T_WLA<152> T_WLA<151> T_WLA<150> T_WLA<149> 
+ T_WLA<148> T_WLA<147> T_WLA<146> T_WLA<145> T_WLA<144> T_WLA<143> T_WLA<142> T_WLA<141> T_WLA<140> 
+ T_WLA<139> T_WLA<138> T_WLA<137> T_WLA<136> T_WLA<135> T_WLA<134> T_WLA<133> T_WLA<132> T_WLA<131> 
+ T_WLA<130> T_WLA<129> T_WLA<128> T_WLA<127> T_WLA<126> T_WLA<125> T_WLA<124> T_WLA<123> T_WLA<122> 
+ T_WLA<121> T_WLA<120> T_WLA<119> T_WLA<118> T_WLA<117> T_WLA<116> T_WLA<115> T_WLA<114> T_WLA<113> 
+ T_WLA<112> T_WLA<111> T_WLA<110> T_WLA<109> T_WLA<108> T_WLA<107> T_WLA<106> T_WLA<105> T_WLA<104> 
+ T_WLA<103> T_WLA<102> T_WLA<101> T_WLA<100> T_WLA<99> T_WLA<98> T_WLA<97> T_WLA<96> T_WLA<95> 
+ T_WLA<94> T_WLA<93> T_WLA<92> T_WLA<91> T_WLA<90> T_WLA<89> T_WLA<88> T_WLA<87> T_WLA<86> 
+ T_WLA<85> T_WLA<84> T_WLA<83> T_WLA<82> T_WLA<81> T_WLA<80> T_WLA<79> T_WLA<78> T_WLA<77> 
+ T_WLA<76> T_WLA<75> T_WLA<74> T_WLA<73> T_WLA<72> T_WLA<71> T_WLA<70> T_WLA<69> T_WLA<68> 
+ T_WLA<67> T_WLA<66> T_WLA<65> T_WLA<64> T_WLA<63> T_WLA<62> T_WLA<61> T_WLA<60> T_WLA<59> 
+ T_WLA<58> T_WLA<57> T_WLA<56> T_WLA<55> T_WLA<54> T_WLA<53> T_WLA<52> T_WLA<51> T_WLA<50> 
+ T_WLA<49> T_WLA<48> T_WLA<47> T_WLA<46> T_WLA<45> T_WLA<44> T_WLA<43> T_WLA<42> T_WLA<41> 
+ T_WLA<40> T_WLA<39> T_WLA<38> T_WLA<37> T_WLA<36> T_WLA<35> T_WLA<34> T_WLA<33> T_WLA<32> 
+ T_WLA<31> T_WLA<30> T_WLA<29> T_WLA<28> T_WLA<27> T_WLA<26> T_WLA<25> T_WLA<24> T_WLA<23> 
+ T_WLA<22> T_WLA<21> T_WLA<20> T_WLA<19> T_WLA<18> T_WLA<17> T_WLA<16> T_WLA<15> T_WLA<14> 
+ T_WLA<13> T_WLA<12> T_WLA<11> T_WLA<10> T_WLA<9> T_WLA<8> T_WLA<7> T_WLA<6> T_WLA<5> 
+ T_WLA<4> T_WLA<3> T_WLA<2> T_WLA<1> T_WLA<0> T_WLB<255> T_WLB<254> T_WLB<253> T_WLB<252> 
+ T_WLB<251> T_WLB<250> T_WLB<249> T_WLB<248> T_WLB<247> T_WLB<246> T_WLB<245> T_WLB<244> T_WLB<243> 
+ T_WLB<242> T_WLB<241> T_WLB<240> T_WLB<239> T_WLB<238> T_WLB<237> T_WLB<236> T_WLB<235> T_WLB<234> 
+ T_WLB<233> T_WLB<232> T_WLB<231> T_WLB<230> T_WLB<229> T_WLB<228> T_WLB<227> T_WLB<226> T_WLB<225> 
+ T_WLB<224> T_WLB<223> T_WLB<222> T_WLB<221> T_WLB<220> T_WLB<219> T_WLB<218> T_WLB<217> T_WLB<216> 
+ T_WLB<215> T_WLB<214> T_WLB<213> T_WLB<212> T_WLB<211> T_WLB<210> T_WLB<209> T_WLB<208> T_WLB<207> 
+ T_WLB<206> T_WLB<205> T_WLB<204> T_WLB<203> T_WLB<202> T_WLB<201> T_WLB<200> T_WLB<199> T_WLB<198> 
+ T_WLB<197> T_WLB<196> T_WLB<195> T_WLB<194> T_WLB<193> T_WLB<192> T_WLB<191> T_WLB<190> T_WLB<189> 
+ T_WLB<188> T_WLB<187> T_WLB<186> T_WLB<185> T_WLB<184> T_WLB<183> T_WLB<182> T_WLB<181> T_WLB<180> 
+ T_WLB<179> T_WLB<178> T_WLB<177> T_WLB<176> T_WLB<175> T_WLB<174> T_WLB<173> T_WLB<172> T_WLB<171> 
+ T_WLB<170> T_WLB<169> T_WLB<168> T_WLB<167> T_WLB<166> T_WLB<165> T_WLB<164> T_WLB<163> T_WLB<162> 
+ T_WLB<161> T_WLB<160> T_WLB<159> T_WLB<158> T_WLB<157> T_WLB<156> T_WLB<155> T_WLB<154> T_WLB<153> 
+ T_WLB<152> T_WLB<151> T_WLB<150> T_WLB<149> T_WLB<148> T_WLB<147> T_WLB<146> T_WLB<145> T_WLB<144> 
+ T_WLB<143> T_WLB<142> T_WLB<141> T_WLB<140> T_WLB<139> T_WLB<138> T_WLB<137> T_WLB<136> T_WLB<135> 
+ T_WLB<134> T_WLB<133> T_WLB<132> T_WLB<131> T_WLB<130> T_WLB<129> T_WLB<128> T_WLB<127> T_WLB<126> 
+ T_WLB<125> T_WLB<124> T_WLB<123> T_WLB<122> T_WLB<121> T_WLB<120> T_WLB<119> T_WLB<118> T_WLB<117> 
+ T_WLB<116> T_WLB<115> T_WLB<114> T_WLB<113> T_WLB<112> T_WLB<111> T_WLB<110> T_WLB<109> T_WLB<108> 
+ T_WLB<107> T_WLB<106> T_WLB<105> T_WLB<104> T_WLB<103> T_WLB<102> T_WLB<101> T_WLB<100> T_WLB<99> 
+ T_WLB<98> T_WLB<97> T_WLB<96> T_WLB<95> T_WLB<94> T_WLB<93> T_WLB<92> T_WLB<91> T_WLB<90> 
+ T_WLB<89> T_WLB<88> T_WLB<87> T_WLB<86> T_WLB<85> T_WLB<84> T_WLB<83> T_WLB<82> T_WLB<81> 
+ T_WLB<80> T_WLB<79> T_WLB<78> T_WLB<77> T_WLB<76> T_WLB<75> T_WLB<74> T_WLB<73> T_WLB<72> 
+ T_WLB<71> T_WLB<70> T_WLB<69> T_WLB<68> T_WLB<67> T_WLB<66> T_WLB<65> T_WLB<64> T_WLB<63> 
+ T_WLB<62> T_WLB<61> T_WLB<60> T_WLB<59> T_WLB<58> T_WLB<57> T_WLB<56> T_WLB<55> T_WLB<54> 
+ T_WLB<53> T_WLB<52> T_WLB<51> T_WLB<50> T_WLB<49> T_WLB<48> T_WLB<47> T_WLB<46> T_WLB<45> 
+ T_WLB<44> T_WLB<43> T_WLB<42> T_WLB<41> T_WLB<40> T_WLB<39> T_WLB<38> T_WLB<37> T_WLB<36> 
+ T_WLB<35> T_WLB<34> T_WLB<33> T_WLB<32> T_WLB<31> T_WLB<30> T_WLB<29> T_WLB<28> T_WLB<27> 
+ T_WLB<26> T_WLB<25> T_WLB<24> T_WLB<23> T_WLB<22> T_WLB<21> T_WLB<20> T_WLB<19> T_WLB<18> 
+ T_WLB<17> T_WLB<16> T_WLB<15> T_WLB<14> T_WLB<13> T_WLB<12> T_WLB<11> T_WLB<10> T_WLB<9> 
+ T_WLB<8> T_WLB<7> T_WLB<6> T_WLB<5> T_WLB<4> T_WLB<3> T_WLB<2> T_WLB<1> T_WLB<0> 
+  / dpram16x4096_AR_COLX8_ROWX256
XAR_BOT<5>
+ B_BLA<11> B_BLA<10> B_BLA_N<11> B_BLA_N<10> B_BLB<11> B_BLB<10> B_BLB_N<11> B_BLB_N<10> VSS 
+ VDD B_WLA<255> B_WLA<254> B_WLA<253> B_WLA<252> B_WLA<251> B_WLA<250> B_WLA<249> B_WLA<248> 
+ B_WLA<247> B_WLA<246> B_WLA<245> B_WLA<244> B_WLA<243> B_WLA<242> B_WLA<241> B_WLA<240> B_WLA<239> 
+ B_WLA<238> B_WLA<237> B_WLA<236> B_WLA<235> B_WLA<234> B_WLA<233> B_WLA<232> B_WLA<231> B_WLA<230> 
+ B_WLA<229> B_WLA<228> B_WLA<227> B_WLA<226> B_WLA<225> B_WLA<224> B_WLA<223> B_WLA<222> B_WLA<221> 
+ B_WLA<220> B_WLA<219> B_WLA<218> B_WLA<217> B_WLA<216> B_WLA<215> B_WLA<214> B_WLA<213> B_WLA<212> 
+ B_WLA<211> B_WLA<210> B_WLA<209> B_WLA<208> B_WLA<207> B_WLA<206> B_WLA<205> B_WLA<204> B_WLA<203> 
+ B_WLA<202> B_WLA<201> B_WLA<200> B_WLA<199> B_WLA<198> B_WLA<197> B_WLA<196> B_WLA<195> B_WLA<194> 
+ B_WLA<193> B_WLA<192> B_WLA<191> B_WLA<190> B_WLA<189> B_WLA<188> B_WLA<187> B_WLA<186> B_WLA<185> 
+ B_WLA<184> B_WLA<183> B_WLA<182> B_WLA<181> B_WLA<180> B_WLA<179> B_WLA<178> B_WLA<177> B_WLA<176> 
+ B_WLA<175> B_WLA<174> B_WLA<173> B_WLA<172> B_WLA<171> B_WLA<170> B_WLA<169> B_WLA<168> B_WLA<167> 
+ B_WLA<166> B_WLA<165> B_WLA<164> B_WLA<163> B_WLA<162> B_WLA<161> B_WLA<160> B_WLA<159> B_WLA<158> 
+ B_WLA<157> B_WLA<156> B_WLA<155> B_WLA<154> B_WLA<153> B_WLA<152> B_WLA<151> B_WLA<150> B_WLA<149> 
+ B_WLA<148> B_WLA<147> B_WLA<146> B_WLA<145> B_WLA<144> B_WLA<143> B_WLA<142> B_WLA<141> B_WLA<140> 
+ B_WLA<139> B_WLA<138> B_WLA<137> B_WLA<136> B_WLA<135> B_WLA<134> B_WLA<133> B_WLA<132> B_WLA<131> 
+ B_WLA<130> B_WLA<129> B_WLA<128> B_WLA<127> B_WLA<126> B_WLA<125> B_WLA<124> B_WLA<123> B_WLA<122> 
+ B_WLA<121> B_WLA<120> B_WLA<119> B_WLA<118> B_WLA<117> B_WLA<116> B_WLA<115> B_WLA<114> B_WLA<113> 
+ B_WLA<112> B_WLA<111> B_WLA<110> B_WLA<109> B_WLA<108> B_WLA<107> B_WLA<106> B_WLA<105> B_WLA<104> 
+ B_WLA<103> B_WLA<102> B_WLA<101> B_WLA<100> B_WLA<99> B_WLA<98> B_WLA<97> B_WLA<96> B_WLA<95> 
+ B_WLA<94> B_WLA<93> B_WLA<92> B_WLA<91> B_WLA<90> B_WLA<89> B_WLA<88> B_WLA<87> B_WLA<86> 
+ B_WLA<85> B_WLA<84> B_WLA<83> B_WLA<82> B_WLA<81> B_WLA<80> B_WLA<79> B_WLA<78> B_WLA<77> 
+ B_WLA<76> B_WLA<75> B_WLA<74> B_WLA<73> B_WLA<72> B_WLA<71> B_WLA<70> B_WLA<69> B_WLA<68> 
+ B_WLA<67> B_WLA<66> B_WLA<65> B_WLA<64> B_WLA<63> B_WLA<62> B_WLA<61> B_WLA<60> B_WLA<59> 
+ B_WLA<58> B_WLA<57> B_WLA<56> B_WLA<55> B_WLA<54> B_WLA<53> B_WLA<52> B_WLA<51> B_WLA<50> 
+ B_WLA<49> B_WLA<48> B_WLA<47> B_WLA<46> B_WLA<45> B_WLA<44> B_WLA<43> B_WLA<42> B_WLA<41> 
+ B_WLA<40> B_WLA<39> B_WLA<38> B_WLA<37> B_WLA<36> B_WLA<35> B_WLA<34> B_WLA<33> B_WLA<32> 
+ B_WLA<31> B_WLA<30> B_WLA<29> B_WLA<28> B_WLA<27> B_WLA<26> B_WLA<25> B_WLA<24> B_WLA<23> 
+ B_WLA<22> B_WLA<21> B_WLA<20> B_WLA<19> B_WLA<18> B_WLA<17> B_WLA<16> B_WLA<15> B_WLA<14> 
+ B_WLA<13> B_WLA<12> B_WLA<11> B_WLA<10> B_WLA<9> B_WLA<8> B_WLA<7> B_WLA<6> B_WLA<5> 
+ B_WLA<4> B_WLA<3> B_WLA<2> B_WLA<1> B_WLA<0> B_WLB<255> B_WLB<254> B_WLB<253> B_WLB<252> 
+ B_WLB<251> B_WLB<250> B_WLB<249> B_WLB<248> B_WLB<247> B_WLB<246> B_WLB<245> B_WLB<244> B_WLB<243> 
+ B_WLB<242> B_WLB<241> B_WLB<240> B_WLB<239> B_WLB<238> B_WLB<237> B_WLB<236> B_WLB<235> B_WLB<234> 
+ B_WLB<233> B_WLB<232> B_WLB<231> B_WLB<230> B_WLB<229> B_WLB<228> B_WLB<227> B_WLB<226> B_WLB<225> 
+ B_WLB<224> B_WLB<223> B_WLB<222> B_WLB<221> B_WLB<220> B_WLB<219> B_WLB<218> B_WLB<217> B_WLB<216> 
+ B_WLB<215> B_WLB<214> B_WLB<213> B_WLB<212> B_WLB<211> B_WLB<210> B_WLB<209> B_WLB<208> B_WLB<207> 
+ B_WLB<206> B_WLB<205> B_WLB<204> B_WLB<203> B_WLB<202> B_WLB<201> B_WLB<200> B_WLB<199> B_WLB<198> 
+ B_WLB<197> B_WLB<196> B_WLB<195> B_WLB<194> B_WLB<193> B_WLB<192> B_WLB<191> B_WLB<190> B_WLB<189> 
+ B_WLB<188> B_WLB<187> B_WLB<186> B_WLB<185> B_WLB<184> B_WLB<183> B_WLB<182> B_WLB<181> B_WLB<180> 
+ B_WLB<179> B_WLB<178> B_WLB<177> B_WLB<176> B_WLB<175> B_WLB<174> B_WLB<173> B_WLB<172> B_WLB<171> 
+ B_WLB<170> B_WLB<169> B_WLB<168> B_WLB<167> B_WLB<166> B_WLB<165> B_WLB<164> B_WLB<163> B_WLB<162> 
+ B_WLB<161> B_WLB<160> B_WLB<159> B_WLB<158> B_WLB<157> B_WLB<156> B_WLB<155> B_WLB<154> B_WLB<153> 
+ B_WLB<152> B_WLB<151> B_WLB<150> B_WLB<149> B_WLB<148> B_WLB<147> B_WLB<146> B_WLB<145> B_WLB<144> 
+ B_WLB<143> B_WLB<142> B_WLB<141> B_WLB<140> B_WLB<139> B_WLB<138> B_WLB<137> B_WLB<136> B_WLB<135> 
+ B_WLB<134> B_WLB<133> B_WLB<132> B_WLB<131> B_WLB<130> B_WLB<129> B_WLB<128> B_WLB<127> B_WLB<126> 
+ B_WLB<125> B_WLB<124> B_WLB<123> B_WLB<122> B_WLB<121> B_WLB<120> B_WLB<119> B_WLB<118> B_WLB<117> 
+ B_WLB<116> B_WLB<115> B_WLB<114> B_WLB<113> B_WLB<112> B_WLB<111> B_WLB<110> B_WLB<109> B_WLB<108> 
+ B_WLB<107> B_WLB<106> B_WLB<105> B_WLB<104> B_WLB<103> B_WLB<102> B_WLB<101> B_WLB<100> B_WLB<99> 
+ B_WLB<98> B_WLB<97> B_WLB<96> B_WLB<95> B_WLB<94> B_WLB<93> B_WLB<92> B_WLB<91> B_WLB<90> 
+ B_WLB<89> B_WLB<88> B_WLB<87> B_WLB<86> B_WLB<85> B_WLB<84> B_WLB<83> B_WLB<82> B_WLB<81> 
+ B_WLB<80> B_WLB<79> B_WLB<78> B_WLB<77> B_WLB<76> B_WLB<75> B_WLB<74> B_WLB<73> B_WLB<72> 
+ B_WLB<71> B_WLB<70> B_WLB<69> B_WLB<68> B_WLB<67> B_WLB<66> B_WLB<65> B_WLB<64> B_WLB<63> 
+ B_WLB<62> B_WLB<61> B_WLB<60> B_WLB<59> B_WLB<58> B_WLB<57> B_WLB<56> B_WLB<55> B_WLB<54> 
+ B_WLB<53> B_WLB<52> B_WLB<51> B_WLB<50> B_WLB<49> B_WLB<48> B_WLB<47> B_WLB<46> B_WLB<45> 
+ B_WLB<44> B_WLB<43> B_WLB<42> B_WLB<41> B_WLB<40> B_WLB<39> B_WLB<38> B_WLB<37> B_WLB<36> 
+ B_WLB<35> B_WLB<34> B_WLB<33> B_WLB<32> B_WLB<31> B_WLB<30> B_WLB<29> B_WLB<28> B_WLB<27> 
+ B_WLB<26> B_WLB<25> B_WLB<24> B_WLB<23> B_WLB<22> B_WLB<21> B_WLB<20> B_WLB<19> B_WLB<18> 
+ B_WLB<17> B_WLB<16> B_WLB<15> B_WLB<14> B_WLB<13> B_WLB<12> B_WLB<11> B_WLB<10> B_WLB<9> 
+ B_WLB<8> B_WLB<7> B_WLB<6> B_WLB<5> B_WLB<4> B_WLB<3> B_WLB<2> B_WLB<1> B_WLB<0> 
+  / dpram16x4096_AR_COLX8_ROWX256
XAR_TOP<4>
+ T_BLA<9> T_BLA<8> T_BLA_N<9> T_BLA_N<8> T_BLB<9> T_BLB<8> T_BLB_N<9> T_BLB_N<8> VSS 
+ VDD T_WLA<255> T_WLA<254> T_WLA<253> T_WLA<252> T_WLA<251> T_WLA<250> T_WLA<249> T_WLA<248> 
+ T_WLA<247> T_WLA<246> T_WLA<245> T_WLA<244> T_WLA<243> T_WLA<242> T_WLA<241> T_WLA<240> T_WLA<239> 
+ T_WLA<238> T_WLA<237> T_WLA<236> T_WLA<235> T_WLA<234> T_WLA<233> T_WLA<232> T_WLA<231> T_WLA<230> 
+ T_WLA<229> T_WLA<228> T_WLA<227> T_WLA<226> T_WLA<225> T_WLA<224> T_WLA<223> T_WLA<222> T_WLA<221> 
+ T_WLA<220> T_WLA<219> T_WLA<218> T_WLA<217> T_WLA<216> T_WLA<215> T_WLA<214> T_WLA<213> T_WLA<212> 
+ T_WLA<211> T_WLA<210> T_WLA<209> T_WLA<208> T_WLA<207> T_WLA<206> T_WLA<205> T_WLA<204> T_WLA<203> 
+ T_WLA<202> T_WLA<201> T_WLA<200> T_WLA<199> T_WLA<198> T_WLA<197> T_WLA<196> T_WLA<195> T_WLA<194> 
+ T_WLA<193> T_WLA<192> T_WLA<191> T_WLA<190> T_WLA<189> T_WLA<188> T_WLA<187> T_WLA<186> T_WLA<185> 
+ T_WLA<184> T_WLA<183> T_WLA<182> T_WLA<181> T_WLA<180> T_WLA<179> T_WLA<178> T_WLA<177> T_WLA<176> 
+ T_WLA<175> T_WLA<174> T_WLA<173> T_WLA<172> T_WLA<171> T_WLA<170> T_WLA<169> T_WLA<168> T_WLA<167> 
+ T_WLA<166> T_WLA<165> T_WLA<164> T_WLA<163> T_WLA<162> T_WLA<161> T_WLA<160> T_WLA<159> T_WLA<158> 
+ T_WLA<157> T_WLA<156> T_WLA<155> T_WLA<154> T_WLA<153> T_WLA<152> T_WLA<151> T_WLA<150> T_WLA<149> 
+ T_WLA<148> T_WLA<147> T_WLA<146> T_WLA<145> T_WLA<144> T_WLA<143> T_WLA<142> T_WLA<141> T_WLA<140> 
+ T_WLA<139> T_WLA<138> T_WLA<137> T_WLA<136> T_WLA<135> T_WLA<134> T_WLA<133> T_WLA<132> T_WLA<131> 
+ T_WLA<130> T_WLA<129> T_WLA<128> T_WLA<127> T_WLA<126> T_WLA<125> T_WLA<124> T_WLA<123> T_WLA<122> 
+ T_WLA<121> T_WLA<120> T_WLA<119> T_WLA<118> T_WLA<117> T_WLA<116> T_WLA<115> T_WLA<114> T_WLA<113> 
+ T_WLA<112> T_WLA<111> T_WLA<110> T_WLA<109> T_WLA<108> T_WLA<107> T_WLA<106> T_WLA<105> T_WLA<104> 
+ T_WLA<103> T_WLA<102> T_WLA<101> T_WLA<100> T_WLA<99> T_WLA<98> T_WLA<97> T_WLA<96> T_WLA<95> 
+ T_WLA<94> T_WLA<93> T_WLA<92> T_WLA<91> T_WLA<90> T_WLA<89> T_WLA<88> T_WLA<87> T_WLA<86> 
+ T_WLA<85> T_WLA<84> T_WLA<83> T_WLA<82> T_WLA<81> T_WLA<80> T_WLA<79> T_WLA<78> T_WLA<77> 
+ T_WLA<76> T_WLA<75> T_WLA<74> T_WLA<73> T_WLA<72> T_WLA<71> T_WLA<70> T_WLA<69> T_WLA<68> 
+ T_WLA<67> T_WLA<66> T_WLA<65> T_WLA<64> T_WLA<63> T_WLA<62> T_WLA<61> T_WLA<60> T_WLA<59> 
+ T_WLA<58> T_WLA<57> T_WLA<56> T_WLA<55> T_WLA<54> T_WLA<53> T_WLA<52> T_WLA<51> T_WLA<50> 
+ T_WLA<49> T_WLA<48> T_WLA<47> T_WLA<46> T_WLA<45> T_WLA<44> T_WLA<43> T_WLA<42> T_WLA<41> 
+ T_WLA<40> T_WLA<39> T_WLA<38> T_WLA<37> T_WLA<36> T_WLA<35> T_WLA<34> T_WLA<33> T_WLA<32> 
+ T_WLA<31> T_WLA<30> T_WLA<29> T_WLA<28> T_WLA<27> T_WLA<26> T_WLA<25> T_WLA<24> T_WLA<23> 
+ T_WLA<22> T_WLA<21> T_WLA<20> T_WLA<19> T_WLA<18> T_WLA<17> T_WLA<16> T_WLA<15> T_WLA<14> 
+ T_WLA<13> T_WLA<12> T_WLA<11> T_WLA<10> T_WLA<9> T_WLA<8> T_WLA<7> T_WLA<6> T_WLA<5> 
+ T_WLA<4> T_WLA<3> T_WLA<2> T_WLA<1> T_WLA<0> T_WLB<255> T_WLB<254> T_WLB<253> T_WLB<252> 
+ T_WLB<251> T_WLB<250> T_WLB<249> T_WLB<248> T_WLB<247> T_WLB<246> T_WLB<245> T_WLB<244> T_WLB<243> 
+ T_WLB<242> T_WLB<241> T_WLB<240> T_WLB<239> T_WLB<238> T_WLB<237> T_WLB<236> T_WLB<235> T_WLB<234> 
+ T_WLB<233> T_WLB<232> T_WLB<231> T_WLB<230> T_WLB<229> T_WLB<228> T_WLB<227> T_WLB<226> T_WLB<225> 
+ T_WLB<224> T_WLB<223> T_WLB<222> T_WLB<221> T_WLB<220> T_WLB<219> T_WLB<218> T_WLB<217> T_WLB<216> 
+ T_WLB<215> T_WLB<214> T_WLB<213> T_WLB<212> T_WLB<211> T_WLB<210> T_WLB<209> T_WLB<208> T_WLB<207> 
+ T_WLB<206> T_WLB<205> T_WLB<204> T_WLB<203> T_WLB<202> T_WLB<201> T_WLB<200> T_WLB<199> T_WLB<198> 
+ T_WLB<197> T_WLB<196> T_WLB<195> T_WLB<194> T_WLB<193> T_WLB<192> T_WLB<191> T_WLB<190> T_WLB<189> 
+ T_WLB<188> T_WLB<187> T_WLB<186> T_WLB<185> T_WLB<184> T_WLB<183> T_WLB<182> T_WLB<181> T_WLB<180> 
+ T_WLB<179> T_WLB<178> T_WLB<177> T_WLB<176> T_WLB<175> T_WLB<174> T_WLB<173> T_WLB<172> T_WLB<171> 
+ T_WLB<170> T_WLB<169> T_WLB<168> T_WLB<167> T_WLB<166> T_WLB<165> T_WLB<164> T_WLB<163> T_WLB<162> 
+ T_WLB<161> T_WLB<160> T_WLB<159> T_WLB<158> T_WLB<157> T_WLB<156> T_WLB<155> T_WLB<154> T_WLB<153> 
+ T_WLB<152> T_WLB<151> T_WLB<150> T_WLB<149> T_WLB<148> T_WLB<147> T_WLB<146> T_WLB<145> T_WLB<144> 
+ T_WLB<143> T_WLB<142> T_WLB<141> T_WLB<140> T_WLB<139> T_WLB<138> T_WLB<137> T_WLB<136> T_WLB<135> 
+ T_WLB<134> T_WLB<133> T_WLB<132> T_WLB<131> T_WLB<130> T_WLB<129> T_WLB<128> T_WLB<127> T_WLB<126> 
+ T_WLB<125> T_WLB<124> T_WLB<123> T_WLB<122> T_WLB<121> T_WLB<120> T_WLB<119> T_WLB<118> T_WLB<117> 
+ T_WLB<116> T_WLB<115> T_WLB<114> T_WLB<113> T_WLB<112> T_WLB<111> T_WLB<110> T_WLB<109> T_WLB<108> 
+ T_WLB<107> T_WLB<106> T_WLB<105> T_WLB<104> T_WLB<103> T_WLB<102> T_WLB<101> T_WLB<100> T_WLB<99> 
+ T_WLB<98> T_WLB<97> T_WLB<96> T_WLB<95> T_WLB<94> T_WLB<93> T_WLB<92> T_WLB<91> T_WLB<90> 
+ T_WLB<89> T_WLB<88> T_WLB<87> T_WLB<86> T_WLB<85> T_WLB<84> T_WLB<83> T_WLB<82> T_WLB<81> 
+ T_WLB<80> T_WLB<79> T_WLB<78> T_WLB<77> T_WLB<76> T_WLB<75> T_WLB<74> T_WLB<73> T_WLB<72> 
+ T_WLB<71> T_WLB<70> T_WLB<69> T_WLB<68> T_WLB<67> T_WLB<66> T_WLB<65> T_WLB<64> T_WLB<63> 
+ T_WLB<62> T_WLB<61> T_WLB<60> T_WLB<59> T_WLB<58> T_WLB<57> T_WLB<56> T_WLB<55> T_WLB<54> 
+ T_WLB<53> T_WLB<52> T_WLB<51> T_WLB<50> T_WLB<49> T_WLB<48> T_WLB<47> T_WLB<46> T_WLB<45> 
+ T_WLB<44> T_WLB<43> T_WLB<42> T_WLB<41> T_WLB<40> T_WLB<39> T_WLB<38> T_WLB<37> T_WLB<36> 
+ T_WLB<35> T_WLB<34> T_WLB<33> T_WLB<32> T_WLB<31> T_WLB<30> T_WLB<29> T_WLB<28> T_WLB<27> 
+ T_WLB<26> T_WLB<25> T_WLB<24> T_WLB<23> T_WLB<22> T_WLB<21> T_WLB<20> T_WLB<19> T_WLB<18> 
+ T_WLB<17> T_WLB<16> T_WLB<15> T_WLB<14> T_WLB<13> T_WLB<12> T_WLB<11> T_WLB<10> T_WLB<9> 
+ T_WLB<8> T_WLB<7> T_WLB<6> T_WLB<5> T_WLB<4> T_WLB<3> T_WLB<2> T_WLB<1> T_WLB<0> 
+  / dpram16x4096_AR_COLX8_ROWX256
XAR_BOT<4>
+ B_BLA<9> B_BLA<8> B_BLA_N<9> B_BLA_N<8> B_BLB<9> B_BLB<8> B_BLB_N<9> B_BLB_N<8> VSS 
+ VDD B_WLA<255> B_WLA<254> B_WLA<253> B_WLA<252> B_WLA<251> B_WLA<250> B_WLA<249> B_WLA<248> 
+ B_WLA<247> B_WLA<246> B_WLA<245> B_WLA<244> B_WLA<243> B_WLA<242> B_WLA<241> B_WLA<240> B_WLA<239> 
+ B_WLA<238> B_WLA<237> B_WLA<236> B_WLA<235> B_WLA<234> B_WLA<233> B_WLA<232> B_WLA<231> B_WLA<230> 
+ B_WLA<229> B_WLA<228> B_WLA<227> B_WLA<226> B_WLA<225> B_WLA<224> B_WLA<223> B_WLA<222> B_WLA<221> 
+ B_WLA<220> B_WLA<219> B_WLA<218> B_WLA<217> B_WLA<216> B_WLA<215> B_WLA<214> B_WLA<213> B_WLA<212> 
+ B_WLA<211> B_WLA<210> B_WLA<209> B_WLA<208> B_WLA<207> B_WLA<206> B_WLA<205> B_WLA<204> B_WLA<203> 
+ B_WLA<202> B_WLA<201> B_WLA<200> B_WLA<199> B_WLA<198> B_WLA<197> B_WLA<196> B_WLA<195> B_WLA<194> 
+ B_WLA<193> B_WLA<192> B_WLA<191> B_WLA<190> B_WLA<189> B_WLA<188> B_WLA<187> B_WLA<186> B_WLA<185> 
+ B_WLA<184> B_WLA<183> B_WLA<182> B_WLA<181> B_WLA<180> B_WLA<179> B_WLA<178> B_WLA<177> B_WLA<176> 
+ B_WLA<175> B_WLA<174> B_WLA<173> B_WLA<172> B_WLA<171> B_WLA<170> B_WLA<169> B_WLA<168> B_WLA<167> 
+ B_WLA<166> B_WLA<165> B_WLA<164> B_WLA<163> B_WLA<162> B_WLA<161> B_WLA<160> B_WLA<159> B_WLA<158> 
+ B_WLA<157> B_WLA<156> B_WLA<155> B_WLA<154> B_WLA<153> B_WLA<152> B_WLA<151> B_WLA<150> B_WLA<149> 
+ B_WLA<148> B_WLA<147> B_WLA<146> B_WLA<145> B_WLA<144> B_WLA<143> B_WLA<142> B_WLA<141> B_WLA<140> 
+ B_WLA<139> B_WLA<138> B_WLA<137> B_WLA<136> B_WLA<135> B_WLA<134> B_WLA<133> B_WLA<132> B_WLA<131> 
+ B_WLA<130> B_WLA<129> B_WLA<128> B_WLA<127> B_WLA<126> B_WLA<125> B_WLA<124> B_WLA<123> B_WLA<122> 
+ B_WLA<121> B_WLA<120> B_WLA<119> B_WLA<118> B_WLA<117> B_WLA<116> B_WLA<115> B_WLA<114> B_WLA<113> 
+ B_WLA<112> B_WLA<111> B_WLA<110> B_WLA<109> B_WLA<108> B_WLA<107> B_WLA<106> B_WLA<105> B_WLA<104> 
+ B_WLA<103> B_WLA<102> B_WLA<101> B_WLA<100> B_WLA<99> B_WLA<98> B_WLA<97> B_WLA<96> B_WLA<95> 
+ B_WLA<94> B_WLA<93> B_WLA<92> B_WLA<91> B_WLA<90> B_WLA<89> B_WLA<88> B_WLA<87> B_WLA<86> 
+ B_WLA<85> B_WLA<84> B_WLA<83> B_WLA<82> B_WLA<81> B_WLA<80> B_WLA<79> B_WLA<78> B_WLA<77> 
+ B_WLA<76> B_WLA<75> B_WLA<74> B_WLA<73> B_WLA<72> B_WLA<71> B_WLA<70> B_WLA<69> B_WLA<68> 
+ B_WLA<67> B_WLA<66> B_WLA<65> B_WLA<64> B_WLA<63> B_WLA<62> B_WLA<61> B_WLA<60> B_WLA<59> 
+ B_WLA<58> B_WLA<57> B_WLA<56> B_WLA<55> B_WLA<54> B_WLA<53> B_WLA<52> B_WLA<51> B_WLA<50> 
+ B_WLA<49> B_WLA<48> B_WLA<47> B_WLA<46> B_WLA<45> B_WLA<44> B_WLA<43> B_WLA<42> B_WLA<41> 
+ B_WLA<40> B_WLA<39> B_WLA<38> B_WLA<37> B_WLA<36> B_WLA<35> B_WLA<34> B_WLA<33> B_WLA<32> 
+ B_WLA<31> B_WLA<30> B_WLA<29> B_WLA<28> B_WLA<27> B_WLA<26> B_WLA<25> B_WLA<24> B_WLA<23> 
+ B_WLA<22> B_WLA<21> B_WLA<20> B_WLA<19> B_WLA<18> B_WLA<17> B_WLA<16> B_WLA<15> B_WLA<14> 
+ B_WLA<13> B_WLA<12> B_WLA<11> B_WLA<10> B_WLA<9> B_WLA<8> B_WLA<7> B_WLA<6> B_WLA<5> 
+ B_WLA<4> B_WLA<3> B_WLA<2> B_WLA<1> B_WLA<0> B_WLB<255> B_WLB<254> B_WLB<253> B_WLB<252> 
+ B_WLB<251> B_WLB<250> B_WLB<249> B_WLB<248> B_WLB<247> B_WLB<246> B_WLB<245> B_WLB<244> B_WLB<243> 
+ B_WLB<242> B_WLB<241> B_WLB<240> B_WLB<239> B_WLB<238> B_WLB<237> B_WLB<236> B_WLB<235> B_WLB<234> 
+ B_WLB<233> B_WLB<232> B_WLB<231> B_WLB<230> B_WLB<229> B_WLB<228> B_WLB<227> B_WLB<226> B_WLB<225> 
+ B_WLB<224> B_WLB<223> B_WLB<222> B_WLB<221> B_WLB<220> B_WLB<219> B_WLB<218> B_WLB<217> B_WLB<216> 
+ B_WLB<215> B_WLB<214> B_WLB<213> B_WLB<212> B_WLB<211> B_WLB<210> B_WLB<209> B_WLB<208> B_WLB<207> 
+ B_WLB<206> B_WLB<205> B_WLB<204> B_WLB<203> B_WLB<202> B_WLB<201> B_WLB<200> B_WLB<199> B_WLB<198> 
+ B_WLB<197> B_WLB<196> B_WLB<195> B_WLB<194> B_WLB<193> B_WLB<192> B_WLB<191> B_WLB<190> B_WLB<189> 
+ B_WLB<188> B_WLB<187> B_WLB<186> B_WLB<185> B_WLB<184> B_WLB<183> B_WLB<182> B_WLB<181> B_WLB<180> 
+ B_WLB<179> B_WLB<178> B_WLB<177> B_WLB<176> B_WLB<175> B_WLB<174> B_WLB<173> B_WLB<172> B_WLB<171> 
+ B_WLB<170> B_WLB<169> B_WLB<168> B_WLB<167> B_WLB<166> B_WLB<165> B_WLB<164> B_WLB<163> B_WLB<162> 
+ B_WLB<161> B_WLB<160> B_WLB<159> B_WLB<158> B_WLB<157> B_WLB<156> B_WLB<155> B_WLB<154> B_WLB<153> 
+ B_WLB<152> B_WLB<151> B_WLB<150> B_WLB<149> B_WLB<148> B_WLB<147> B_WLB<146> B_WLB<145> B_WLB<144> 
+ B_WLB<143> B_WLB<142> B_WLB<141> B_WLB<140> B_WLB<139> B_WLB<138> B_WLB<137> B_WLB<136> B_WLB<135> 
+ B_WLB<134> B_WLB<133> B_WLB<132> B_WLB<131> B_WLB<130> B_WLB<129> B_WLB<128> B_WLB<127> B_WLB<126> 
+ B_WLB<125> B_WLB<124> B_WLB<123> B_WLB<122> B_WLB<121> B_WLB<120> B_WLB<119> B_WLB<118> B_WLB<117> 
+ B_WLB<116> B_WLB<115> B_WLB<114> B_WLB<113> B_WLB<112> B_WLB<111> B_WLB<110> B_WLB<109> B_WLB<108> 
+ B_WLB<107> B_WLB<106> B_WLB<105> B_WLB<104> B_WLB<103> B_WLB<102> B_WLB<101> B_WLB<100> B_WLB<99> 
+ B_WLB<98> B_WLB<97> B_WLB<96> B_WLB<95> B_WLB<94> B_WLB<93> B_WLB<92> B_WLB<91> B_WLB<90> 
+ B_WLB<89> B_WLB<88> B_WLB<87> B_WLB<86> B_WLB<85> B_WLB<84> B_WLB<83> B_WLB<82> B_WLB<81> 
+ B_WLB<80> B_WLB<79> B_WLB<78> B_WLB<77> B_WLB<76> B_WLB<75> B_WLB<74> B_WLB<73> B_WLB<72> 
+ B_WLB<71> B_WLB<70> B_WLB<69> B_WLB<68> B_WLB<67> B_WLB<66> B_WLB<65> B_WLB<64> B_WLB<63> 
+ B_WLB<62> B_WLB<61> B_WLB<60> B_WLB<59> B_WLB<58> B_WLB<57> B_WLB<56> B_WLB<55> B_WLB<54> 
+ B_WLB<53> B_WLB<52> B_WLB<51> B_WLB<50> B_WLB<49> B_WLB<48> B_WLB<47> B_WLB<46> B_WLB<45> 
+ B_WLB<44> B_WLB<43> B_WLB<42> B_WLB<41> B_WLB<40> B_WLB<39> B_WLB<38> B_WLB<37> B_WLB<36> 
+ B_WLB<35> B_WLB<34> B_WLB<33> B_WLB<32> B_WLB<31> B_WLB<30> B_WLB<29> B_WLB<28> B_WLB<27> 
+ B_WLB<26> B_WLB<25> B_WLB<24> B_WLB<23> B_WLB<22> B_WLB<21> B_WLB<20> B_WLB<19> B_WLB<18> 
+ B_WLB<17> B_WLB<16> B_WLB<15> B_WLB<14> B_WLB<13> B_WLB<12> B_WLB<11> B_WLB<10> B_WLB<9> 
+ B_WLB<8> B_WLB<7> B_WLB<6> B_WLB<5> B_WLB<4> B_WLB<3> B_WLB<2> B_WLB<1> B_WLB<0> 
+  / dpram16x4096_AR_COLX8_ROWX256
XAR_TOP<3>
+ T_BLA<7> T_BLA<6> T_BLA_N<7> T_BLA_N<6> T_BLB<7> T_BLB<6> T_BLB_N<7> T_BLB_N<6> VSS 
+ VDD T_WLA<255> T_WLA<254> T_WLA<253> T_WLA<252> T_WLA<251> T_WLA<250> T_WLA<249> T_WLA<248> 
+ T_WLA<247> T_WLA<246> T_WLA<245> T_WLA<244> T_WLA<243> T_WLA<242> T_WLA<241> T_WLA<240> T_WLA<239> 
+ T_WLA<238> T_WLA<237> T_WLA<236> T_WLA<235> T_WLA<234> T_WLA<233> T_WLA<232> T_WLA<231> T_WLA<230> 
+ T_WLA<229> T_WLA<228> T_WLA<227> T_WLA<226> T_WLA<225> T_WLA<224> T_WLA<223> T_WLA<222> T_WLA<221> 
+ T_WLA<220> T_WLA<219> T_WLA<218> T_WLA<217> T_WLA<216> T_WLA<215> T_WLA<214> T_WLA<213> T_WLA<212> 
+ T_WLA<211> T_WLA<210> T_WLA<209> T_WLA<208> T_WLA<207> T_WLA<206> T_WLA<205> T_WLA<204> T_WLA<203> 
+ T_WLA<202> T_WLA<201> T_WLA<200> T_WLA<199> T_WLA<198> T_WLA<197> T_WLA<196> T_WLA<195> T_WLA<194> 
+ T_WLA<193> T_WLA<192> T_WLA<191> T_WLA<190> T_WLA<189> T_WLA<188> T_WLA<187> T_WLA<186> T_WLA<185> 
+ T_WLA<184> T_WLA<183> T_WLA<182> T_WLA<181> T_WLA<180> T_WLA<179> T_WLA<178> T_WLA<177> T_WLA<176> 
+ T_WLA<175> T_WLA<174> T_WLA<173> T_WLA<172> T_WLA<171> T_WLA<170> T_WLA<169> T_WLA<168> T_WLA<167> 
+ T_WLA<166> T_WLA<165> T_WLA<164> T_WLA<163> T_WLA<162> T_WLA<161> T_WLA<160> T_WLA<159> T_WLA<158> 
+ T_WLA<157> T_WLA<156> T_WLA<155> T_WLA<154> T_WLA<153> T_WLA<152> T_WLA<151> T_WLA<150> T_WLA<149> 
+ T_WLA<148> T_WLA<147> T_WLA<146> T_WLA<145> T_WLA<144> T_WLA<143> T_WLA<142> T_WLA<141> T_WLA<140> 
+ T_WLA<139> T_WLA<138> T_WLA<137> T_WLA<136> T_WLA<135> T_WLA<134> T_WLA<133> T_WLA<132> T_WLA<131> 
+ T_WLA<130> T_WLA<129> T_WLA<128> T_WLA<127> T_WLA<126> T_WLA<125> T_WLA<124> T_WLA<123> T_WLA<122> 
+ T_WLA<121> T_WLA<120> T_WLA<119> T_WLA<118> T_WLA<117> T_WLA<116> T_WLA<115> T_WLA<114> T_WLA<113> 
+ T_WLA<112> T_WLA<111> T_WLA<110> T_WLA<109> T_WLA<108> T_WLA<107> T_WLA<106> T_WLA<105> T_WLA<104> 
+ T_WLA<103> T_WLA<102> T_WLA<101> T_WLA<100> T_WLA<99> T_WLA<98> T_WLA<97> T_WLA<96> T_WLA<95> 
+ T_WLA<94> T_WLA<93> T_WLA<92> T_WLA<91> T_WLA<90> T_WLA<89> T_WLA<88> T_WLA<87> T_WLA<86> 
+ T_WLA<85> T_WLA<84> T_WLA<83> T_WLA<82> T_WLA<81> T_WLA<80> T_WLA<79> T_WLA<78> T_WLA<77> 
+ T_WLA<76> T_WLA<75> T_WLA<74> T_WLA<73> T_WLA<72> T_WLA<71> T_WLA<70> T_WLA<69> T_WLA<68> 
+ T_WLA<67> T_WLA<66> T_WLA<65> T_WLA<64> T_WLA<63> T_WLA<62> T_WLA<61> T_WLA<60> T_WLA<59> 
+ T_WLA<58> T_WLA<57> T_WLA<56> T_WLA<55> T_WLA<54> T_WLA<53> T_WLA<52> T_WLA<51> T_WLA<50> 
+ T_WLA<49> T_WLA<48> T_WLA<47> T_WLA<46> T_WLA<45> T_WLA<44> T_WLA<43> T_WLA<42> T_WLA<41> 
+ T_WLA<40> T_WLA<39> T_WLA<38> T_WLA<37> T_WLA<36> T_WLA<35> T_WLA<34> T_WLA<33> T_WLA<32> 
+ T_WLA<31> T_WLA<30> T_WLA<29> T_WLA<28> T_WLA<27> T_WLA<26> T_WLA<25> T_WLA<24> T_WLA<23> 
+ T_WLA<22> T_WLA<21> T_WLA<20> T_WLA<19> T_WLA<18> T_WLA<17> T_WLA<16> T_WLA<15> T_WLA<14> 
+ T_WLA<13> T_WLA<12> T_WLA<11> T_WLA<10> T_WLA<9> T_WLA<8> T_WLA<7> T_WLA<6> T_WLA<5> 
+ T_WLA<4> T_WLA<3> T_WLA<2> T_WLA<1> T_WLA<0> T_WLB<255> T_WLB<254> T_WLB<253> T_WLB<252> 
+ T_WLB<251> T_WLB<250> T_WLB<249> T_WLB<248> T_WLB<247> T_WLB<246> T_WLB<245> T_WLB<244> T_WLB<243> 
+ T_WLB<242> T_WLB<241> T_WLB<240> T_WLB<239> T_WLB<238> T_WLB<237> T_WLB<236> T_WLB<235> T_WLB<234> 
+ T_WLB<233> T_WLB<232> T_WLB<231> T_WLB<230> T_WLB<229> T_WLB<228> T_WLB<227> T_WLB<226> T_WLB<225> 
+ T_WLB<224> T_WLB<223> T_WLB<222> T_WLB<221> T_WLB<220> T_WLB<219> T_WLB<218> T_WLB<217> T_WLB<216> 
+ T_WLB<215> T_WLB<214> T_WLB<213> T_WLB<212> T_WLB<211> T_WLB<210> T_WLB<209> T_WLB<208> T_WLB<207> 
+ T_WLB<206> T_WLB<205> T_WLB<204> T_WLB<203> T_WLB<202> T_WLB<201> T_WLB<200> T_WLB<199> T_WLB<198> 
+ T_WLB<197> T_WLB<196> T_WLB<195> T_WLB<194> T_WLB<193> T_WLB<192> T_WLB<191> T_WLB<190> T_WLB<189> 
+ T_WLB<188> T_WLB<187> T_WLB<186> T_WLB<185> T_WLB<184> T_WLB<183> T_WLB<182> T_WLB<181> T_WLB<180> 
+ T_WLB<179> T_WLB<178> T_WLB<177> T_WLB<176> T_WLB<175> T_WLB<174> T_WLB<173> T_WLB<172> T_WLB<171> 
+ T_WLB<170> T_WLB<169> T_WLB<168> T_WLB<167> T_WLB<166> T_WLB<165> T_WLB<164> T_WLB<163> T_WLB<162> 
+ T_WLB<161> T_WLB<160> T_WLB<159> T_WLB<158> T_WLB<157> T_WLB<156> T_WLB<155> T_WLB<154> T_WLB<153> 
+ T_WLB<152> T_WLB<151> T_WLB<150> T_WLB<149> T_WLB<148> T_WLB<147> T_WLB<146> T_WLB<145> T_WLB<144> 
+ T_WLB<143> T_WLB<142> T_WLB<141> T_WLB<140> T_WLB<139> T_WLB<138> T_WLB<137> T_WLB<136> T_WLB<135> 
+ T_WLB<134> T_WLB<133> T_WLB<132> T_WLB<131> T_WLB<130> T_WLB<129> T_WLB<128> T_WLB<127> T_WLB<126> 
+ T_WLB<125> T_WLB<124> T_WLB<123> T_WLB<122> T_WLB<121> T_WLB<120> T_WLB<119> T_WLB<118> T_WLB<117> 
+ T_WLB<116> T_WLB<115> T_WLB<114> T_WLB<113> T_WLB<112> T_WLB<111> T_WLB<110> T_WLB<109> T_WLB<108> 
+ T_WLB<107> T_WLB<106> T_WLB<105> T_WLB<104> T_WLB<103> T_WLB<102> T_WLB<101> T_WLB<100> T_WLB<99> 
+ T_WLB<98> T_WLB<97> T_WLB<96> T_WLB<95> T_WLB<94> T_WLB<93> T_WLB<92> T_WLB<91> T_WLB<90> 
+ T_WLB<89> T_WLB<88> T_WLB<87> T_WLB<86> T_WLB<85> T_WLB<84> T_WLB<83> T_WLB<82> T_WLB<81> 
+ T_WLB<80> T_WLB<79> T_WLB<78> T_WLB<77> T_WLB<76> T_WLB<75> T_WLB<74> T_WLB<73> T_WLB<72> 
+ T_WLB<71> T_WLB<70> T_WLB<69> T_WLB<68> T_WLB<67> T_WLB<66> T_WLB<65> T_WLB<64> T_WLB<63> 
+ T_WLB<62> T_WLB<61> T_WLB<60> T_WLB<59> T_WLB<58> T_WLB<57> T_WLB<56> T_WLB<55> T_WLB<54> 
+ T_WLB<53> T_WLB<52> T_WLB<51> T_WLB<50> T_WLB<49> T_WLB<48> T_WLB<47> T_WLB<46> T_WLB<45> 
+ T_WLB<44> T_WLB<43> T_WLB<42> T_WLB<41> T_WLB<40> T_WLB<39> T_WLB<38> T_WLB<37> T_WLB<36> 
+ T_WLB<35> T_WLB<34> T_WLB<33> T_WLB<32> T_WLB<31> T_WLB<30> T_WLB<29> T_WLB<28> T_WLB<27> 
+ T_WLB<26> T_WLB<25> T_WLB<24> T_WLB<23> T_WLB<22> T_WLB<21> T_WLB<20> T_WLB<19> T_WLB<18> 
+ T_WLB<17> T_WLB<16> T_WLB<15> T_WLB<14> T_WLB<13> T_WLB<12> T_WLB<11> T_WLB<10> T_WLB<9> 
+ T_WLB<8> T_WLB<7> T_WLB<6> T_WLB<5> T_WLB<4> T_WLB<3> T_WLB<2> T_WLB<1> T_WLB<0> 
+  / dpram16x4096_AR_COLX8_ROWX256
XAR_BOT<3>
+ B_BLA<7> B_BLA<6> B_BLA_N<7> B_BLA_N<6> B_BLB<7> B_BLB<6> B_BLB_N<7> B_BLB_N<6> VSS 
+ VDD B_WLA<255> B_WLA<254> B_WLA<253> B_WLA<252> B_WLA<251> B_WLA<250> B_WLA<249> B_WLA<248> 
+ B_WLA<247> B_WLA<246> B_WLA<245> B_WLA<244> B_WLA<243> B_WLA<242> B_WLA<241> B_WLA<240> B_WLA<239> 
+ B_WLA<238> B_WLA<237> B_WLA<236> B_WLA<235> B_WLA<234> B_WLA<233> B_WLA<232> B_WLA<231> B_WLA<230> 
+ B_WLA<229> B_WLA<228> B_WLA<227> B_WLA<226> B_WLA<225> B_WLA<224> B_WLA<223> B_WLA<222> B_WLA<221> 
+ B_WLA<220> B_WLA<219> B_WLA<218> B_WLA<217> B_WLA<216> B_WLA<215> B_WLA<214> B_WLA<213> B_WLA<212> 
+ B_WLA<211> B_WLA<210> B_WLA<209> B_WLA<208> B_WLA<207> B_WLA<206> B_WLA<205> B_WLA<204> B_WLA<203> 
+ B_WLA<202> B_WLA<201> B_WLA<200> B_WLA<199> B_WLA<198> B_WLA<197> B_WLA<196> B_WLA<195> B_WLA<194> 
+ B_WLA<193> B_WLA<192> B_WLA<191> B_WLA<190> B_WLA<189> B_WLA<188> B_WLA<187> B_WLA<186> B_WLA<185> 
+ B_WLA<184> B_WLA<183> B_WLA<182> B_WLA<181> B_WLA<180> B_WLA<179> B_WLA<178> B_WLA<177> B_WLA<176> 
+ B_WLA<175> B_WLA<174> B_WLA<173> B_WLA<172> B_WLA<171> B_WLA<170> B_WLA<169> B_WLA<168> B_WLA<167> 
+ B_WLA<166> B_WLA<165> B_WLA<164> B_WLA<163> B_WLA<162> B_WLA<161> B_WLA<160> B_WLA<159> B_WLA<158> 
+ B_WLA<157> B_WLA<156> B_WLA<155> B_WLA<154> B_WLA<153> B_WLA<152> B_WLA<151> B_WLA<150> B_WLA<149> 
+ B_WLA<148> B_WLA<147> B_WLA<146> B_WLA<145> B_WLA<144> B_WLA<143> B_WLA<142> B_WLA<141> B_WLA<140> 
+ B_WLA<139> B_WLA<138> B_WLA<137> B_WLA<136> B_WLA<135> B_WLA<134> B_WLA<133> B_WLA<132> B_WLA<131> 
+ B_WLA<130> B_WLA<129> B_WLA<128> B_WLA<127> B_WLA<126> B_WLA<125> B_WLA<124> B_WLA<123> B_WLA<122> 
+ B_WLA<121> B_WLA<120> B_WLA<119> B_WLA<118> B_WLA<117> B_WLA<116> B_WLA<115> B_WLA<114> B_WLA<113> 
+ B_WLA<112> B_WLA<111> B_WLA<110> B_WLA<109> B_WLA<108> B_WLA<107> B_WLA<106> B_WLA<105> B_WLA<104> 
+ B_WLA<103> B_WLA<102> B_WLA<101> B_WLA<100> B_WLA<99> B_WLA<98> B_WLA<97> B_WLA<96> B_WLA<95> 
+ B_WLA<94> B_WLA<93> B_WLA<92> B_WLA<91> B_WLA<90> B_WLA<89> B_WLA<88> B_WLA<87> B_WLA<86> 
+ B_WLA<85> B_WLA<84> B_WLA<83> B_WLA<82> B_WLA<81> B_WLA<80> B_WLA<79> B_WLA<78> B_WLA<77> 
+ B_WLA<76> B_WLA<75> B_WLA<74> B_WLA<73> B_WLA<72> B_WLA<71> B_WLA<70> B_WLA<69> B_WLA<68> 
+ B_WLA<67> B_WLA<66> B_WLA<65> B_WLA<64> B_WLA<63> B_WLA<62> B_WLA<61> B_WLA<60> B_WLA<59> 
+ B_WLA<58> B_WLA<57> B_WLA<56> B_WLA<55> B_WLA<54> B_WLA<53> B_WLA<52> B_WLA<51> B_WLA<50> 
+ B_WLA<49> B_WLA<48> B_WLA<47> B_WLA<46> B_WLA<45> B_WLA<44> B_WLA<43> B_WLA<42> B_WLA<41> 
+ B_WLA<40> B_WLA<39> B_WLA<38> B_WLA<37> B_WLA<36> B_WLA<35> B_WLA<34> B_WLA<33> B_WLA<32> 
+ B_WLA<31> B_WLA<30> B_WLA<29> B_WLA<28> B_WLA<27> B_WLA<26> B_WLA<25> B_WLA<24> B_WLA<23> 
+ B_WLA<22> B_WLA<21> B_WLA<20> B_WLA<19> B_WLA<18> B_WLA<17> B_WLA<16> B_WLA<15> B_WLA<14> 
+ B_WLA<13> B_WLA<12> B_WLA<11> B_WLA<10> B_WLA<9> B_WLA<8> B_WLA<7> B_WLA<6> B_WLA<5> 
+ B_WLA<4> B_WLA<3> B_WLA<2> B_WLA<1> B_WLA<0> B_WLB<255> B_WLB<254> B_WLB<253> B_WLB<252> 
+ B_WLB<251> B_WLB<250> B_WLB<249> B_WLB<248> B_WLB<247> B_WLB<246> B_WLB<245> B_WLB<244> B_WLB<243> 
+ B_WLB<242> B_WLB<241> B_WLB<240> B_WLB<239> B_WLB<238> B_WLB<237> B_WLB<236> B_WLB<235> B_WLB<234> 
+ B_WLB<233> B_WLB<232> B_WLB<231> B_WLB<230> B_WLB<229> B_WLB<228> B_WLB<227> B_WLB<226> B_WLB<225> 
+ B_WLB<224> B_WLB<223> B_WLB<222> B_WLB<221> B_WLB<220> B_WLB<219> B_WLB<218> B_WLB<217> B_WLB<216> 
+ B_WLB<215> B_WLB<214> B_WLB<213> B_WLB<212> B_WLB<211> B_WLB<210> B_WLB<209> B_WLB<208> B_WLB<207> 
+ B_WLB<206> B_WLB<205> B_WLB<204> B_WLB<203> B_WLB<202> B_WLB<201> B_WLB<200> B_WLB<199> B_WLB<198> 
+ B_WLB<197> B_WLB<196> B_WLB<195> B_WLB<194> B_WLB<193> B_WLB<192> B_WLB<191> B_WLB<190> B_WLB<189> 
+ B_WLB<188> B_WLB<187> B_WLB<186> B_WLB<185> B_WLB<184> B_WLB<183> B_WLB<182> B_WLB<181> B_WLB<180> 
+ B_WLB<179> B_WLB<178> B_WLB<177> B_WLB<176> B_WLB<175> B_WLB<174> B_WLB<173> B_WLB<172> B_WLB<171> 
+ B_WLB<170> B_WLB<169> B_WLB<168> B_WLB<167> B_WLB<166> B_WLB<165> B_WLB<164> B_WLB<163> B_WLB<162> 
+ B_WLB<161> B_WLB<160> B_WLB<159> B_WLB<158> B_WLB<157> B_WLB<156> B_WLB<155> B_WLB<154> B_WLB<153> 
+ B_WLB<152> B_WLB<151> B_WLB<150> B_WLB<149> B_WLB<148> B_WLB<147> B_WLB<146> B_WLB<145> B_WLB<144> 
+ B_WLB<143> B_WLB<142> B_WLB<141> B_WLB<140> B_WLB<139> B_WLB<138> B_WLB<137> B_WLB<136> B_WLB<135> 
+ B_WLB<134> B_WLB<133> B_WLB<132> B_WLB<131> B_WLB<130> B_WLB<129> B_WLB<128> B_WLB<127> B_WLB<126> 
+ B_WLB<125> B_WLB<124> B_WLB<123> B_WLB<122> B_WLB<121> B_WLB<120> B_WLB<119> B_WLB<118> B_WLB<117> 
+ B_WLB<116> B_WLB<115> B_WLB<114> B_WLB<113> B_WLB<112> B_WLB<111> B_WLB<110> B_WLB<109> B_WLB<108> 
+ B_WLB<107> B_WLB<106> B_WLB<105> B_WLB<104> B_WLB<103> B_WLB<102> B_WLB<101> B_WLB<100> B_WLB<99> 
+ B_WLB<98> B_WLB<97> B_WLB<96> B_WLB<95> B_WLB<94> B_WLB<93> B_WLB<92> B_WLB<91> B_WLB<90> 
+ B_WLB<89> B_WLB<88> B_WLB<87> B_WLB<86> B_WLB<85> B_WLB<84> B_WLB<83> B_WLB<82> B_WLB<81> 
+ B_WLB<80> B_WLB<79> B_WLB<78> B_WLB<77> B_WLB<76> B_WLB<75> B_WLB<74> B_WLB<73> B_WLB<72> 
+ B_WLB<71> B_WLB<70> B_WLB<69> B_WLB<68> B_WLB<67> B_WLB<66> B_WLB<65> B_WLB<64> B_WLB<63> 
+ B_WLB<62> B_WLB<61> B_WLB<60> B_WLB<59> B_WLB<58> B_WLB<57> B_WLB<56> B_WLB<55> B_WLB<54> 
+ B_WLB<53> B_WLB<52> B_WLB<51> B_WLB<50> B_WLB<49> B_WLB<48> B_WLB<47> B_WLB<46> B_WLB<45> 
+ B_WLB<44> B_WLB<43> B_WLB<42> B_WLB<41> B_WLB<40> B_WLB<39> B_WLB<38> B_WLB<37> B_WLB<36> 
+ B_WLB<35> B_WLB<34> B_WLB<33> B_WLB<32> B_WLB<31> B_WLB<30> B_WLB<29> B_WLB<28> B_WLB<27> 
+ B_WLB<26> B_WLB<25> B_WLB<24> B_WLB<23> B_WLB<22> B_WLB<21> B_WLB<20> B_WLB<19> B_WLB<18> 
+ B_WLB<17> B_WLB<16> B_WLB<15> B_WLB<14> B_WLB<13> B_WLB<12> B_WLB<11> B_WLB<10> B_WLB<9> 
+ B_WLB<8> B_WLB<7> B_WLB<6> B_WLB<5> B_WLB<4> B_WLB<3> B_WLB<2> B_WLB<1> B_WLB<0> 
+  / dpram16x4096_AR_COLX8_ROWX256
XAR_TOP<2>
+ T_BLA<5> T_BLA<4> T_BLA_N<5> T_BLA_N<4> T_BLB<5> T_BLB<4> T_BLB_N<5> T_BLB_N<4> VSS 
+ VDD T_WLA<255> T_WLA<254> T_WLA<253> T_WLA<252> T_WLA<251> T_WLA<250> T_WLA<249> T_WLA<248> 
+ T_WLA<247> T_WLA<246> T_WLA<245> T_WLA<244> T_WLA<243> T_WLA<242> T_WLA<241> T_WLA<240> T_WLA<239> 
+ T_WLA<238> T_WLA<237> T_WLA<236> T_WLA<235> T_WLA<234> T_WLA<233> T_WLA<232> T_WLA<231> T_WLA<230> 
+ T_WLA<229> T_WLA<228> T_WLA<227> T_WLA<226> T_WLA<225> T_WLA<224> T_WLA<223> T_WLA<222> T_WLA<221> 
+ T_WLA<220> T_WLA<219> T_WLA<218> T_WLA<217> T_WLA<216> T_WLA<215> T_WLA<214> T_WLA<213> T_WLA<212> 
+ T_WLA<211> T_WLA<210> T_WLA<209> T_WLA<208> T_WLA<207> T_WLA<206> T_WLA<205> T_WLA<204> T_WLA<203> 
+ T_WLA<202> T_WLA<201> T_WLA<200> T_WLA<199> T_WLA<198> T_WLA<197> T_WLA<196> T_WLA<195> T_WLA<194> 
+ T_WLA<193> T_WLA<192> T_WLA<191> T_WLA<190> T_WLA<189> T_WLA<188> T_WLA<187> T_WLA<186> T_WLA<185> 
+ T_WLA<184> T_WLA<183> T_WLA<182> T_WLA<181> T_WLA<180> T_WLA<179> T_WLA<178> T_WLA<177> T_WLA<176> 
+ T_WLA<175> T_WLA<174> T_WLA<173> T_WLA<172> T_WLA<171> T_WLA<170> T_WLA<169> T_WLA<168> T_WLA<167> 
+ T_WLA<166> T_WLA<165> T_WLA<164> T_WLA<163> T_WLA<162> T_WLA<161> T_WLA<160> T_WLA<159> T_WLA<158> 
+ T_WLA<157> T_WLA<156> T_WLA<155> T_WLA<154> T_WLA<153> T_WLA<152> T_WLA<151> T_WLA<150> T_WLA<149> 
+ T_WLA<148> T_WLA<147> T_WLA<146> T_WLA<145> T_WLA<144> T_WLA<143> T_WLA<142> T_WLA<141> T_WLA<140> 
+ T_WLA<139> T_WLA<138> T_WLA<137> T_WLA<136> T_WLA<135> T_WLA<134> T_WLA<133> T_WLA<132> T_WLA<131> 
+ T_WLA<130> T_WLA<129> T_WLA<128> T_WLA<127> T_WLA<126> T_WLA<125> T_WLA<124> T_WLA<123> T_WLA<122> 
+ T_WLA<121> T_WLA<120> T_WLA<119> T_WLA<118> T_WLA<117> T_WLA<116> T_WLA<115> T_WLA<114> T_WLA<113> 
+ T_WLA<112> T_WLA<111> T_WLA<110> T_WLA<109> T_WLA<108> T_WLA<107> T_WLA<106> T_WLA<105> T_WLA<104> 
+ T_WLA<103> T_WLA<102> T_WLA<101> T_WLA<100> T_WLA<99> T_WLA<98> T_WLA<97> T_WLA<96> T_WLA<95> 
+ T_WLA<94> T_WLA<93> T_WLA<92> T_WLA<91> T_WLA<90> T_WLA<89> T_WLA<88> T_WLA<87> T_WLA<86> 
+ T_WLA<85> T_WLA<84> T_WLA<83> T_WLA<82> T_WLA<81> T_WLA<80> T_WLA<79> T_WLA<78> T_WLA<77> 
+ T_WLA<76> T_WLA<75> T_WLA<74> T_WLA<73> T_WLA<72> T_WLA<71> T_WLA<70> T_WLA<69> T_WLA<68> 
+ T_WLA<67> T_WLA<66> T_WLA<65> T_WLA<64> T_WLA<63> T_WLA<62> T_WLA<61> T_WLA<60> T_WLA<59> 
+ T_WLA<58> T_WLA<57> T_WLA<56> T_WLA<55> T_WLA<54> T_WLA<53> T_WLA<52> T_WLA<51> T_WLA<50> 
+ T_WLA<49> T_WLA<48> T_WLA<47> T_WLA<46> T_WLA<45> T_WLA<44> T_WLA<43> T_WLA<42> T_WLA<41> 
+ T_WLA<40> T_WLA<39> T_WLA<38> T_WLA<37> T_WLA<36> T_WLA<35> T_WLA<34> T_WLA<33> T_WLA<32> 
+ T_WLA<31> T_WLA<30> T_WLA<29> T_WLA<28> T_WLA<27> T_WLA<26> T_WLA<25> T_WLA<24> T_WLA<23> 
+ T_WLA<22> T_WLA<21> T_WLA<20> T_WLA<19> T_WLA<18> T_WLA<17> T_WLA<16> T_WLA<15> T_WLA<14> 
+ T_WLA<13> T_WLA<12> T_WLA<11> T_WLA<10> T_WLA<9> T_WLA<8> T_WLA<7> T_WLA<6> T_WLA<5> 
+ T_WLA<4> T_WLA<3> T_WLA<2> T_WLA<1> T_WLA<0> T_WLB<255> T_WLB<254> T_WLB<253> T_WLB<252> 
+ T_WLB<251> T_WLB<250> T_WLB<249> T_WLB<248> T_WLB<247> T_WLB<246> T_WLB<245> T_WLB<244> T_WLB<243> 
+ T_WLB<242> T_WLB<241> T_WLB<240> T_WLB<239> T_WLB<238> T_WLB<237> T_WLB<236> T_WLB<235> T_WLB<234> 
+ T_WLB<233> T_WLB<232> T_WLB<231> T_WLB<230> T_WLB<229> T_WLB<228> T_WLB<227> T_WLB<226> T_WLB<225> 
+ T_WLB<224> T_WLB<223> T_WLB<222> T_WLB<221> T_WLB<220> T_WLB<219> T_WLB<218> T_WLB<217> T_WLB<216> 
+ T_WLB<215> T_WLB<214> T_WLB<213> T_WLB<212> T_WLB<211> T_WLB<210> T_WLB<209> T_WLB<208> T_WLB<207> 
+ T_WLB<206> T_WLB<205> T_WLB<204> T_WLB<203> T_WLB<202> T_WLB<201> T_WLB<200> T_WLB<199> T_WLB<198> 
+ T_WLB<197> T_WLB<196> T_WLB<195> T_WLB<194> T_WLB<193> T_WLB<192> T_WLB<191> T_WLB<190> T_WLB<189> 
+ T_WLB<188> T_WLB<187> T_WLB<186> T_WLB<185> T_WLB<184> T_WLB<183> T_WLB<182> T_WLB<181> T_WLB<180> 
+ T_WLB<179> T_WLB<178> T_WLB<177> T_WLB<176> T_WLB<175> T_WLB<174> T_WLB<173> T_WLB<172> T_WLB<171> 
+ T_WLB<170> T_WLB<169> T_WLB<168> T_WLB<167> T_WLB<166> T_WLB<165> T_WLB<164> T_WLB<163> T_WLB<162> 
+ T_WLB<161> T_WLB<160> T_WLB<159> T_WLB<158> T_WLB<157> T_WLB<156> T_WLB<155> T_WLB<154> T_WLB<153> 
+ T_WLB<152> T_WLB<151> T_WLB<150> T_WLB<149> T_WLB<148> T_WLB<147> T_WLB<146> T_WLB<145> T_WLB<144> 
+ T_WLB<143> T_WLB<142> T_WLB<141> T_WLB<140> T_WLB<139> T_WLB<138> T_WLB<137> T_WLB<136> T_WLB<135> 
+ T_WLB<134> T_WLB<133> T_WLB<132> T_WLB<131> T_WLB<130> T_WLB<129> T_WLB<128> T_WLB<127> T_WLB<126> 
+ T_WLB<125> T_WLB<124> T_WLB<123> T_WLB<122> T_WLB<121> T_WLB<120> T_WLB<119> T_WLB<118> T_WLB<117> 
+ T_WLB<116> T_WLB<115> T_WLB<114> T_WLB<113> T_WLB<112> T_WLB<111> T_WLB<110> T_WLB<109> T_WLB<108> 
+ T_WLB<107> T_WLB<106> T_WLB<105> T_WLB<104> T_WLB<103> T_WLB<102> T_WLB<101> T_WLB<100> T_WLB<99> 
+ T_WLB<98> T_WLB<97> T_WLB<96> T_WLB<95> T_WLB<94> T_WLB<93> T_WLB<92> T_WLB<91> T_WLB<90> 
+ T_WLB<89> T_WLB<88> T_WLB<87> T_WLB<86> T_WLB<85> T_WLB<84> T_WLB<83> T_WLB<82> T_WLB<81> 
+ T_WLB<80> T_WLB<79> T_WLB<78> T_WLB<77> T_WLB<76> T_WLB<75> T_WLB<74> T_WLB<73> T_WLB<72> 
+ T_WLB<71> T_WLB<70> T_WLB<69> T_WLB<68> T_WLB<67> T_WLB<66> T_WLB<65> T_WLB<64> T_WLB<63> 
+ T_WLB<62> T_WLB<61> T_WLB<60> T_WLB<59> T_WLB<58> T_WLB<57> T_WLB<56> T_WLB<55> T_WLB<54> 
+ T_WLB<53> T_WLB<52> T_WLB<51> T_WLB<50> T_WLB<49> T_WLB<48> T_WLB<47> T_WLB<46> T_WLB<45> 
+ T_WLB<44> T_WLB<43> T_WLB<42> T_WLB<41> T_WLB<40> T_WLB<39> T_WLB<38> T_WLB<37> T_WLB<36> 
+ T_WLB<35> T_WLB<34> T_WLB<33> T_WLB<32> T_WLB<31> T_WLB<30> T_WLB<29> T_WLB<28> T_WLB<27> 
+ T_WLB<26> T_WLB<25> T_WLB<24> T_WLB<23> T_WLB<22> T_WLB<21> T_WLB<20> T_WLB<19> T_WLB<18> 
+ T_WLB<17> T_WLB<16> T_WLB<15> T_WLB<14> T_WLB<13> T_WLB<12> T_WLB<11> T_WLB<10> T_WLB<9> 
+ T_WLB<8> T_WLB<7> T_WLB<6> T_WLB<5> T_WLB<4> T_WLB<3> T_WLB<2> T_WLB<1> T_WLB<0> 
+  / dpram16x4096_AR_COLX8_ROWX256
XAR_BOT<2>
+ B_BLA<5> B_BLA<4> B_BLA_N<5> B_BLA_N<4> B_BLB<5> B_BLB<4> B_BLB_N<5> B_BLB_N<4> VSS 
+ VDD B_WLA<255> B_WLA<254> B_WLA<253> B_WLA<252> B_WLA<251> B_WLA<250> B_WLA<249> B_WLA<248> 
+ B_WLA<247> B_WLA<246> B_WLA<245> B_WLA<244> B_WLA<243> B_WLA<242> B_WLA<241> B_WLA<240> B_WLA<239> 
+ B_WLA<238> B_WLA<237> B_WLA<236> B_WLA<235> B_WLA<234> B_WLA<233> B_WLA<232> B_WLA<231> B_WLA<230> 
+ B_WLA<229> B_WLA<228> B_WLA<227> B_WLA<226> B_WLA<225> B_WLA<224> B_WLA<223> B_WLA<222> B_WLA<221> 
+ B_WLA<220> B_WLA<219> B_WLA<218> B_WLA<217> B_WLA<216> B_WLA<215> B_WLA<214> B_WLA<213> B_WLA<212> 
+ B_WLA<211> B_WLA<210> B_WLA<209> B_WLA<208> B_WLA<207> B_WLA<206> B_WLA<205> B_WLA<204> B_WLA<203> 
+ B_WLA<202> B_WLA<201> B_WLA<200> B_WLA<199> B_WLA<198> B_WLA<197> B_WLA<196> B_WLA<195> B_WLA<194> 
+ B_WLA<193> B_WLA<192> B_WLA<191> B_WLA<190> B_WLA<189> B_WLA<188> B_WLA<187> B_WLA<186> B_WLA<185> 
+ B_WLA<184> B_WLA<183> B_WLA<182> B_WLA<181> B_WLA<180> B_WLA<179> B_WLA<178> B_WLA<177> B_WLA<176> 
+ B_WLA<175> B_WLA<174> B_WLA<173> B_WLA<172> B_WLA<171> B_WLA<170> B_WLA<169> B_WLA<168> B_WLA<167> 
+ B_WLA<166> B_WLA<165> B_WLA<164> B_WLA<163> B_WLA<162> B_WLA<161> B_WLA<160> B_WLA<159> B_WLA<158> 
+ B_WLA<157> B_WLA<156> B_WLA<155> B_WLA<154> B_WLA<153> B_WLA<152> B_WLA<151> B_WLA<150> B_WLA<149> 
+ B_WLA<148> B_WLA<147> B_WLA<146> B_WLA<145> B_WLA<144> B_WLA<143> B_WLA<142> B_WLA<141> B_WLA<140> 
+ B_WLA<139> B_WLA<138> B_WLA<137> B_WLA<136> B_WLA<135> B_WLA<134> B_WLA<133> B_WLA<132> B_WLA<131> 
+ B_WLA<130> B_WLA<129> B_WLA<128> B_WLA<127> B_WLA<126> B_WLA<125> B_WLA<124> B_WLA<123> B_WLA<122> 
+ B_WLA<121> B_WLA<120> B_WLA<119> B_WLA<118> B_WLA<117> B_WLA<116> B_WLA<115> B_WLA<114> B_WLA<113> 
+ B_WLA<112> B_WLA<111> B_WLA<110> B_WLA<109> B_WLA<108> B_WLA<107> B_WLA<106> B_WLA<105> B_WLA<104> 
+ B_WLA<103> B_WLA<102> B_WLA<101> B_WLA<100> B_WLA<99> B_WLA<98> B_WLA<97> B_WLA<96> B_WLA<95> 
+ B_WLA<94> B_WLA<93> B_WLA<92> B_WLA<91> B_WLA<90> B_WLA<89> B_WLA<88> B_WLA<87> B_WLA<86> 
+ B_WLA<85> B_WLA<84> B_WLA<83> B_WLA<82> B_WLA<81> B_WLA<80> B_WLA<79> B_WLA<78> B_WLA<77> 
+ B_WLA<76> B_WLA<75> B_WLA<74> B_WLA<73> B_WLA<72> B_WLA<71> B_WLA<70> B_WLA<69> B_WLA<68> 
+ B_WLA<67> B_WLA<66> B_WLA<65> B_WLA<64> B_WLA<63> B_WLA<62> B_WLA<61> B_WLA<60> B_WLA<59> 
+ B_WLA<58> B_WLA<57> B_WLA<56> B_WLA<55> B_WLA<54> B_WLA<53> B_WLA<52> B_WLA<51> B_WLA<50> 
+ B_WLA<49> B_WLA<48> B_WLA<47> B_WLA<46> B_WLA<45> B_WLA<44> B_WLA<43> B_WLA<42> B_WLA<41> 
+ B_WLA<40> B_WLA<39> B_WLA<38> B_WLA<37> B_WLA<36> B_WLA<35> B_WLA<34> B_WLA<33> B_WLA<32> 
+ B_WLA<31> B_WLA<30> B_WLA<29> B_WLA<28> B_WLA<27> B_WLA<26> B_WLA<25> B_WLA<24> B_WLA<23> 
+ B_WLA<22> B_WLA<21> B_WLA<20> B_WLA<19> B_WLA<18> B_WLA<17> B_WLA<16> B_WLA<15> B_WLA<14> 
+ B_WLA<13> B_WLA<12> B_WLA<11> B_WLA<10> B_WLA<9> B_WLA<8> B_WLA<7> B_WLA<6> B_WLA<5> 
+ B_WLA<4> B_WLA<3> B_WLA<2> B_WLA<1> B_WLA<0> B_WLB<255> B_WLB<254> B_WLB<253> B_WLB<252> 
+ B_WLB<251> B_WLB<250> B_WLB<249> B_WLB<248> B_WLB<247> B_WLB<246> B_WLB<245> B_WLB<244> B_WLB<243> 
+ B_WLB<242> B_WLB<241> B_WLB<240> B_WLB<239> B_WLB<238> B_WLB<237> B_WLB<236> B_WLB<235> B_WLB<234> 
+ B_WLB<233> B_WLB<232> B_WLB<231> B_WLB<230> B_WLB<229> B_WLB<228> B_WLB<227> B_WLB<226> B_WLB<225> 
+ B_WLB<224> B_WLB<223> B_WLB<222> B_WLB<221> B_WLB<220> B_WLB<219> B_WLB<218> B_WLB<217> B_WLB<216> 
+ B_WLB<215> B_WLB<214> B_WLB<213> B_WLB<212> B_WLB<211> B_WLB<210> B_WLB<209> B_WLB<208> B_WLB<207> 
+ B_WLB<206> B_WLB<205> B_WLB<204> B_WLB<203> B_WLB<202> B_WLB<201> B_WLB<200> B_WLB<199> B_WLB<198> 
+ B_WLB<197> B_WLB<196> B_WLB<195> B_WLB<194> B_WLB<193> B_WLB<192> B_WLB<191> B_WLB<190> B_WLB<189> 
+ B_WLB<188> B_WLB<187> B_WLB<186> B_WLB<185> B_WLB<184> B_WLB<183> B_WLB<182> B_WLB<181> B_WLB<180> 
+ B_WLB<179> B_WLB<178> B_WLB<177> B_WLB<176> B_WLB<175> B_WLB<174> B_WLB<173> B_WLB<172> B_WLB<171> 
+ B_WLB<170> B_WLB<169> B_WLB<168> B_WLB<167> B_WLB<166> B_WLB<165> B_WLB<164> B_WLB<163> B_WLB<162> 
+ B_WLB<161> B_WLB<160> B_WLB<159> B_WLB<158> B_WLB<157> B_WLB<156> B_WLB<155> B_WLB<154> B_WLB<153> 
+ B_WLB<152> B_WLB<151> B_WLB<150> B_WLB<149> B_WLB<148> B_WLB<147> B_WLB<146> B_WLB<145> B_WLB<144> 
+ B_WLB<143> B_WLB<142> B_WLB<141> B_WLB<140> B_WLB<139> B_WLB<138> B_WLB<137> B_WLB<136> B_WLB<135> 
+ B_WLB<134> B_WLB<133> B_WLB<132> B_WLB<131> B_WLB<130> B_WLB<129> B_WLB<128> B_WLB<127> B_WLB<126> 
+ B_WLB<125> B_WLB<124> B_WLB<123> B_WLB<122> B_WLB<121> B_WLB<120> B_WLB<119> B_WLB<118> B_WLB<117> 
+ B_WLB<116> B_WLB<115> B_WLB<114> B_WLB<113> B_WLB<112> B_WLB<111> B_WLB<110> B_WLB<109> B_WLB<108> 
+ B_WLB<107> B_WLB<106> B_WLB<105> B_WLB<104> B_WLB<103> B_WLB<102> B_WLB<101> B_WLB<100> B_WLB<99> 
+ B_WLB<98> B_WLB<97> B_WLB<96> B_WLB<95> B_WLB<94> B_WLB<93> B_WLB<92> B_WLB<91> B_WLB<90> 
+ B_WLB<89> B_WLB<88> B_WLB<87> B_WLB<86> B_WLB<85> B_WLB<84> B_WLB<83> B_WLB<82> B_WLB<81> 
+ B_WLB<80> B_WLB<79> B_WLB<78> B_WLB<77> B_WLB<76> B_WLB<75> B_WLB<74> B_WLB<73> B_WLB<72> 
+ B_WLB<71> B_WLB<70> B_WLB<69> B_WLB<68> B_WLB<67> B_WLB<66> B_WLB<65> B_WLB<64> B_WLB<63> 
+ B_WLB<62> B_WLB<61> B_WLB<60> B_WLB<59> B_WLB<58> B_WLB<57> B_WLB<56> B_WLB<55> B_WLB<54> 
+ B_WLB<53> B_WLB<52> B_WLB<51> B_WLB<50> B_WLB<49> B_WLB<48> B_WLB<47> B_WLB<46> B_WLB<45> 
+ B_WLB<44> B_WLB<43> B_WLB<42> B_WLB<41> B_WLB<40> B_WLB<39> B_WLB<38> B_WLB<37> B_WLB<36> 
+ B_WLB<35> B_WLB<34> B_WLB<33> B_WLB<32> B_WLB<31> B_WLB<30> B_WLB<29> B_WLB<28> B_WLB<27> 
+ B_WLB<26> B_WLB<25> B_WLB<24> B_WLB<23> B_WLB<22> B_WLB<21> B_WLB<20> B_WLB<19> B_WLB<18> 
+ B_WLB<17> B_WLB<16> B_WLB<15> B_WLB<14> B_WLB<13> B_WLB<12> B_WLB<11> B_WLB<10> B_WLB<9> 
+ B_WLB<8> B_WLB<7> B_WLB<6> B_WLB<5> B_WLB<4> B_WLB<3> B_WLB<2> B_WLB<1> B_WLB<0> 
+  / dpram16x4096_AR_COLX8_ROWX256
XAR_TOP<1>
+ T_BLA<3> T_BLA<2> T_BLA_N<3> T_BLA_N<2> T_BLB<3> T_BLB<2> T_BLB_N<3> T_BLB_N<2> VSS 
+ VDD T_WLA<255> T_WLA<254> T_WLA<253> T_WLA<252> T_WLA<251> T_WLA<250> T_WLA<249> T_WLA<248> 
+ T_WLA<247> T_WLA<246> T_WLA<245> T_WLA<244> T_WLA<243> T_WLA<242> T_WLA<241> T_WLA<240> T_WLA<239> 
+ T_WLA<238> T_WLA<237> T_WLA<236> T_WLA<235> T_WLA<234> T_WLA<233> T_WLA<232> T_WLA<231> T_WLA<230> 
+ T_WLA<229> T_WLA<228> T_WLA<227> T_WLA<226> T_WLA<225> T_WLA<224> T_WLA<223> T_WLA<222> T_WLA<221> 
+ T_WLA<220> T_WLA<219> T_WLA<218> T_WLA<217> T_WLA<216> T_WLA<215> T_WLA<214> T_WLA<213> T_WLA<212> 
+ T_WLA<211> T_WLA<210> T_WLA<209> T_WLA<208> T_WLA<207> T_WLA<206> T_WLA<205> T_WLA<204> T_WLA<203> 
+ T_WLA<202> T_WLA<201> T_WLA<200> T_WLA<199> T_WLA<198> T_WLA<197> T_WLA<196> T_WLA<195> T_WLA<194> 
+ T_WLA<193> T_WLA<192> T_WLA<191> T_WLA<190> T_WLA<189> T_WLA<188> T_WLA<187> T_WLA<186> T_WLA<185> 
+ T_WLA<184> T_WLA<183> T_WLA<182> T_WLA<181> T_WLA<180> T_WLA<179> T_WLA<178> T_WLA<177> T_WLA<176> 
+ T_WLA<175> T_WLA<174> T_WLA<173> T_WLA<172> T_WLA<171> T_WLA<170> T_WLA<169> T_WLA<168> T_WLA<167> 
+ T_WLA<166> T_WLA<165> T_WLA<164> T_WLA<163> T_WLA<162> T_WLA<161> T_WLA<160> T_WLA<159> T_WLA<158> 
+ T_WLA<157> T_WLA<156> T_WLA<155> T_WLA<154> T_WLA<153> T_WLA<152> T_WLA<151> T_WLA<150> T_WLA<149> 
+ T_WLA<148> T_WLA<147> T_WLA<146> T_WLA<145> T_WLA<144> T_WLA<143> T_WLA<142> T_WLA<141> T_WLA<140> 
+ T_WLA<139> T_WLA<138> T_WLA<137> T_WLA<136> T_WLA<135> T_WLA<134> T_WLA<133> T_WLA<132> T_WLA<131> 
+ T_WLA<130> T_WLA<129> T_WLA<128> T_WLA<127> T_WLA<126> T_WLA<125> T_WLA<124> T_WLA<123> T_WLA<122> 
+ T_WLA<121> T_WLA<120> T_WLA<119> T_WLA<118> T_WLA<117> T_WLA<116> T_WLA<115> T_WLA<114> T_WLA<113> 
+ T_WLA<112> T_WLA<111> T_WLA<110> T_WLA<109> T_WLA<108> T_WLA<107> T_WLA<106> T_WLA<105> T_WLA<104> 
+ T_WLA<103> T_WLA<102> T_WLA<101> T_WLA<100> T_WLA<99> T_WLA<98> T_WLA<97> T_WLA<96> T_WLA<95> 
+ T_WLA<94> T_WLA<93> T_WLA<92> T_WLA<91> T_WLA<90> T_WLA<89> T_WLA<88> T_WLA<87> T_WLA<86> 
+ T_WLA<85> T_WLA<84> T_WLA<83> T_WLA<82> T_WLA<81> T_WLA<80> T_WLA<79> T_WLA<78> T_WLA<77> 
+ T_WLA<76> T_WLA<75> T_WLA<74> T_WLA<73> T_WLA<72> T_WLA<71> T_WLA<70> T_WLA<69> T_WLA<68> 
+ T_WLA<67> T_WLA<66> T_WLA<65> T_WLA<64> T_WLA<63> T_WLA<62> T_WLA<61> T_WLA<60> T_WLA<59> 
+ T_WLA<58> T_WLA<57> T_WLA<56> T_WLA<55> T_WLA<54> T_WLA<53> T_WLA<52> T_WLA<51> T_WLA<50> 
+ T_WLA<49> T_WLA<48> T_WLA<47> T_WLA<46> T_WLA<45> T_WLA<44> T_WLA<43> T_WLA<42> T_WLA<41> 
+ T_WLA<40> T_WLA<39> T_WLA<38> T_WLA<37> T_WLA<36> T_WLA<35> T_WLA<34> T_WLA<33> T_WLA<32> 
+ T_WLA<31> T_WLA<30> T_WLA<29> T_WLA<28> T_WLA<27> T_WLA<26> T_WLA<25> T_WLA<24> T_WLA<23> 
+ T_WLA<22> T_WLA<21> T_WLA<20> T_WLA<19> T_WLA<18> T_WLA<17> T_WLA<16> T_WLA<15> T_WLA<14> 
+ T_WLA<13> T_WLA<12> T_WLA<11> T_WLA<10> T_WLA<9> T_WLA<8> T_WLA<7> T_WLA<6> T_WLA<5> 
+ T_WLA<4> T_WLA<3> T_WLA<2> T_WLA<1> T_WLA<0> T_WLB<255> T_WLB<254> T_WLB<253> T_WLB<252> 
+ T_WLB<251> T_WLB<250> T_WLB<249> T_WLB<248> T_WLB<247> T_WLB<246> T_WLB<245> T_WLB<244> T_WLB<243> 
+ T_WLB<242> T_WLB<241> T_WLB<240> T_WLB<239> T_WLB<238> T_WLB<237> T_WLB<236> T_WLB<235> T_WLB<234> 
+ T_WLB<233> T_WLB<232> T_WLB<231> T_WLB<230> T_WLB<229> T_WLB<228> T_WLB<227> T_WLB<226> T_WLB<225> 
+ T_WLB<224> T_WLB<223> T_WLB<222> T_WLB<221> T_WLB<220> T_WLB<219> T_WLB<218> T_WLB<217> T_WLB<216> 
+ T_WLB<215> T_WLB<214> T_WLB<213> T_WLB<212> T_WLB<211> T_WLB<210> T_WLB<209> T_WLB<208> T_WLB<207> 
+ T_WLB<206> T_WLB<205> T_WLB<204> T_WLB<203> T_WLB<202> T_WLB<201> T_WLB<200> T_WLB<199> T_WLB<198> 
+ T_WLB<197> T_WLB<196> T_WLB<195> T_WLB<194> T_WLB<193> T_WLB<192> T_WLB<191> T_WLB<190> T_WLB<189> 
+ T_WLB<188> T_WLB<187> T_WLB<186> T_WLB<185> T_WLB<184> T_WLB<183> T_WLB<182> T_WLB<181> T_WLB<180> 
+ T_WLB<179> T_WLB<178> T_WLB<177> T_WLB<176> T_WLB<175> T_WLB<174> T_WLB<173> T_WLB<172> T_WLB<171> 
+ T_WLB<170> T_WLB<169> T_WLB<168> T_WLB<167> T_WLB<166> T_WLB<165> T_WLB<164> T_WLB<163> T_WLB<162> 
+ T_WLB<161> T_WLB<160> T_WLB<159> T_WLB<158> T_WLB<157> T_WLB<156> T_WLB<155> T_WLB<154> T_WLB<153> 
+ T_WLB<152> T_WLB<151> T_WLB<150> T_WLB<149> T_WLB<148> T_WLB<147> T_WLB<146> T_WLB<145> T_WLB<144> 
+ T_WLB<143> T_WLB<142> T_WLB<141> T_WLB<140> T_WLB<139> T_WLB<138> T_WLB<137> T_WLB<136> T_WLB<135> 
+ T_WLB<134> T_WLB<133> T_WLB<132> T_WLB<131> T_WLB<130> T_WLB<129> T_WLB<128> T_WLB<127> T_WLB<126> 
+ T_WLB<125> T_WLB<124> T_WLB<123> T_WLB<122> T_WLB<121> T_WLB<120> T_WLB<119> T_WLB<118> T_WLB<117> 
+ T_WLB<116> T_WLB<115> T_WLB<114> T_WLB<113> T_WLB<112> T_WLB<111> T_WLB<110> T_WLB<109> T_WLB<108> 
+ T_WLB<107> T_WLB<106> T_WLB<105> T_WLB<104> T_WLB<103> T_WLB<102> T_WLB<101> T_WLB<100> T_WLB<99> 
+ T_WLB<98> T_WLB<97> T_WLB<96> T_WLB<95> T_WLB<94> T_WLB<93> T_WLB<92> T_WLB<91> T_WLB<90> 
+ T_WLB<89> T_WLB<88> T_WLB<87> T_WLB<86> T_WLB<85> T_WLB<84> T_WLB<83> T_WLB<82> T_WLB<81> 
+ T_WLB<80> T_WLB<79> T_WLB<78> T_WLB<77> T_WLB<76> T_WLB<75> T_WLB<74> T_WLB<73> T_WLB<72> 
+ T_WLB<71> T_WLB<70> T_WLB<69> T_WLB<68> T_WLB<67> T_WLB<66> T_WLB<65> T_WLB<64> T_WLB<63> 
+ T_WLB<62> T_WLB<61> T_WLB<60> T_WLB<59> T_WLB<58> T_WLB<57> T_WLB<56> T_WLB<55> T_WLB<54> 
+ T_WLB<53> T_WLB<52> T_WLB<51> T_WLB<50> T_WLB<49> T_WLB<48> T_WLB<47> T_WLB<46> T_WLB<45> 
+ T_WLB<44> T_WLB<43> T_WLB<42> T_WLB<41> T_WLB<40> T_WLB<39> T_WLB<38> T_WLB<37> T_WLB<36> 
+ T_WLB<35> T_WLB<34> T_WLB<33> T_WLB<32> T_WLB<31> T_WLB<30> T_WLB<29> T_WLB<28> T_WLB<27> 
+ T_WLB<26> T_WLB<25> T_WLB<24> T_WLB<23> T_WLB<22> T_WLB<21> T_WLB<20> T_WLB<19> T_WLB<18> 
+ T_WLB<17> T_WLB<16> T_WLB<15> T_WLB<14> T_WLB<13> T_WLB<12> T_WLB<11> T_WLB<10> T_WLB<9> 
+ T_WLB<8> T_WLB<7> T_WLB<6> T_WLB<5> T_WLB<4> T_WLB<3> T_WLB<2> T_WLB<1> T_WLB<0> 
+  / dpram16x4096_AR_COLX8_ROWX256
XAR_BOT<1>
+ B_BLA<3> B_BLA<2> B_BLA_N<3> B_BLA_N<2> B_BLB<3> B_BLB<2> B_BLB_N<3> B_BLB_N<2> VSS 
+ VDD B_WLA<255> B_WLA<254> B_WLA<253> B_WLA<252> B_WLA<251> B_WLA<250> B_WLA<249> B_WLA<248> 
+ B_WLA<247> B_WLA<246> B_WLA<245> B_WLA<244> B_WLA<243> B_WLA<242> B_WLA<241> B_WLA<240> B_WLA<239> 
+ B_WLA<238> B_WLA<237> B_WLA<236> B_WLA<235> B_WLA<234> B_WLA<233> B_WLA<232> B_WLA<231> B_WLA<230> 
+ B_WLA<229> B_WLA<228> B_WLA<227> B_WLA<226> B_WLA<225> B_WLA<224> B_WLA<223> B_WLA<222> B_WLA<221> 
+ B_WLA<220> B_WLA<219> B_WLA<218> B_WLA<217> B_WLA<216> B_WLA<215> B_WLA<214> B_WLA<213> B_WLA<212> 
+ B_WLA<211> B_WLA<210> B_WLA<209> B_WLA<208> B_WLA<207> B_WLA<206> B_WLA<205> B_WLA<204> B_WLA<203> 
+ B_WLA<202> B_WLA<201> B_WLA<200> B_WLA<199> B_WLA<198> B_WLA<197> B_WLA<196> B_WLA<195> B_WLA<194> 
+ B_WLA<193> B_WLA<192> B_WLA<191> B_WLA<190> B_WLA<189> B_WLA<188> B_WLA<187> B_WLA<186> B_WLA<185> 
+ B_WLA<184> B_WLA<183> B_WLA<182> B_WLA<181> B_WLA<180> B_WLA<179> B_WLA<178> B_WLA<177> B_WLA<176> 
+ B_WLA<175> B_WLA<174> B_WLA<173> B_WLA<172> B_WLA<171> B_WLA<170> B_WLA<169> B_WLA<168> B_WLA<167> 
+ B_WLA<166> B_WLA<165> B_WLA<164> B_WLA<163> B_WLA<162> B_WLA<161> B_WLA<160> B_WLA<159> B_WLA<158> 
+ B_WLA<157> B_WLA<156> B_WLA<155> B_WLA<154> B_WLA<153> B_WLA<152> B_WLA<151> B_WLA<150> B_WLA<149> 
+ B_WLA<148> B_WLA<147> B_WLA<146> B_WLA<145> B_WLA<144> B_WLA<143> B_WLA<142> B_WLA<141> B_WLA<140> 
+ B_WLA<139> B_WLA<138> B_WLA<137> B_WLA<136> B_WLA<135> B_WLA<134> B_WLA<133> B_WLA<132> B_WLA<131> 
+ B_WLA<130> B_WLA<129> B_WLA<128> B_WLA<127> B_WLA<126> B_WLA<125> B_WLA<124> B_WLA<123> B_WLA<122> 
+ B_WLA<121> B_WLA<120> B_WLA<119> B_WLA<118> B_WLA<117> B_WLA<116> B_WLA<115> B_WLA<114> B_WLA<113> 
+ B_WLA<112> B_WLA<111> B_WLA<110> B_WLA<109> B_WLA<108> B_WLA<107> B_WLA<106> B_WLA<105> B_WLA<104> 
+ B_WLA<103> B_WLA<102> B_WLA<101> B_WLA<100> B_WLA<99> B_WLA<98> B_WLA<97> B_WLA<96> B_WLA<95> 
+ B_WLA<94> B_WLA<93> B_WLA<92> B_WLA<91> B_WLA<90> B_WLA<89> B_WLA<88> B_WLA<87> B_WLA<86> 
+ B_WLA<85> B_WLA<84> B_WLA<83> B_WLA<82> B_WLA<81> B_WLA<80> B_WLA<79> B_WLA<78> B_WLA<77> 
+ B_WLA<76> B_WLA<75> B_WLA<74> B_WLA<73> B_WLA<72> B_WLA<71> B_WLA<70> B_WLA<69> B_WLA<68> 
+ B_WLA<67> B_WLA<66> B_WLA<65> B_WLA<64> B_WLA<63> B_WLA<62> B_WLA<61> B_WLA<60> B_WLA<59> 
+ B_WLA<58> B_WLA<57> B_WLA<56> B_WLA<55> B_WLA<54> B_WLA<53> B_WLA<52> B_WLA<51> B_WLA<50> 
+ B_WLA<49> B_WLA<48> B_WLA<47> B_WLA<46> B_WLA<45> B_WLA<44> B_WLA<43> B_WLA<42> B_WLA<41> 
+ B_WLA<40> B_WLA<39> B_WLA<38> B_WLA<37> B_WLA<36> B_WLA<35> B_WLA<34> B_WLA<33> B_WLA<32> 
+ B_WLA<31> B_WLA<30> B_WLA<29> B_WLA<28> B_WLA<27> B_WLA<26> B_WLA<25> B_WLA<24> B_WLA<23> 
+ B_WLA<22> B_WLA<21> B_WLA<20> B_WLA<19> B_WLA<18> B_WLA<17> B_WLA<16> B_WLA<15> B_WLA<14> 
+ B_WLA<13> B_WLA<12> B_WLA<11> B_WLA<10> B_WLA<9> B_WLA<8> B_WLA<7> B_WLA<6> B_WLA<5> 
+ B_WLA<4> B_WLA<3> B_WLA<2> B_WLA<1> B_WLA<0> B_WLB<255> B_WLB<254> B_WLB<253> B_WLB<252> 
+ B_WLB<251> B_WLB<250> B_WLB<249> B_WLB<248> B_WLB<247> B_WLB<246> B_WLB<245> B_WLB<244> B_WLB<243> 
+ B_WLB<242> B_WLB<241> B_WLB<240> B_WLB<239> B_WLB<238> B_WLB<237> B_WLB<236> B_WLB<235> B_WLB<234> 
+ B_WLB<233> B_WLB<232> B_WLB<231> B_WLB<230> B_WLB<229> B_WLB<228> B_WLB<227> B_WLB<226> B_WLB<225> 
+ B_WLB<224> B_WLB<223> B_WLB<222> B_WLB<221> B_WLB<220> B_WLB<219> B_WLB<218> B_WLB<217> B_WLB<216> 
+ B_WLB<215> B_WLB<214> B_WLB<213> B_WLB<212> B_WLB<211> B_WLB<210> B_WLB<209> B_WLB<208> B_WLB<207> 
+ B_WLB<206> B_WLB<205> B_WLB<204> B_WLB<203> B_WLB<202> B_WLB<201> B_WLB<200> B_WLB<199> B_WLB<198> 
+ B_WLB<197> B_WLB<196> B_WLB<195> B_WLB<194> B_WLB<193> B_WLB<192> B_WLB<191> B_WLB<190> B_WLB<189> 
+ B_WLB<188> B_WLB<187> B_WLB<186> B_WLB<185> B_WLB<184> B_WLB<183> B_WLB<182> B_WLB<181> B_WLB<180> 
+ B_WLB<179> B_WLB<178> B_WLB<177> B_WLB<176> B_WLB<175> B_WLB<174> B_WLB<173> B_WLB<172> B_WLB<171> 
+ B_WLB<170> B_WLB<169> B_WLB<168> B_WLB<167> B_WLB<166> B_WLB<165> B_WLB<164> B_WLB<163> B_WLB<162> 
+ B_WLB<161> B_WLB<160> B_WLB<159> B_WLB<158> B_WLB<157> B_WLB<156> B_WLB<155> B_WLB<154> B_WLB<153> 
+ B_WLB<152> B_WLB<151> B_WLB<150> B_WLB<149> B_WLB<148> B_WLB<147> B_WLB<146> B_WLB<145> B_WLB<144> 
+ B_WLB<143> B_WLB<142> B_WLB<141> B_WLB<140> B_WLB<139> B_WLB<138> B_WLB<137> B_WLB<136> B_WLB<135> 
+ B_WLB<134> B_WLB<133> B_WLB<132> B_WLB<131> B_WLB<130> B_WLB<129> B_WLB<128> B_WLB<127> B_WLB<126> 
+ B_WLB<125> B_WLB<124> B_WLB<123> B_WLB<122> B_WLB<121> B_WLB<120> B_WLB<119> B_WLB<118> B_WLB<117> 
+ B_WLB<116> B_WLB<115> B_WLB<114> B_WLB<113> B_WLB<112> B_WLB<111> B_WLB<110> B_WLB<109> B_WLB<108> 
+ B_WLB<107> B_WLB<106> B_WLB<105> B_WLB<104> B_WLB<103> B_WLB<102> B_WLB<101> B_WLB<100> B_WLB<99> 
+ B_WLB<98> B_WLB<97> B_WLB<96> B_WLB<95> B_WLB<94> B_WLB<93> B_WLB<92> B_WLB<91> B_WLB<90> 
+ B_WLB<89> B_WLB<88> B_WLB<87> B_WLB<86> B_WLB<85> B_WLB<84> B_WLB<83> B_WLB<82> B_WLB<81> 
+ B_WLB<80> B_WLB<79> B_WLB<78> B_WLB<77> B_WLB<76> B_WLB<75> B_WLB<74> B_WLB<73> B_WLB<72> 
+ B_WLB<71> B_WLB<70> B_WLB<69> B_WLB<68> B_WLB<67> B_WLB<66> B_WLB<65> B_WLB<64> B_WLB<63> 
+ B_WLB<62> B_WLB<61> B_WLB<60> B_WLB<59> B_WLB<58> B_WLB<57> B_WLB<56> B_WLB<55> B_WLB<54> 
+ B_WLB<53> B_WLB<52> B_WLB<51> B_WLB<50> B_WLB<49> B_WLB<48> B_WLB<47> B_WLB<46> B_WLB<45> 
+ B_WLB<44> B_WLB<43> B_WLB<42> B_WLB<41> B_WLB<40> B_WLB<39> B_WLB<38> B_WLB<37> B_WLB<36> 
+ B_WLB<35> B_WLB<34> B_WLB<33> B_WLB<32> B_WLB<31> B_WLB<30> B_WLB<29> B_WLB<28> B_WLB<27> 
+ B_WLB<26> B_WLB<25> B_WLB<24> B_WLB<23> B_WLB<22> B_WLB<21> B_WLB<20> B_WLB<19> B_WLB<18> 
+ B_WLB<17> B_WLB<16> B_WLB<15> B_WLB<14> B_WLB<13> B_WLB<12> B_WLB<11> B_WLB<10> B_WLB<9> 
+ B_WLB<8> B_WLB<7> B_WLB<6> B_WLB<5> B_WLB<4> B_WLB<3> B_WLB<2> B_WLB<1> B_WLB<0> 
+  / dpram16x4096_AR_COLX8_ROWX256
XAR_TOP<0>
+ T_BLA<1> T_BLA<0> T_BLA_N<1> T_BLA_N<0> T_BLB<1> T_BLB<0> T_BLB_N<1> T_BLB_N<0> VSS 
+ VDD T_WLA<255> T_WLA<254> T_WLA<253> T_WLA<252> T_WLA<251> T_WLA<250> T_WLA<249> T_WLA<248> 
+ T_WLA<247> T_WLA<246> T_WLA<245> T_WLA<244> T_WLA<243> T_WLA<242> T_WLA<241> T_WLA<240> T_WLA<239> 
+ T_WLA<238> T_WLA<237> T_WLA<236> T_WLA<235> T_WLA<234> T_WLA<233> T_WLA<232> T_WLA<231> T_WLA<230> 
+ T_WLA<229> T_WLA<228> T_WLA<227> T_WLA<226> T_WLA<225> T_WLA<224> T_WLA<223> T_WLA<222> T_WLA<221> 
+ T_WLA<220> T_WLA<219> T_WLA<218> T_WLA<217> T_WLA<216> T_WLA<215> T_WLA<214> T_WLA<213> T_WLA<212> 
+ T_WLA<211> T_WLA<210> T_WLA<209> T_WLA<208> T_WLA<207> T_WLA<206> T_WLA<205> T_WLA<204> T_WLA<203> 
+ T_WLA<202> T_WLA<201> T_WLA<200> T_WLA<199> T_WLA<198> T_WLA<197> T_WLA<196> T_WLA<195> T_WLA<194> 
+ T_WLA<193> T_WLA<192> T_WLA<191> T_WLA<190> T_WLA<189> T_WLA<188> T_WLA<187> T_WLA<186> T_WLA<185> 
+ T_WLA<184> T_WLA<183> T_WLA<182> T_WLA<181> T_WLA<180> T_WLA<179> T_WLA<178> T_WLA<177> T_WLA<176> 
+ T_WLA<175> T_WLA<174> T_WLA<173> T_WLA<172> T_WLA<171> T_WLA<170> T_WLA<169> T_WLA<168> T_WLA<167> 
+ T_WLA<166> T_WLA<165> T_WLA<164> T_WLA<163> T_WLA<162> T_WLA<161> T_WLA<160> T_WLA<159> T_WLA<158> 
+ T_WLA<157> T_WLA<156> T_WLA<155> T_WLA<154> T_WLA<153> T_WLA<152> T_WLA<151> T_WLA<150> T_WLA<149> 
+ T_WLA<148> T_WLA<147> T_WLA<146> T_WLA<145> T_WLA<144> T_WLA<143> T_WLA<142> T_WLA<141> T_WLA<140> 
+ T_WLA<139> T_WLA<138> T_WLA<137> T_WLA<136> T_WLA<135> T_WLA<134> T_WLA<133> T_WLA<132> T_WLA<131> 
+ T_WLA<130> T_WLA<129> T_WLA<128> T_WLA<127> T_WLA<126> T_WLA<125> T_WLA<124> T_WLA<123> T_WLA<122> 
+ T_WLA<121> T_WLA<120> T_WLA<119> T_WLA<118> T_WLA<117> T_WLA<116> T_WLA<115> T_WLA<114> T_WLA<113> 
+ T_WLA<112> T_WLA<111> T_WLA<110> T_WLA<109> T_WLA<108> T_WLA<107> T_WLA<106> T_WLA<105> T_WLA<104> 
+ T_WLA<103> T_WLA<102> T_WLA<101> T_WLA<100> T_WLA<99> T_WLA<98> T_WLA<97> T_WLA<96> T_WLA<95> 
+ T_WLA<94> T_WLA<93> T_WLA<92> T_WLA<91> T_WLA<90> T_WLA<89> T_WLA<88> T_WLA<87> T_WLA<86> 
+ T_WLA<85> T_WLA<84> T_WLA<83> T_WLA<82> T_WLA<81> T_WLA<80> T_WLA<79> T_WLA<78> T_WLA<77> 
+ T_WLA<76> T_WLA<75> T_WLA<74> T_WLA<73> T_WLA<72> T_WLA<71> T_WLA<70> T_WLA<69> T_WLA<68> 
+ T_WLA<67> T_WLA<66> T_WLA<65> T_WLA<64> T_WLA<63> T_WLA<62> T_WLA<61> T_WLA<60> T_WLA<59> 
+ T_WLA<58> T_WLA<57> T_WLA<56> T_WLA<55> T_WLA<54> T_WLA<53> T_WLA<52> T_WLA<51> T_WLA<50> 
+ T_WLA<49> T_WLA<48> T_WLA<47> T_WLA<46> T_WLA<45> T_WLA<44> T_WLA<43> T_WLA<42> T_WLA<41> 
+ T_WLA<40> T_WLA<39> T_WLA<38> T_WLA<37> T_WLA<36> T_WLA<35> T_WLA<34> T_WLA<33> T_WLA<32> 
+ T_WLA<31> T_WLA<30> T_WLA<29> T_WLA<28> T_WLA<27> T_WLA<26> T_WLA<25> T_WLA<24> T_WLA<23> 
+ T_WLA<22> T_WLA<21> T_WLA<20> T_WLA<19> T_WLA<18> T_WLA<17> T_WLA<16> T_WLA<15> T_WLA<14> 
+ T_WLA<13> T_WLA<12> T_WLA<11> T_WLA<10> T_WLA<9> T_WLA<8> T_WLA<7> T_WLA<6> T_WLA<5> 
+ T_WLA<4> T_WLA<3> T_WLA<2> T_WLA<1> T_WLA<0> T_WLB<255> T_WLB<254> T_WLB<253> T_WLB<252> 
+ T_WLB<251> T_WLB<250> T_WLB<249> T_WLB<248> T_WLB<247> T_WLB<246> T_WLB<245> T_WLB<244> T_WLB<243> 
+ T_WLB<242> T_WLB<241> T_WLB<240> T_WLB<239> T_WLB<238> T_WLB<237> T_WLB<236> T_WLB<235> T_WLB<234> 
+ T_WLB<233> T_WLB<232> T_WLB<231> T_WLB<230> T_WLB<229> T_WLB<228> T_WLB<227> T_WLB<226> T_WLB<225> 
+ T_WLB<224> T_WLB<223> T_WLB<222> T_WLB<221> T_WLB<220> T_WLB<219> T_WLB<218> T_WLB<217> T_WLB<216> 
+ T_WLB<215> T_WLB<214> T_WLB<213> T_WLB<212> T_WLB<211> T_WLB<210> T_WLB<209> T_WLB<208> T_WLB<207> 
+ T_WLB<206> T_WLB<205> T_WLB<204> T_WLB<203> T_WLB<202> T_WLB<201> T_WLB<200> T_WLB<199> T_WLB<198> 
+ T_WLB<197> T_WLB<196> T_WLB<195> T_WLB<194> T_WLB<193> T_WLB<192> T_WLB<191> T_WLB<190> T_WLB<189> 
+ T_WLB<188> T_WLB<187> T_WLB<186> T_WLB<185> T_WLB<184> T_WLB<183> T_WLB<182> T_WLB<181> T_WLB<180> 
+ T_WLB<179> T_WLB<178> T_WLB<177> T_WLB<176> T_WLB<175> T_WLB<174> T_WLB<173> T_WLB<172> T_WLB<171> 
+ T_WLB<170> T_WLB<169> T_WLB<168> T_WLB<167> T_WLB<166> T_WLB<165> T_WLB<164> T_WLB<163> T_WLB<162> 
+ T_WLB<161> T_WLB<160> T_WLB<159> T_WLB<158> T_WLB<157> T_WLB<156> T_WLB<155> T_WLB<154> T_WLB<153> 
+ T_WLB<152> T_WLB<151> T_WLB<150> T_WLB<149> T_WLB<148> T_WLB<147> T_WLB<146> T_WLB<145> T_WLB<144> 
+ T_WLB<143> T_WLB<142> T_WLB<141> T_WLB<140> T_WLB<139> T_WLB<138> T_WLB<137> T_WLB<136> T_WLB<135> 
+ T_WLB<134> T_WLB<133> T_WLB<132> T_WLB<131> T_WLB<130> T_WLB<129> T_WLB<128> T_WLB<127> T_WLB<126> 
+ T_WLB<125> T_WLB<124> T_WLB<123> T_WLB<122> T_WLB<121> T_WLB<120> T_WLB<119> T_WLB<118> T_WLB<117> 
+ T_WLB<116> T_WLB<115> T_WLB<114> T_WLB<113> T_WLB<112> T_WLB<111> T_WLB<110> T_WLB<109> T_WLB<108> 
+ T_WLB<107> T_WLB<106> T_WLB<105> T_WLB<104> T_WLB<103> T_WLB<102> T_WLB<101> T_WLB<100> T_WLB<99> 
+ T_WLB<98> T_WLB<97> T_WLB<96> T_WLB<95> T_WLB<94> T_WLB<93> T_WLB<92> T_WLB<91> T_WLB<90> 
+ T_WLB<89> T_WLB<88> T_WLB<87> T_WLB<86> T_WLB<85> T_WLB<84> T_WLB<83> T_WLB<82> T_WLB<81> 
+ T_WLB<80> T_WLB<79> T_WLB<78> T_WLB<77> T_WLB<76> T_WLB<75> T_WLB<74> T_WLB<73> T_WLB<72> 
+ T_WLB<71> T_WLB<70> T_WLB<69> T_WLB<68> T_WLB<67> T_WLB<66> T_WLB<65> T_WLB<64> T_WLB<63> 
+ T_WLB<62> T_WLB<61> T_WLB<60> T_WLB<59> T_WLB<58> T_WLB<57> T_WLB<56> T_WLB<55> T_WLB<54> 
+ T_WLB<53> T_WLB<52> T_WLB<51> T_WLB<50> T_WLB<49> T_WLB<48> T_WLB<47> T_WLB<46> T_WLB<45> 
+ T_WLB<44> T_WLB<43> T_WLB<42> T_WLB<41> T_WLB<40> T_WLB<39> T_WLB<38> T_WLB<37> T_WLB<36> 
+ T_WLB<35> T_WLB<34> T_WLB<33> T_WLB<32> T_WLB<31> T_WLB<30> T_WLB<29> T_WLB<28> T_WLB<27> 
+ T_WLB<26> T_WLB<25> T_WLB<24> T_WLB<23> T_WLB<22> T_WLB<21> T_WLB<20> T_WLB<19> T_WLB<18> 
+ T_WLB<17> T_WLB<16> T_WLB<15> T_WLB<14> T_WLB<13> T_WLB<12> T_WLB<11> T_WLB<10> T_WLB<9> 
+ T_WLB<8> T_WLB<7> T_WLB<6> T_WLB<5> T_WLB<4> T_WLB<3> T_WLB<2> T_WLB<1> T_WLB<0> 
+  / dpram16x4096_AR_COLX8_ROWX256
XAR_BOT<0>
+ B_BLA<1> B_BLA<0> B_BLA_N<1> B_BLA_N<0> B_BLB<1> B_BLB<0> B_BLB_N<1> B_BLB_N<0> VSS 
+ VDD B_WLA<255> B_WLA<254> B_WLA<253> B_WLA<252> B_WLA<251> B_WLA<250> B_WLA<249> B_WLA<248> 
+ B_WLA<247> B_WLA<246> B_WLA<245> B_WLA<244> B_WLA<243> B_WLA<242> B_WLA<241> B_WLA<240> B_WLA<239> 
+ B_WLA<238> B_WLA<237> B_WLA<236> B_WLA<235> B_WLA<234> B_WLA<233> B_WLA<232> B_WLA<231> B_WLA<230> 
+ B_WLA<229> B_WLA<228> B_WLA<227> B_WLA<226> B_WLA<225> B_WLA<224> B_WLA<223> B_WLA<222> B_WLA<221> 
+ B_WLA<220> B_WLA<219> B_WLA<218> B_WLA<217> B_WLA<216> B_WLA<215> B_WLA<214> B_WLA<213> B_WLA<212> 
+ B_WLA<211> B_WLA<210> B_WLA<209> B_WLA<208> B_WLA<207> B_WLA<206> B_WLA<205> B_WLA<204> B_WLA<203> 
+ B_WLA<202> B_WLA<201> B_WLA<200> B_WLA<199> B_WLA<198> B_WLA<197> B_WLA<196> B_WLA<195> B_WLA<194> 
+ B_WLA<193> B_WLA<192> B_WLA<191> B_WLA<190> B_WLA<189> B_WLA<188> B_WLA<187> B_WLA<186> B_WLA<185> 
+ B_WLA<184> B_WLA<183> B_WLA<182> B_WLA<181> B_WLA<180> B_WLA<179> B_WLA<178> B_WLA<177> B_WLA<176> 
+ B_WLA<175> B_WLA<174> B_WLA<173> B_WLA<172> B_WLA<171> B_WLA<170> B_WLA<169> B_WLA<168> B_WLA<167> 
+ B_WLA<166> B_WLA<165> B_WLA<164> B_WLA<163> B_WLA<162> B_WLA<161> B_WLA<160> B_WLA<159> B_WLA<158> 
+ B_WLA<157> B_WLA<156> B_WLA<155> B_WLA<154> B_WLA<153> B_WLA<152> B_WLA<151> B_WLA<150> B_WLA<149> 
+ B_WLA<148> B_WLA<147> B_WLA<146> B_WLA<145> B_WLA<144> B_WLA<143> B_WLA<142> B_WLA<141> B_WLA<140> 
+ B_WLA<139> B_WLA<138> B_WLA<137> B_WLA<136> B_WLA<135> B_WLA<134> B_WLA<133> B_WLA<132> B_WLA<131> 
+ B_WLA<130> B_WLA<129> B_WLA<128> B_WLA<127> B_WLA<126> B_WLA<125> B_WLA<124> B_WLA<123> B_WLA<122> 
+ B_WLA<121> B_WLA<120> B_WLA<119> B_WLA<118> B_WLA<117> B_WLA<116> B_WLA<115> B_WLA<114> B_WLA<113> 
+ B_WLA<112> B_WLA<111> B_WLA<110> B_WLA<109> B_WLA<108> B_WLA<107> B_WLA<106> B_WLA<105> B_WLA<104> 
+ B_WLA<103> B_WLA<102> B_WLA<101> B_WLA<100> B_WLA<99> B_WLA<98> B_WLA<97> B_WLA<96> B_WLA<95> 
+ B_WLA<94> B_WLA<93> B_WLA<92> B_WLA<91> B_WLA<90> B_WLA<89> B_WLA<88> B_WLA<87> B_WLA<86> 
+ B_WLA<85> B_WLA<84> B_WLA<83> B_WLA<82> B_WLA<81> B_WLA<80> B_WLA<79> B_WLA<78> B_WLA<77> 
+ B_WLA<76> B_WLA<75> B_WLA<74> B_WLA<73> B_WLA<72> B_WLA<71> B_WLA<70> B_WLA<69> B_WLA<68> 
+ B_WLA<67> B_WLA<66> B_WLA<65> B_WLA<64> B_WLA<63> B_WLA<62> B_WLA<61> B_WLA<60> B_WLA<59> 
+ B_WLA<58> B_WLA<57> B_WLA<56> B_WLA<55> B_WLA<54> B_WLA<53> B_WLA<52> B_WLA<51> B_WLA<50> 
+ B_WLA<49> B_WLA<48> B_WLA<47> B_WLA<46> B_WLA<45> B_WLA<44> B_WLA<43> B_WLA<42> B_WLA<41> 
+ B_WLA<40> B_WLA<39> B_WLA<38> B_WLA<37> B_WLA<36> B_WLA<35> B_WLA<34> B_WLA<33> B_WLA<32> 
+ B_WLA<31> B_WLA<30> B_WLA<29> B_WLA<28> B_WLA<27> B_WLA<26> B_WLA<25> B_WLA<24> B_WLA<23> 
+ B_WLA<22> B_WLA<21> B_WLA<20> B_WLA<19> B_WLA<18> B_WLA<17> B_WLA<16> B_WLA<15> B_WLA<14> 
+ B_WLA<13> B_WLA<12> B_WLA<11> B_WLA<10> B_WLA<9> B_WLA<8> B_WLA<7> B_WLA<6> B_WLA<5> 
+ B_WLA<4> B_WLA<3> B_WLA<2> B_WLA<1> B_WLA<0> B_WLB<255> B_WLB<254> B_WLB<253> B_WLB<252> 
+ B_WLB<251> B_WLB<250> B_WLB<249> B_WLB<248> B_WLB<247> B_WLB<246> B_WLB<245> B_WLB<244> B_WLB<243> 
+ B_WLB<242> B_WLB<241> B_WLB<240> B_WLB<239> B_WLB<238> B_WLB<237> B_WLB<236> B_WLB<235> B_WLB<234> 
+ B_WLB<233> B_WLB<232> B_WLB<231> B_WLB<230> B_WLB<229> B_WLB<228> B_WLB<227> B_WLB<226> B_WLB<225> 
+ B_WLB<224> B_WLB<223> B_WLB<222> B_WLB<221> B_WLB<220> B_WLB<219> B_WLB<218> B_WLB<217> B_WLB<216> 
+ B_WLB<215> B_WLB<214> B_WLB<213> B_WLB<212> B_WLB<211> B_WLB<210> B_WLB<209> B_WLB<208> B_WLB<207> 
+ B_WLB<206> B_WLB<205> B_WLB<204> B_WLB<203> B_WLB<202> B_WLB<201> B_WLB<200> B_WLB<199> B_WLB<198> 
+ B_WLB<197> B_WLB<196> B_WLB<195> B_WLB<194> B_WLB<193> B_WLB<192> B_WLB<191> B_WLB<190> B_WLB<189> 
+ B_WLB<188> B_WLB<187> B_WLB<186> B_WLB<185> B_WLB<184> B_WLB<183> B_WLB<182> B_WLB<181> B_WLB<180> 
+ B_WLB<179> B_WLB<178> B_WLB<177> B_WLB<176> B_WLB<175> B_WLB<174> B_WLB<173> B_WLB<172> B_WLB<171> 
+ B_WLB<170> B_WLB<169> B_WLB<168> B_WLB<167> B_WLB<166> B_WLB<165> B_WLB<164> B_WLB<163> B_WLB<162> 
+ B_WLB<161> B_WLB<160> B_WLB<159> B_WLB<158> B_WLB<157> B_WLB<156> B_WLB<155> B_WLB<154> B_WLB<153> 
+ B_WLB<152> B_WLB<151> B_WLB<150> B_WLB<149> B_WLB<148> B_WLB<147> B_WLB<146> B_WLB<145> B_WLB<144> 
+ B_WLB<143> B_WLB<142> B_WLB<141> B_WLB<140> B_WLB<139> B_WLB<138> B_WLB<137> B_WLB<136> B_WLB<135> 
+ B_WLB<134> B_WLB<133> B_WLB<132> B_WLB<131> B_WLB<130> B_WLB<129> B_WLB<128> B_WLB<127> B_WLB<126> 
+ B_WLB<125> B_WLB<124> B_WLB<123> B_WLB<122> B_WLB<121> B_WLB<120> B_WLB<119> B_WLB<118> B_WLB<117> 
+ B_WLB<116> B_WLB<115> B_WLB<114> B_WLB<113> B_WLB<112> B_WLB<111> B_WLB<110> B_WLB<109> B_WLB<108> 
+ B_WLB<107> B_WLB<106> B_WLB<105> B_WLB<104> B_WLB<103> B_WLB<102> B_WLB<101> B_WLB<100> B_WLB<99> 
+ B_WLB<98> B_WLB<97> B_WLB<96> B_WLB<95> B_WLB<94> B_WLB<93> B_WLB<92> B_WLB<91> B_WLB<90> 
+ B_WLB<89> B_WLB<88> B_WLB<87> B_WLB<86> B_WLB<85> B_WLB<84> B_WLB<83> B_WLB<82> B_WLB<81> 
+ B_WLB<80> B_WLB<79> B_WLB<78> B_WLB<77> B_WLB<76> B_WLB<75> B_WLB<74> B_WLB<73> B_WLB<72> 
+ B_WLB<71> B_WLB<70> B_WLB<69> B_WLB<68> B_WLB<67> B_WLB<66> B_WLB<65> B_WLB<64> B_WLB<63> 
+ B_WLB<62> B_WLB<61> B_WLB<60> B_WLB<59> B_WLB<58> B_WLB<57> B_WLB<56> B_WLB<55> B_WLB<54> 
+ B_WLB<53> B_WLB<52> B_WLB<51> B_WLB<50> B_WLB<49> B_WLB<48> B_WLB<47> B_WLB<46> B_WLB<45> 
+ B_WLB<44> B_WLB<43> B_WLB<42> B_WLB<41> B_WLB<40> B_WLB<39> B_WLB<38> B_WLB<37> B_WLB<36> 
+ B_WLB<35> B_WLB<34> B_WLB<33> B_WLB<32> B_WLB<31> B_WLB<30> B_WLB<29> B_WLB<28> B_WLB<27> 
+ B_WLB<26> B_WLB<25> B_WLB<24> B_WLB<23> B_WLB<22> B_WLB<21> B_WLB<20> B_WLB<19> B_WLB<18> 
+ B_WLB<17> B_WLB<16> B_WLB<15> B_WLB<14> B_WLB<13> B_WLB<12> B_WLB<11> B_WLB<10> B_WLB<9> 
+ B_WLB<8> B_WLB<7> B_WLB<6> B_WLB<5> B_WLB<4> B_WLB<3> B_WLB<2> B_WLB<1> B_WLB<0> 
+  / dpram16x4096_AR_COLX8_ROWX256
XBUF0
+ BWENA<0> BWENA_INT<0> BWENB<0> BWENB_INT<0> DA<0> DA_INT<0> DB<0> DB_INT<0> QA<0> 
+ QA_INT<0> QB<0> QB_INT<0> VDD VSS  / xmc55_dps_collar_dq_8_bw
XBUF1
+ BWENA<1> BWENA_INT<1> BWENB<1> BWENB_INT<1> DA<1> DA_INT<1> DB<1> DB_INT<1> QA<1> 
+ QA_INT<1> QB<1> QB_INT<1> VDD VSS  / xmc55_dps_collar_dq_8_bw
.ENDS

************************************************************************
* Cell Name:    dpram16x4096_XDECX256
* View Name:    schematic
************************************************************************
.SUBCKT dpram16x4096_XDECX256
+ PXAA<3> PXAA<2> PXAA<1> PXAA<0> PXAB<3> PXAB<2> PXAB<1> PXAB<0> PXBA_N<7> 
+ PXBA_N<6> PXBA_N<5> PXBA_N<4> PXBA_N<3> PXBA_N<2> PXBA_N<1> PXBA_N<0> PXBB_N<7> PXBB_N<6> 
+ PXBB_N<5> PXBB_N<4> PXBB_N<3> PXBB_N<2> PXBB_N<1> PXBB_N<0> PXCA_N<7> PXCA_N<6> PXCA_N<5> 
+ PXCA_N<4> PXCA_N<3> PXCA_N<2> PXCA_N<1> PXCA_N<0> PXCB_N<7> PXCB_N<6> PXCB_N<5> PXCB_N<4> 
+ PXCB_N<3> PXCB_N<2> PXCB_N<1> PXCB_N<0> VDD VSS WLA<255> WLA<254> WLA<253> 
+ WLA<252> WLA<251> WLA<250> WLA<249> WLA<248> WLA<247> WLA<246> WLA<245> WLA<244> 
+ WLA<243> WLA<242> WLA<241> WLA<240> WLA<239> WLA<238> WLA<237> WLA<236> WLA<235> 
+ WLA<234> WLA<233> WLA<232> WLA<231> WLA<230> WLA<229> WLA<228> WLA<227> WLA<226> 
+ WLA<225> WLA<224> WLA<223> WLA<222> WLA<221> WLA<220> WLA<219> WLA<218> WLA<217> 
+ WLA<216> WLA<215> WLA<214> WLA<213> WLA<212> WLA<211> WLA<210> WLA<209> WLA<208> 
+ WLA<207> WLA<206> WLA<205> WLA<204> WLA<203> WLA<202> WLA<201> WLA<200> WLA<199> 
+ WLA<198> WLA<197> WLA<196> WLA<195> WLA<194> WLA<193> WLA<192> WLA<191> WLA<190> 
+ WLA<189> WLA<188> WLA<187> WLA<186> WLA<185> WLA<184> WLA<183> WLA<182> WLA<181> 
+ WLA<180> WLA<179> WLA<178> WLA<177> WLA<176> WLA<175> WLA<174> WLA<173> WLA<172> 
+ WLA<171> WLA<170> WLA<169> WLA<168> WLA<167> WLA<166> WLA<165> WLA<164> WLA<163> 
+ WLA<162> WLA<161> WLA<160> WLA<159> WLA<158> WLA<157> WLA<156> WLA<155> WLA<154> 
+ WLA<153> WLA<152> WLA<151> WLA<150> WLA<149> WLA<148> WLA<147> WLA<146> WLA<145> 
+ WLA<144> WLA<143> WLA<142> WLA<141> WLA<140> WLA<139> WLA<138> WLA<137> WLA<136> 
+ WLA<135> WLA<134> WLA<133> WLA<132> WLA<131> WLA<130> WLA<129> WLA<128> WLA<127> 
+ WLA<126> WLA<125> WLA<124> WLA<123> WLA<122> WLA<121> WLA<120> WLA<119> WLA<118> 
+ WLA<117> WLA<116> WLA<115> WLA<114> WLA<113> WLA<112> WLA<111> WLA<110> WLA<109> 
+ WLA<108> WLA<107> WLA<106> WLA<105> WLA<104> WLA<103> WLA<102> WLA<101> WLA<100> 
+ WLA<99> WLA<98> WLA<97> WLA<96> WLA<95> WLA<94> WLA<93> WLA<92> WLA<91> 
+ WLA<90> WLA<89> WLA<88> WLA<87> WLA<86> WLA<85> WLA<84> WLA<83> WLA<82> 
+ WLA<81> WLA<80> WLA<79> WLA<78> WLA<77> WLA<76> WLA<75> WLA<74> WLA<73> 
+ WLA<72> WLA<71> WLA<70> WLA<69> WLA<68> WLA<67> WLA<66> WLA<65> WLA<64> 
+ WLA<63> WLA<62> WLA<61> WLA<60> WLA<59> WLA<58> WLA<57> WLA<56> WLA<55> 
+ WLA<54> WLA<53> WLA<52> WLA<51> WLA<50> WLA<49> WLA<48> WLA<47> WLA<46> 
+ WLA<45> WLA<44> WLA<43> WLA<42> WLA<41> WLA<40> WLA<39> WLA<38> WLA<37> 
+ WLA<36> WLA<35> WLA<34> WLA<33> WLA<32> WLA<31> WLA<30> WLA<29> WLA<28> 
+ WLA<27> WLA<26> WLA<25> WLA<24> WLA<23> WLA<22> WLA<21> WLA<20> WLA<19> 
+ WLA<18> WLA<17> WLA<16> WLA<15> WLA<14> WLA<13> WLA<12> WLA<11> WLA<10> 
+ WLA<9> WLA<8> WLA<7> WLA<6> WLA<5> WLA<4> WLA<3> WLA<2> WLA<1> 
+ WLA<0> WLB<255> WLB<254> WLB<253> WLB<252> WLB<251> WLB<250> WLB<249> WLB<248> 
+ WLB<247> WLB<246> WLB<245> WLB<244> WLB<243> WLB<242> WLB<241> WLB<240> WLB<239> 
+ WLB<238> WLB<237> WLB<236> WLB<235> WLB<234> WLB<233> WLB<232> WLB<231> WLB<230> 
+ WLB<229> WLB<228> WLB<227> WLB<226> WLB<225> WLB<224> WLB<223> WLB<222> WLB<221> 
+ WLB<220> WLB<219> WLB<218> WLB<217> WLB<216> WLB<215> WLB<214> WLB<213> WLB<212> 
+ WLB<211> WLB<210> WLB<209> WLB<208> WLB<207> WLB<206> WLB<205> WLB<204> WLB<203> 
+ WLB<202> WLB<201> WLB<200> WLB<199> WLB<198> WLB<197> WLB<196> WLB<195> WLB<194> 
+ WLB<193> WLB<192> WLB<191> WLB<190> WLB<189> WLB<188> WLB<187> WLB<186> WLB<185> 
+ WLB<184> WLB<183> WLB<182> WLB<181> WLB<180> WLB<179> WLB<178> WLB<177> WLB<176> 
+ WLB<175> WLB<174> WLB<173> WLB<172> WLB<171> WLB<170> WLB<169> WLB<168> WLB<167> 
+ WLB<166> WLB<165> WLB<164> WLB<163> WLB<162> WLB<161> WLB<160> WLB<159> WLB<158> 
+ WLB<157> WLB<156> WLB<155> WLB<154> WLB<153> WLB<152> WLB<151> WLB<150> WLB<149> 
+ WLB<148> WLB<147> WLB<146> WLB<145> WLB<144> WLB<143> WLB<142> WLB<141> WLB<140> 
+ WLB<139> WLB<138> WLB<137> WLB<136> WLB<135> WLB<134> WLB<133> WLB<132> WLB<131> 
+ WLB<130> WLB<129> WLB<128> WLB<127> WLB<126> WLB<125> WLB<124> WLB<123> WLB<122> 
+ WLB<121> WLB<120> WLB<119> WLB<118> WLB<117> WLB<116> WLB<115> WLB<114> WLB<113> 
+ WLB<112> WLB<111> WLB<110> WLB<109> WLB<108> WLB<107> WLB<106> WLB<105> WLB<104> 
+ WLB<103> WLB<102> WLB<101> WLB<100> WLB<99> WLB<98> WLB<97> WLB<96> WLB<95> 
+ WLB<94> WLB<93> WLB<92> WLB<91> WLB<90> WLB<89> WLB<88> WLB<87> WLB<86> 
+ WLB<85> WLB<84> WLB<83> WLB<82> WLB<81> WLB<80> WLB<79> WLB<78> WLB<77> 
+ WLB<76> WLB<75> WLB<74> WLB<73> WLB<72> WLB<71> WLB<70> WLB<69> WLB<68> 
+ WLB<67> WLB<66> WLB<65> WLB<64> WLB<63> WLB<62> WLB<61> WLB<60> WLB<59> 
+ WLB<58> WLB<57> WLB<56> WLB<55> WLB<54> WLB<53> WLB<52> WLB<51> WLB<50> 
+ WLB<49> WLB<48> WLB<47> WLB<46> WLB<45> WLB<44> WLB<43> WLB<42> WLB<41> 
+ WLB<40> WLB<39> WLB<38> WLB<37> WLB<36> WLB<35> WLB<34> WLB<33> WLB<32> 
+ WLB<31> WLB<30> WLB<29> WLB<28> WLB<27> WLB<26> WLB<25> WLB<24> WLB<23> 
+ WLB<22> WLB<21> WLB<20> WLB<19> WLB<18> WLB<17> WLB<16> WLB<15> WLB<14> 
+ WLB<13> WLB<12> WLB<11> WLB<10> WLB<9> WLB<8> WLB<7> WLB<6> WLB<5> 
+ WLB<4> WLB<3> WLB<2> WLB<1> WLB<0> 
XDUMMY_IN
+ VDD VSS  / xmc55_dps_xdec1_dummy_in
XDUMMY_OUT
+ VDD VSS  / xmc55_dps_xdec1_dummy_out
XDUM<1>
+ VDD VSS  / xmc55_dps_xdec1_dummy
XXDEC<63>
+ PXAA<3> PXAA<2> PXAA<1> PXAA<0> PXAB<3> PXAB<2> PXAB<1> PXAB<0> PXBA_N<7> 
+ PXBB_N<7> PXCA_N<7> PXCB_N<7> VDD VSS WLA<255> WLA<254> WLA<253> WLA<252> 
+ WLB<255> WLB<254> WLB<253> WLB<252>  / xmc55_dps_xdec4
XXDEC<62>
+ PXAA<3> PXAA<2> PXAA<1> PXAA<0> PXAB<3> PXAB<2> PXAB<1> PXAB<0> PXBA_N<6> 
+ PXBB_N<6> PXCA_N<7> PXCB_N<7> VDD VSS WLA<251> WLA<250> WLA<249> WLA<248> 
+ WLB<251> WLB<250> WLB<249> WLB<248>  / xmc55_dps_xdec4
XXDEC<61>
+ PXAA<3> PXAA<2> PXAA<1> PXAA<0> PXAB<3> PXAB<2> PXAB<1> PXAB<0> PXBA_N<5> 
+ PXBB_N<5> PXCA_N<7> PXCB_N<7> VDD VSS WLA<247> WLA<246> WLA<245> WLA<244> 
+ WLB<247> WLB<246> WLB<245> WLB<244>  / xmc55_dps_xdec4
XXDEC<60>
+ PXAA<3> PXAA<2> PXAA<1> PXAA<0> PXAB<3> PXAB<2> PXAB<1> PXAB<0> PXBA_N<4> 
+ PXBB_N<4> PXCA_N<7> PXCB_N<7> VDD VSS WLA<243> WLA<242> WLA<241> WLA<240> 
+ WLB<243> WLB<242> WLB<241> WLB<240>  / xmc55_dps_xdec4
XXDEC<59>
+ PXAA<3> PXAA<2> PXAA<1> PXAA<0> PXAB<3> PXAB<2> PXAB<1> PXAB<0> PXBA_N<3> 
+ PXBB_N<3> PXCA_N<7> PXCB_N<7> VDD VSS WLA<239> WLA<238> WLA<237> WLA<236> 
+ WLB<239> WLB<238> WLB<237> WLB<236>  / xmc55_dps_xdec4
XXDEC<58>
+ PXAA<3> PXAA<2> PXAA<1> PXAA<0> PXAB<3> PXAB<2> PXAB<1> PXAB<0> PXBA_N<2> 
+ PXBB_N<2> PXCA_N<7> PXCB_N<7> VDD VSS WLA<235> WLA<234> WLA<233> WLA<232> 
+ WLB<235> WLB<234> WLB<233> WLB<232>  / xmc55_dps_xdec4
XXDEC<57>
+ PXAA<3> PXAA<2> PXAA<1> PXAA<0> PXAB<3> PXAB<2> PXAB<1> PXAB<0> PXBA_N<1> 
+ PXBB_N<1> PXCA_N<7> PXCB_N<7> VDD VSS WLA<231> WLA<230> WLA<229> WLA<228> 
+ WLB<231> WLB<230> WLB<229> WLB<228>  / xmc55_dps_xdec4
XXDEC<56>
+ PXAA<3> PXAA<2> PXAA<1> PXAA<0> PXAB<3> PXAB<2> PXAB<1> PXAB<0> PXBA_N<0> 
+ PXBB_N<0> PXCA_N<7> PXCB_N<7> VDD VSS WLA<227> WLA<226> WLA<225> WLA<224> 
+ WLB<227> WLB<226> WLB<225> WLB<224>  / xmc55_dps_xdec4
XXDEC<55>
+ PXAA<3> PXAA<2> PXAA<1> PXAA<0> PXAB<3> PXAB<2> PXAB<1> PXAB<0> PXBA_N<7> 
+ PXBB_N<7> PXCA_N<6> PXCB_N<6> VDD VSS WLA<223> WLA<222> WLA<221> WLA<220> 
+ WLB<223> WLB<222> WLB<221> WLB<220>  / xmc55_dps_xdec4
XXDEC<54>
+ PXAA<3> PXAA<2> PXAA<1> PXAA<0> PXAB<3> PXAB<2> PXAB<1> PXAB<0> PXBA_N<6> 
+ PXBB_N<6> PXCA_N<6> PXCB_N<6> VDD VSS WLA<219> WLA<218> WLA<217> WLA<216> 
+ WLB<219> WLB<218> WLB<217> WLB<216>  / xmc55_dps_xdec4
XXDEC<53>
+ PXAA<3> PXAA<2> PXAA<1> PXAA<0> PXAB<3> PXAB<2> PXAB<1> PXAB<0> PXBA_N<5> 
+ PXBB_N<5> PXCA_N<6> PXCB_N<6> VDD VSS WLA<215> WLA<214> WLA<213> WLA<212> 
+ WLB<215> WLB<214> WLB<213> WLB<212>  / xmc55_dps_xdec4
XXDEC<52>
+ PXAA<3> PXAA<2> PXAA<1> PXAA<0> PXAB<3> PXAB<2> PXAB<1> PXAB<0> PXBA_N<4> 
+ PXBB_N<4> PXCA_N<6> PXCB_N<6> VDD VSS WLA<211> WLA<210> WLA<209> WLA<208> 
+ WLB<211> WLB<210> WLB<209> WLB<208>  / xmc55_dps_xdec4
XXDEC<51>
+ PXAA<3> PXAA<2> PXAA<1> PXAA<0> PXAB<3> PXAB<2> PXAB<1> PXAB<0> PXBA_N<3> 
+ PXBB_N<3> PXCA_N<6> PXCB_N<6> VDD VSS WLA<207> WLA<206> WLA<205> WLA<204> 
+ WLB<207> WLB<206> WLB<205> WLB<204>  / xmc55_dps_xdec4
XXDEC<50>
+ PXAA<3> PXAA<2> PXAA<1> PXAA<0> PXAB<3> PXAB<2> PXAB<1> PXAB<0> PXBA_N<2> 
+ PXBB_N<2> PXCA_N<6> PXCB_N<6> VDD VSS WLA<203> WLA<202> WLA<201> WLA<200> 
+ WLB<203> WLB<202> WLB<201> WLB<200>  / xmc55_dps_xdec4
XXDEC<49>
+ PXAA<3> PXAA<2> PXAA<1> PXAA<0> PXAB<3> PXAB<2> PXAB<1> PXAB<0> PXBA_N<1> 
+ PXBB_N<1> PXCA_N<6> PXCB_N<6> VDD VSS WLA<199> WLA<198> WLA<197> WLA<196> 
+ WLB<199> WLB<198> WLB<197> WLB<196>  / xmc55_dps_xdec4
XXDEC<48>
+ PXAA<3> PXAA<2> PXAA<1> PXAA<0> PXAB<3> PXAB<2> PXAB<1> PXAB<0> PXBA_N<0> 
+ PXBB_N<0> PXCA_N<6> PXCB_N<6> VDD VSS WLA<195> WLA<194> WLA<193> WLA<192> 
+ WLB<195> WLB<194> WLB<193> WLB<192>  / xmc55_dps_xdec4
XXDEC<47>
+ PXAA<3> PXAA<2> PXAA<1> PXAA<0> PXAB<3> PXAB<2> PXAB<1> PXAB<0> PXBA_N<7> 
+ PXBB_N<7> PXCA_N<5> PXCB_N<5> VDD VSS WLA<191> WLA<190> WLA<189> WLA<188> 
+ WLB<191> WLB<190> WLB<189> WLB<188>  / xmc55_dps_xdec4
XXDEC<46>
+ PXAA<3> PXAA<2> PXAA<1> PXAA<0> PXAB<3> PXAB<2> PXAB<1> PXAB<0> PXBA_N<6> 
+ PXBB_N<6> PXCA_N<5> PXCB_N<5> VDD VSS WLA<187> WLA<186> WLA<185> WLA<184> 
+ WLB<187> WLB<186> WLB<185> WLB<184>  / xmc55_dps_xdec4
XXDEC<45>
+ PXAA<3> PXAA<2> PXAA<1> PXAA<0> PXAB<3> PXAB<2> PXAB<1> PXAB<0> PXBA_N<5> 
+ PXBB_N<5> PXCA_N<5> PXCB_N<5> VDD VSS WLA<183> WLA<182> WLA<181> WLA<180> 
+ WLB<183> WLB<182> WLB<181> WLB<180>  / xmc55_dps_xdec4
XXDEC<44>
+ PXAA<3> PXAA<2> PXAA<1> PXAA<0> PXAB<3> PXAB<2> PXAB<1> PXAB<0> PXBA_N<4> 
+ PXBB_N<4> PXCA_N<5> PXCB_N<5> VDD VSS WLA<179> WLA<178> WLA<177> WLA<176> 
+ WLB<179> WLB<178> WLB<177> WLB<176>  / xmc55_dps_xdec4
XXDEC<43>
+ PXAA<3> PXAA<2> PXAA<1> PXAA<0> PXAB<3> PXAB<2> PXAB<1> PXAB<0> PXBA_N<3> 
+ PXBB_N<3> PXCA_N<5> PXCB_N<5> VDD VSS WLA<175> WLA<174> WLA<173> WLA<172> 
+ WLB<175> WLB<174> WLB<173> WLB<172>  / xmc55_dps_xdec4
XXDEC<42>
+ PXAA<3> PXAA<2> PXAA<1> PXAA<0> PXAB<3> PXAB<2> PXAB<1> PXAB<0> PXBA_N<2> 
+ PXBB_N<2> PXCA_N<5> PXCB_N<5> VDD VSS WLA<171> WLA<170> WLA<169> WLA<168> 
+ WLB<171> WLB<170> WLB<169> WLB<168>  / xmc55_dps_xdec4
XXDEC<41>
+ PXAA<3> PXAA<2> PXAA<1> PXAA<0> PXAB<3> PXAB<2> PXAB<1> PXAB<0> PXBA_N<1> 
+ PXBB_N<1> PXCA_N<5> PXCB_N<5> VDD VSS WLA<167> WLA<166> WLA<165> WLA<164> 
+ WLB<167> WLB<166> WLB<165> WLB<164>  / xmc55_dps_xdec4
XXDEC<40>
+ PXAA<3> PXAA<2> PXAA<1> PXAA<0> PXAB<3> PXAB<2> PXAB<1> PXAB<0> PXBA_N<0> 
+ PXBB_N<0> PXCA_N<5> PXCB_N<5> VDD VSS WLA<163> WLA<162> WLA<161> WLA<160> 
+ WLB<163> WLB<162> WLB<161> WLB<160>  / xmc55_dps_xdec4
XXDEC<39>
+ PXAA<3> PXAA<2> PXAA<1> PXAA<0> PXAB<3> PXAB<2> PXAB<1> PXAB<0> PXBA_N<7> 
+ PXBB_N<7> PXCA_N<4> PXCB_N<4> VDD VSS WLA<159> WLA<158> WLA<157> WLA<156> 
+ WLB<159> WLB<158> WLB<157> WLB<156>  / xmc55_dps_xdec4
XXDEC<38>
+ PXAA<3> PXAA<2> PXAA<1> PXAA<0> PXAB<3> PXAB<2> PXAB<1> PXAB<0> PXBA_N<6> 
+ PXBB_N<6> PXCA_N<4> PXCB_N<4> VDD VSS WLA<155> WLA<154> WLA<153> WLA<152> 
+ WLB<155> WLB<154> WLB<153> WLB<152>  / xmc55_dps_xdec4
XXDEC<37>
+ PXAA<3> PXAA<2> PXAA<1> PXAA<0> PXAB<3> PXAB<2> PXAB<1> PXAB<0> PXBA_N<5> 
+ PXBB_N<5> PXCA_N<4> PXCB_N<4> VDD VSS WLA<151> WLA<150> WLA<149> WLA<148> 
+ WLB<151> WLB<150> WLB<149> WLB<148>  / xmc55_dps_xdec4
XXDEC<36>
+ PXAA<3> PXAA<2> PXAA<1> PXAA<0> PXAB<3> PXAB<2> PXAB<1> PXAB<0> PXBA_N<4> 
+ PXBB_N<4> PXCA_N<4> PXCB_N<4> VDD VSS WLA<147> WLA<146> WLA<145> WLA<144> 
+ WLB<147> WLB<146> WLB<145> WLB<144>  / xmc55_dps_xdec4
XXDEC<35>
+ PXAA<3> PXAA<2> PXAA<1> PXAA<0> PXAB<3> PXAB<2> PXAB<1> PXAB<0> PXBA_N<3> 
+ PXBB_N<3> PXCA_N<4> PXCB_N<4> VDD VSS WLA<143> WLA<142> WLA<141> WLA<140> 
+ WLB<143> WLB<142> WLB<141> WLB<140>  / xmc55_dps_xdec4
XXDEC<34>
+ PXAA<3> PXAA<2> PXAA<1> PXAA<0> PXAB<3> PXAB<2> PXAB<1> PXAB<0> PXBA_N<2> 
+ PXBB_N<2> PXCA_N<4> PXCB_N<4> VDD VSS WLA<139> WLA<138> WLA<137> WLA<136> 
+ WLB<139> WLB<138> WLB<137> WLB<136>  / xmc55_dps_xdec4
XXDEC<33>
+ PXAA<3> PXAA<2> PXAA<1> PXAA<0> PXAB<3> PXAB<2> PXAB<1> PXAB<0> PXBA_N<1> 
+ PXBB_N<1> PXCA_N<4> PXCB_N<4> VDD VSS WLA<135> WLA<134> WLA<133> WLA<132> 
+ WLB<135> WLB<134> WLB<133> WLB<132>  / xmc55_dps_xdec4
XXDEC<32>
+ PXAA<3> PXAA<2> PXAA<1> PXAA<0> PXAB<3> PXAB<2> PXAB<1> PXAB<0> PXBA_N<0> 
+ PXBB_N<0> PXCA_N<4> PXCB_N<4> VDD VSS WLA<131> WLA<130> WLA<129> WLA<128> 
+ WLB<131> WLB<130> WLB<129> WLB<128>  / xmc55_dps_xdec4
XXDEC<31>
+ PXAA<3> PXAA<2> PXAA<1> PXAA<0> PXAB<3> PXAB<2> PXAB<1> PXAB<0> PXBA_N<7> 
+ PXBB_N<7> PXCA_N<3> PXCB_N<3> VDD VSS WLA<127> WLA<126> WLA<125> WLA<124> 
+ WLB<127> WLB<126> WLB<125> WLB<124>  / xmc55_dps_xdec4
XXDEC<30>
+ PXAA<3> PXAA<2> PXAA<1> PXAA<0> PXAB<3> PXAB<2> PXAB<1> PXAB<0> PXBA_N<6> 
+ PXBB_N<6> PXCA_N<3> PXCB_N<3> VDD VSS WLA<123> WLA<122> WLA<121> WLA<120> 
+ WLB<123> WLB<122> WLB<121> WLB<120>  / xmc55_dps_xdec4
XXDEC<29>
+ PXAA<3> PXAA<2> PXAA<1> PXAA<0> PXAB<3> PXAB<2> PXAB<1> PXAB<0> PXBA_N<5> 
+ PXBB_N<5> PXCA_N<3> PXCB_N<3> VDD VSS WLA<119> WLA<118> WLA<117> WLA<116> 
+ WLB<119> WLB<118> WLB<117> WLB<116>  / xmc55_dps_xdec4
XXDEC<28>
+ PXAA<3> PXAA<2> PXAA<1> PXAA<0> PXAB<3> PXAB<2> PXAB<1> PXAB<0> PXBA_N<4> 
+ PXBB_N<4> PXCA_N<3> PXCB_N<3> VDD VSS WLA<115> WLA<114> WLA<113> WLA<112> 
+ WLB<115> WLB<114> WLB<113> WLB<112>  / xmc55_dps_xdec4
XXDEC<27>
+ PXAA<3> PXAA<2> PXAA<1> PXAA<0> PXAB<3> PXAB<2> PXAB<1> PXAB<0> PXBA_N<3> 
+ PXBB_N<3> PXCA_N<3> PXCB_N<3> VDD VSS WLA<111> WLA<110> WLA<109> WLA<108> 
+ WLB<111> WLB<110> WLB<109> WLB<108>  / xmc55_dps_xdec4
XXDEC<26>
+ PXAA<3> PXAA<2> PXAA<1> PXAA<0> PXAB<3> PXAB<2> PXAB<1> PXAB<0> PXBA_N<2> 
+ PXBB_N<2> PXCA_N<3> PXCB_N<3> VDD VSS WLA<107> WLA<106> WLA<105> WLA<104> 
+ WLB<107> WLB<106> WLB<105> WLB<104>  / xmc55_dps_xdec4
XXDEC<25>
+ PXAA<3> PXAA<2> PXAA<1> PXAA<0> PXAB<3> PXAB<2> PXAB<1> PXAB<0> PXBA_N<1> 
+ PXBB_N<1> PXCA_N<3> PXCB_N<3> VDD VSS WLA<103> WLA<102> WLA<101> WLA<100> 
+ WLB<103> WLB<102> WLB<101> WLB<100>  / xmc55_dps_xdec4
XXDEC<24>
+ PXAA<3> PXAA<2> PXAA<1> PXAA<0> PXAB<3> PXAB<2> PXAB<1> PXAB<0> PXBA_N<0> 
+ PXBB_N<0> PXCA_N<3> PXCB_N<3> VDD VSS WLA<99> WLA<98> WLA<97> WLA<96> 
+ WLB<99> WLB<98> WLB<97> WLB<96>  / xmc55_dps_xdec4
XXDEC<23>
+ PXAA<3> PXAA<2> PXAA<1> PXAA<0> PXAB<3> PXAB<2> PXAB<1> PXAB<0> PXBA_N<7> 
+ PXBB_N<7> PXCA_N<2> PXCB_N<2> VDD VSS WLA<95> WLA<94> WLA<93> WLA<92> 
+ WLB<95> WLB<94> WLB<93> WLB<92>  / xmc55_dps_xdec4
XXDEC<22>
+ PXAA<3> PXAA<2> PXAA<1> PXAA<0> PXAB<3> PXAB<2> PXAB<1> PXAB<0> PXBA_N<6> 
+ PXBB_N<6> PXCA_N<2> PXCB_N<2> VDD VSS WLA<91> WLA<90> WLA<89> WLA<88> 
+ WLB<91> WLB<90> WLB<89> WLB<88>  / xmc55_dps_xdec4
XXDEC<21>
+ PXAA<3> PXAA<2> PXAA<1> PXAA<0> PXAB<3> PXAB<2> PXAB<1> PXAB<0> PXBA_N<5> 
+ PXBB_N<5> PXCA_N<2> PXCB_N<2> VDD VSS WLA<87> WLA<86> WLA<85> WLA<84> 
+ WLB<87> WLB<86> WLB<85> WLB<84>  / xmc55_dps_xdec4
XXDEC<20>
+ PXAA<3> PXAA<2> PXAA<1> PXAA<0> PXAB<3> PXAB<2> PXAB<1> PXAB<0> PXBA_N<4> 
+ PXBB_N<4> PXCA_N<2> PXCB_N<2> VDD VSS WLA<83> WLA<82> WLA<81> WLA<80> 
+ WLB<83> WLB<82> WLB<81> WLB<80>  / xmc55_dps_xdec4
XXDEC<19>
+ PXAA<3> PXAA<2> PXAA<1> PXAA<0> PXAB<3> PXAB<2> PXAB<1> PXAB<0> PXBA_N<3> 
+ PXBB_N<3> PXCA_N<2> PXCB_N<2> VDD VSS WLA<79> WLA<78> WLA<77> WLA<76> 
+ WLB<79> WLB<78> WLB<77> WLB<76>  / xmc55_dps_xdec4
XXDEC<18>
+ PXAA<3> PXAA<2> PXAA<1> PXAA<0> PXAB<3> PXAB<2> PXAB<1> PXAB<0> PXBA_N<2> 
+ PXBB_N<2> PXCA_N<2> PXCB_N<2> VDD VSS WLA<75> WLA<74> WLA<73> WLA<72> 
+ WLB<75> WLB<74> WLB<73> WLB<72>  / xmc55_dps_xdec4
XXDEC<17>
+ PXAA<3> PXAA<2> PXAA<1> PXAA<0> PXAB<3> PXAB<2> PXAB<1> PXAB<0> PXBA_N<1> 
+ PXBB_N<1> PXCA_N<2> PXCB_N<2> VDD VSS WLA<71> WLA<70> WLA<69> WLA<68> 
+ WLB<71> WLB<70> WLB<69> WLB<68>  / xmc55_dps_xdec4
XXDEC<16>
+ PXAA<3> PXAA<2> PXAA<1> PXAA<0> PXAB<3> PXAB<2> PXAB<1> PXAB<0> PXBA_N<0> 
+ PXBB_N<0> PXCA_N<2> PXCB_N<2> VDD VSS WLA<67> WLA<66> WLA<65> WLA<64> 
+ WLB<67> WLB<66> WLB<65> WLB<64>  / xmc55_dps_xdec4
XXDEC<15>
+ PXAA<3> PXAA<2> PXAA<1> PXAA<0> PXAB<3> PXAB<2> PXAB<1> PXAB<0> PXBA_N<7> 
+ PXBB_N<7> PXCA_N<1> PXCB_N<1> VDD VSS WLA<63> WLA<62> WLA<61> WLA<60> 
+ WLB<63> WLB<62> WLB<61> WLB<60>  / xmc55_dps_xdec4
XXDEC<14>
+ PXAA<3> PXAA<2> PXAA<1> PXAA<0> PXAB<3> PXAB<2> PXAB<1> PXAB<0> PXBA_N<6> 
+ PXBB_N<6> PXCA_N<1> PXCB_N<1> VDD VSS WLA<59> WLA<58> WLA<57> WLA<56> 
+ WLB<59> WLB<58> WLB<57> WLB<56>  / xmc55_dps_xdec4
XXDEC<13>
+ PXAA<3> PXAA<2> PXAA<1> PXAA<0> PXAB<3> PXAB<2> PXAB<1> PXAB<0> PXBA_N<5> 
+ PXBB_N<5> PXCA_N<1> PXCB_N<1> VDD VSS WLA<55> WLA<54> WLA<53> WLA<52> 
+ WLB<55> WLB<54> WLB<53> WLB<52>  / xmc55_dps_xdec4
XXDEC<12>
+ PXAA<3> PXAA<2> PXAA<1> PXAA<0> PXAB<3> PXAB<2> PXAB<1> PXAB<0> PXBA_N<4> 
+ PXBB_N<4> PXCA_N<1> PXCB_N<1> VDD VSS WLA<51> WLA<50> WLA<49> WLA<48> 
+ WLB<51> WLB<50> WLB<49> WLB<48>  / xmc55_dps_xdec4
XXDEC<11>
+ PXAA<3> PXAA<2> PXAA<1> PXAA<0> PXAB<3> PXAB<2> PXAB<1> PXAB<0> PXBA_N<3> 
+ PXBB_N<3> PXCA_N<1> PXCB_N<1> VDD VSS WLA<47> WLA<46> WLA<45> WLA<44> 
+ WLB<47> WLB<46> WLB<45> WLB<44>  / xmc55_dps_xdec4
XXDEC<10>
+ PXAA<3> PXAA<2> PXAA<1> PXAA<0> PXAB<3> PXAB<2> PXAB<1> PXAB<0> PXBA_N<2> 
+ PXBB_N<2> PXCA_N<1> PXCB_N<1> VDD VSS WLA<43> WLA<42> WLA<41> WLA<40> 
+ WLB<43> WLB<42> WLB<41> WLB<40>  / xmc55_dps_xdec4
XXDEC<9>
+ PXAA<3> PXAA<2> PXAA<1> PXAA<0> PXAB<3> PXAB<2> PXAB<1> PXAB<0> PXBA_N<1> 
+ PXBB_N<1> PXCA_N<1> PXCB_N<1> VDD VSS WLA<39> WLA<38> WLA<37> WLA<36> 
+ WLB<39> WLB<38> WLB<37> WLB<36>  / xmc55_dps_xdec4
XXDEC<8>
+ PXAA<3> PXAA<2> PXAA<1> PXAA<0> PXAB<3> PXAB<2> PXAB<1> PXAB<0> PXBA_N<0> 
+ PXBB_N<0> PXCA_N<1> PXCB_N<1> VDD VSS WLA<35> WLA<34> WLA<33> WLA<32> 
+ WLB<35> WLB<34> WLB<33> WLB<32>  / xmc55_dps_xdec4
XXDEC<7>
+ PXAA<3> PXAA<2> PXAA<1> PXAA<0> PXAB<3> PXAB<2> PXAB<1> PXAB<0> PXBA_N<7> 
+ PXBB_N<7> PXCA_N<0> PXCB_N<0> VDD VSS WLA<31> WLA<30> WLA<29> WLA<28> 
+ WLB<31> WLB<30> WLB<29> WLB<28>  / xmc55_dps_xdec4
XXDEC<6>
+ PXAA<3> PXAA<2> PXAA<1> PXAA<0> PXAB<3> PXAB<2> PXAB<1> PXAB<0> PXBA_N<6> 
+ PXBB_N<6> PXCA_N<0> PXCB_N<0> VDD VSS WLA<27> WLA<26> WLA<25> WLA<24> 
+ WLB<27> WLB<26> WLB<25> WLB<24>  / xmc55_dps_xdec4
XXDEC<5>
+ PXAA<3> PXAA<2> PXAA<1> PXAA<0> PXAB<3> PXAB<2> PXAB<1> PXAB<0> PXBA_N<5> 
+ PXBB_N<5> PXCA_N<0> PXCB_N<0> VDD VSS WLA<23> WLA<22> WLA<21> WLA<20> 
+ WLB<23> WLB<22> WLB<21> WLB<20>  / xmc55_dps_xdec4
XXDEC<4>
+ PXAA<3> PXAA<2> PXAA<1> PXAA<0> PXAB<3> PXAB<2> PXAB<1> PXAB<0> PXBA_N<4> 
+ PXBB_N<4> PXCA_N<0> PXCB_N<0> VDD VSS WLA<19> WLA<18> WLA<17> WLA<16> 
+ WLB<19> WLB<18> WLB<17> WLB<16>  / xmc55_dps_xdec4
XXDEC<3>
+ PXAA<3> PXAA<2> PXAA<1> PXAA<0> PXAB<3> PXAB<2> PXAB<1> PXAB<0> PXBA_N<3> 
+ PXBB_N<3> PXCA_N<0> PXCB_N<0> VDD VSS WLA<15> WLA<14> WLA<13> WLA<12> 
+ WLB<15> WLB<14> WLB<13> WLB<12>  / xmc55_dps_xdec4
XXDEC<2>
+ PXAA<3> PXAA<2> PXAA<1> PXAA<0> PXAB<3> PXAB<2> PXAB<1> PXAB<0> PXBA_N<2> 
+ PXBB_N<2> PXCA_N<0> PXCB_N<0> VDD VSS WLA<11> WLA<10> WLA<9> WLA<8> 
+ WLB<11> WLB<10> WLB<9> WLB<8>  / xmc55_dps_xdec4
XXDEC<1>
+ PXAA<3> PXAA<2> PXAA<1> PXAA<0> PXAB<3> PXAB<2> PXAB<1> PXAB<0> PXBA_N<1> 
+ PXBB_N<1> PXCA_N<0> PXCB_N<0> VDD VSS WLA<7> WLA<6> WLA<5> WLA<4> 
+ WLB<7> WLB<6> WLB<5> WLB<4>  / xmc55_dps_xdec4
XXDEC<0>
+ PXAA<3> PXAA<2> PXAA<1> PXAA<0> PXAB<3> PXAB<2> PXAB<1> PXAB<0> PXBA_N<0> 
+ PXBB_N<0> PXCA_N<0> PXCB_N<0> VDD VSS WLA<3> WLA<2> WLA<1> WLA<0> 
+ WLB<3> WLB<2> WLB<1> WLB<0>  / xmc55_dps_xdec4
.ENDS

************************************************************************
* Cell Name:    dpram16x4096_MIDX8_ROWX256
* View Name:    schematic
************************************************************************
.SUBCKT dpram16x4096_MIDX8_ROWX256
+ AA<12> AA<11> AA<10> AA<9> AA<8> AA<7> AA<6> AA<5> AA<4> 
+ AA<3> AA<2> AA<1> AA<0> AB<12> AB<11> AB<10> AB<9> AB<8> 
+ AB<7> AB<6> AB<5> AB<4> AB<3> AB<2> AB<1> AB<0> B_WLA<255> 
+ B_WLA<254> B_WLA<253> B_WLA<252> B_WLA<251> B_WLA<250> B_WLA<249> B_WLA<248> B_WLA<247> B_WLA<246> 
+ B_WLA<245> B_WLA<244> B_WLA<243> B_WLA<242> B_WLA<241> B_WLA<240> B_WLA<239> B_WLA<238> B_WLA<237> 
+ B_WLA<236> B_WLA<235> B_WLA<234> B_WLA<233> B_WLA<232> B_WLA<231> B_WLA<230> B_WLA<229> B_WLA<228> 
+ B_WLA<227> B_WLA<226> B_WLA<225> B_WLA<224> B_WLA<223> B_WLA<222> B_WLA<221> B_WLA<220> B_WLA<219> 
+ B_WLA<218> B_WLA<217> B_WLA<216> B_WLA<215> B_WLA<214> B_WLA<213> B_WLA<212> B_WLA<211> B_WLA<210> 
+ B_WLA<209> B_WLA<208> B_WLA<207> B_WLA<206> B_WLA<205> B_WLA<204> B_WLA<203> B_WLA<202> B_WLA<201> 
+ B_WLA<200> B_WLA<199> B_WLA<198> B_WLA<197> B_WLA<196> B_WLA<195> B_WLA<194> B_WLA<193> B_WLA<192> 
+ B_WLA<191> B_WLA<190> B_WLA<189> B_WLA<188> B_WLA<187> B_WLA<186> B_WLA<185> B_WLA<184> B_WLA<183> 
+ B_WLA<182> B_WLA<181> B_WLA<180> B_WLA<179> B_WLA<178> B_WLA<177> B_WLA<176> B_WLA<175> B_WLA<174> 
+ B_WLA<173> B_WLA<172> B_WLA<171> B_WLA<170> B_WLA<169> B_WLA<168> B_WLA<167> B_WLA<166> B_WLA<165> 
+ B_WLA<164> B_WLA<163> B_WLA<162> B_WLA<161> B_WLA<160> B_WLA<159> B_WLA<158> B_WLA<157> B_WLA<156> 
+ B_WLA<155> B_WLA<154> B_WLA<153> B_WLA<152> B_WLA<151> B_WLA<150> B_WLA<149> B_WLA<148> B_WLA<147> 
+ B_WLA<146> B_WLA<145> B_WLA<144> B_WLA<143> B_WLA<142> B_WLA<141> B_WLA<140> B_WLA<139> B_WLA<138> 
+ B_WLA<137> B_WLA<136> B_WLA<135> B_WLA<134> B_WLA<133> B_WLA<132> B_WLA<131> B_WLA<130> B_WLA<129> 
+ B_WLA<128> B_WLA<127> B_WLA<126> B_WLA<125> B_WLA<124> B_WLA<123> B_WLA<122> B_WLA<121> B_WLA<120> 
+ B_WLA<119> B_WLA<118> B_WLA<117> B_WLA<116> B_WLA<115> B_WLA<114> B_WLA<113> B_WLA<112> B_WLA<111> 
+ B_WLA<110> B_WLA<109> B_WLA<108> B_WLA<107> B_WLA<106> B_WLA<105> B_WLA<104> B_WLA<103> B_WLA<102> 
+ B_WLA<101> B_WLA<100> B_WLA<99> B_WLA<98> B_WLA<97> B_WLA<96> B_WLA<95> B_WLA<94> B_WLA<93> 
+ B_WLA<92> B_WLA<91> B_WLA<90> B_WLA<89> B_WLA<88> B_WLA<87> B_WLA<86> B_WLA<85> B_WLA<84> 
+ B_WLA<83> B_WLA<82> B_WLA<81> B_WLA<80> B_WLA<79> B_WLA<78> B_WLA<77> B_WLA<76> B_WLA<75> 
+ B_WLA<74> B_WLA<73> B_WLA<72> B_WLA<71> B_WLA<70> B_WLA<69> B_WLA<68> B_WLA<67> B_WLA<66> 
+ B_WLA<65> B_WLA<64> B_WLA<63> B_WLA<62> B_WLA<61> B_WLA<60> B_WLA<59> B_WLA<58> B_WLA<57> 
+ B_WLA<56> B_WLA<55> B_WLA<54> B_WLA<53> B_WLA<52> B_WLA<51> B_WLA<50> B_WLA<49> B_WLA<48> 
+ B_WLA<47> B_WLA<46> B_WLA<45> B_WLA<44> B_WLA<43> B_WLA<42> B_WLA<41> B_WLA<40> B_WLA<39> 
+ B_WLA<38> B_WLA<37> B_WLA<36> B_WLA<35> B_WLA<34> B_WLA<33> B_WLA<32> B_WLA<31> B_WLA<30> 
+ B_WLA<29> B_WLA<28> B_WLA<27> B_WLA<26> B_WLA<25> B_WLA<24> B_WLA<23> B_WLA<22> B_WLA<21> 
+ B_WLA<20> B_WLA<19> B_WLA<18> B_WLA<17> B_WLA<16> B_WLA<15> B_WLA<14> B_WLA<13> B_WLA<12> 
+ B_WLA<11> B_WLA<10> B_WLA<9> B_WLA<8> B_WLA<7> B_WLA<6> B_WLA<5> B_WLA<4> B_WLA<3> 
+ B_WLA<2> B_WLA<1> B_WLA<0> B_WLB<255> B_WLB<254> B_WLB<253> B_WLB<252> B_WLB<251> B_WLB<250> 
+ B_WLB<249> B_WLB<248> B_WLB<247> B_WLB<246> B_WLB<245> B_WLB<244> B_WLB<243> B_WLB<242> B_WLB<241> 
+ B_WLB<240> B_WLB<239> B_WLB<238> B_WLB<237> B_WLB<236> B_WLB<235> B_WLB<234> B_WLB<233> B_WLB<232> 
+ B_WLB<231> B_WLB<230> B_WLB<229> B_WLB<228> B_WLB<227> B_WLB<226> B_WLB<225> B_WLB<224> B_WLB<223> 
+ B_WLB<222> B_WLB<221> B_WLB<220> B_WLB<219> B_WLB<218> B_WLB<217> B_WLB<216> B_WLB<215> B_WLB<214> 
+ B_WLB<213> B_WLB<212> B_WLB<211> B_WLB<210> B_WLB<209> B_WLB<208> B_WLB<207> B_WLB<206> B_WLB<205> 
+ B_WLB<204> B_WLB<203> B_WLB<202> B_WLB<201> B_WLB<200> B_WLB<199> B_WLB<198> B_WLB<197> B_WLB<196> 
+ B_WLB<195> B_WLB<194> B_WLB<193> B_WLB<192> B_WLB<191> B_WLB<190> B_WLB<189> B_WLB<188> B_WLB<187> 
+ B_WLB<186> B_WLB<185> B_WLB<184> B_WLB<183> B_WLB<182> B_WLB<181> B_WLB<180> B_WLB<179> B_WLB<178> 
+ B_WLB<177> B_WLB<176> B_WLB<175> B_WLB<174> B_WLB<173> B_WLB<172> B_WLB<171> B_WLB<170> B_WLB<169> 
+ B_WLB<168> B_WLB<167> B_WLB<166> B_WLB<165> B_WLB<164> B_WLB<163> B_WLB<162> B_WLB<161> B_WLB<160> 
+ B_WLB<159> B_WLB<158> B_WLB<157> B_WLB<156> B_WLB<155> B_WLB<154> B_WLB<153> B_WLB<152> B_WLB<151> 
+ B_WLB<150> B_WLB<149> B_WLB<148> B_WLB<147> B_WLB<146> B_WLB<145> B_WLB<144> B_WLB<143> B_WLB<142> 
+ B_WLB<141> B_WLB<140> B_WLB<139> B_WLB<138> B_WLB<137> B_WLB<136> B_WLB<135> B_WLB<134> B_WLB<133> 
+ B_WLB<132> B_WLB<131> B_WLB<130> B_WLB<129> B_WLB<128> B_WLB<127> B_WLB<126> B_WLB<125> B_WLB<124> 
+ B_WLB<123> B_WLB<122> B_WLB<121> B_WLB<120> B_WLB<119> B_WLB<118> B_WLB<117> B_WLB<116> B_WLB<115> 
+ B_WLB<114> B_WLB<113> B_WLB<112> B_WLB<111> B_WLB<110> B_WLB<109> B_WLB<108> B_WLB<107> B_WLB<106> 
+ B_WLB<105> B_WLB<104> B_WLB<103> B_WLB<102> B_WLB<101> B_WLB<100> B_WLB<99> B_WLB<98> B_WLB<97> 
+ B_WLB<96> B_WLB<95> B_WLB<94> B_WLB<93> B_WLB<92> B_WLB<91> B_WLB<90> B_WLB<89> B_WLB<88> 
+ B_WLB<87> B_WLB<86> B_WLB<85> B_WLB<84> B_WLB<83> B_WLB<82> B_WLB<81> B_WLB<80> B_WLB<79> 
+ B_WLB<78> B_WLB<77> B_WLB<76> B_WLB<75> B_WLB<74> B_WLB<73> B_WLB<72> B_WLB<71> B_WLB<70> 
+ B_WLB<69> B_WLB<68> B_WLB<67> B_WLB<66> B_WLB<65> B_WLB<64> B_WLB<63> B_WLB<62> B_WLB<61> 
+ B_WLB<60> B_WLB<59> B_WLB<58> B_WLB<57> B_WLB<56> B_WLB<55> B_WLB<54> B_WLB<53> B_WLB<52> 
+ B_WLB<51> B_WLB<50> B_WLB<49> B_WLB<48> B_WLB<47> B_WLB<46> B_WLB<45> B_WLB<44> B_WLB<43> 
+ B_WLB<42> B_WLB<41> B_WLB<40> B_WLB<39> B_WLB<38> B_WLB<37> B_WLB<36> B_WLB<35> B_WLB<34> 
+ B_WLB<33> B_WLB<32> B_WLB<31> B_WLB<30> B_WLB<29> B_WLB<28> B_WLB<27> B_WLB<26> B_WLB<25> 
+ B_WLB<24> B_WLB<23> B_WLB<22> B_WLB<21> B_WLB<20> B_WLB<19> B_WLB<18> B_WLB<17> B_WLB<16> 
+ B_WLB<15> B_WLB<14> B_WLB<13> B_WLB<12> B_WLB<11> B_WLB<10> B_WLB<9> B_WLB<8> B_WLB<7> 
+ B_WLB<6> B_WLB<5> B_WLB<4> B_WLB<3> B_WLB<2> B_WLB<1> B_WLB<0> CENA CENB 
+ CLKA CLKB DBL_PD_N<3> DBL_PD_N<2> DBL_PD_N<1> DBL_PD_N<0> DDQA DDQA_N DDQB 
+ DDQB_N DWLA<1> DWLA<0> DWLB<1> DWLB<0> L_CLK_DQA L_CLK_DQA_N L_CLK_DQB L_CLK_DQB_N 
+ L_LWEA L_LWEB L_SA_PREA_N L_SA_PREB_N L_SAEA_N L_SAEB_N LB_CA<3> LB_CA<2> LB_CA<1> 
+ LB_CA<0> LB_CB<3> LB_CB<2> LB_CB<1> LB_CB<0> LB_MA<3> LB_MA<2> LB_MA<1> LB_MA<0> 
+ LB_MB<3> LB_MB<2> LB_MB<1> LB_MB<0> LB_TM_PREA_N LB_TM_PREB_N LT_CA<3> LT_CA<2> LT_CA<1> 
+ LT_CA<0> LT_CB<3> LT_CB<2> LT_CB<1> LT_CB<0> LT_MA<3> LT_MA<2> LT_MA<1> LT_MA<0> 
+ LT_MB<3> LT_MB<2> LT_MB<1> LT_MB<0> LT_TM_PREA_N LT_TM_PREB_N R_CLK_DQA R_CLK_DQA_N R_CLK_DQB 
+ R_CLK_DQB_N R_LWEA R_LWEB R_SA_PREA_N R_SA_PREB_N R_SAEA_N R_SAEB_N RB_CA<3> RB_CA<2> 
+ RB_CA<1> RB_CA<0> RB_CB<3> RB_CB<2> RB_CB<1> RB_CB<0> RB_MA<3> RB_MA<2> RB_MA<1> 
+ RB_MA<0> RB_MB<3> RB_MB<2> RB_MB<1> RB_MB<0> RB_TM_PREA_N RB_TM_PREB_N RT_CA<3> RT_CA<2> 
+ RT_CA<1> RT_CA<0> RT_CB<3> RT_CB<2> RT_CB<1> RT_CB<0> RT_MA<3> RT_MA<2> RT_MA<1> 
+ RT_MA<0> RT_MB<3> RT_MB<2> RT_MB<1> RT_MB<0> RT_TM_PREA_N RT_TM_PREB_N STCLKA STCLKB 
+ T_WLA<255> T_WLA<254> T_WLA<253> T_WLA<252> T_WLA<251> T_WLA<250> T_WLA<249> T_WLA<248> T_WLA<247> 
+ T_WLA<246> T_WLA<245> T_WLA<244> T_WLA<243> T_WLA<242> T_WLA<241> T_WLA<240> T_WLA<239> T_WLA<238> 
+ T_WLA<237> T_WLA<236> T_WLA<235> T_WLA<234> T_WLA<233> T_WLA<232> T_WLA<231> T_WLA<230> T_WLA<229> 
+ T_WLA<228> T_WLA<227> T_WLA<226> T_WLA<225> T_WLA<224> T_WLA<223> T_WLA<222> T_WLA<221> T_WLA<220> 
+ T_WLA<219> T_WLA<218> T_WLA<217> T_WLA<216> T_WLA<215> T_WLA<214> T_WLA<213> T_WLA<212> T_WLA<211> 
+ T_WLA<210> T_WLA<209> T_WLA<208> T_WLA<207> T_WLA<206> T_WLA<205> T_WLA<204> T_WLA<203> T_WLA<202> 
+ T_WLA<201> T_WLA<200> T_WLA<199> T_WLA<198> T_WLA<197> T_WLA<196> T_WLA<195> T_WLA<194> T_WLA<193> 
+ T_WLA<192> T_WLA<191> T_WLA<190> T_WLA<189> T_WLA<188> T_WLA<187> T_WLA<186> T_WLA<185> T_WLA<184> 
+ T_WLA<183> T_WLA<182> T_WLA<181> T_WLA<180> T_WLA<179> T_WLA<178> T_WLA<177> T_WLA<176> T_WLA<175> 
+ T_WLA<174> T_WLA<173> T_WLA<172> T_WLA<171> T_WLA<170> T_WLA<169> T_WLA<168> T_WLA<167> T_WLA<166> 
+ T_WLA<165> T_WLA<164> T_WLA<163> T_WLA<162> T_WLA<161> T_WLA<160> T_WLA<159> T_WLA<158> T_WLA<157> 
+ T_WLA<156> T_WLA<155> T_WLA<154> T_WLA<153> T_WLA<152> T_WLA<151> T_WLA<150> T_WLA<149> T_WLA<148> 
+ T_WLA<147> T_WLA<146> T_WLA<145> T_WLA<144> T_WLA<143> T_WLA<142> T_WLA<141> T_WLA<140> T_WLA<139> 
+ T_WLA<138> T_WLA<137> T_WLA<136> T_WLA<135> T_WLA<134> T_WLA<133> T_WLA<132> T_WLA<131> T_WLA<130> 
+ T_WLA<129> T_WLA<128> T_WLA<127> T_WLA<126> T_WLA<125> T_WLA<124> T_WLA<123> T_WLA<122> T_WLA<121> 
+ T_WLA<120> T_WLA<119> T_WLA<118> T_WLA<117> T_WLA<116> T_WLA<115> T_WLA<114> T_WLA<113> T_WLA<112> 
+ T_WLA<111> T_WLA<110> T_WLA<109> T_WLA<108> T_WLA<107> T_WLA<106> T_WLA<105> T_WLA<104> T_WLA<103> 
+ T_WLA<102> T_WLA<101> T_WLA<100> T_WLA<99> T_WLA<98> T_WLA<97> T_WLA<96> T_WLA<95> T_WLA<94> 
+ T_WLA<93> T_WLA<92> T_WLA<91> T_WLA<90> T_WLA<89> T_WLA<88> T_WLA<87> T_WLA<86> T_WLA<85> 
+ T_WLA<84> T_WLA<83> T_WLA<82> T_WLA<81> T_WLA<80> T_WLA<79> T_WLA<78> T_WLA<77> T_WLA<76> 
+ T_WLA<75> T_WLA<74> T_WLA<73> T_WLA<72> T_WLA<71> T_WLA<70> T_WLA<69> T_WLA<68> T_WLA<67> 
+ T_WLA<66> T_WLA<65> T_WLA<64> T_WLA<63> T_WLA<62> T_WLA<61> T_WLA<60> T_WLA<59> T_WLA<58> 
+ T_WLA<57> T_WLA<56> T_WLA<55> T_WLA<54> T_WLA<53> T_WLA<52> T_WLA<51> T_WLA<50> T_WLA<49> 
+ T_WLA<48> T_WLA<47> T_WLA<46> T_WLA<45> T_WLA<44> T_WLA<43> T_WLA<42> T_WLA<41> T_WLA<40> 
+ T_WLA<39> T_WLA<38> T_WLA<37> T_WLA<36> T_WLA<35> T_WLA<34> T_WLA<33> T_WLA<32> T_WLA<31> 
+ T_WLA<30> T_WLA<29> T_WLA<28> T_WLA<27> T_WLA<26> T_WLA<25> T_WLA<24> T_WLA<23> T_WLA<22> 
+ T_WLA<21> T_WLA<20> T_WLA<19> T_WLA<18> T_WLA<17> T_WLA<16> T_WLA<15> T_WLA<14> T_WLA<13> 
+ T_WLA<12> T_WLA<11> T_WLA<10> T_WLA<9> T_WLA<8> T_WLA<7> T_WLA<6> T_WLA<5> T_WLA<4> 
+ T_WLA<3> T_WLA<2> T_WLA<1> T_WLA<0> T_WLB<255> T_WLB<254> T_WLB<253> T_WLB<252> T_WLB<251> 
+ T_WLB<250> T_WLB<249> T_WLB<248> T_WLB<247> T_WLB<246> T_WLB<245> T_WLB<244> T_WLB<243> T_WLB<242> 
+ T_WLB<241> T_WLB<240> T_WLB<239> T_WLB<238> T_WLB<237> T_WLB<236> T_WLB<235> T_WLB<234> T_WLB<233> 
+ T_WLB<232> T_WLB<231> T_WLB<230> T_WLB<229> T_WLB<228> T_WLB<227> T_WLB<226> T_WLB<225> T_WLB<224> 
+ T_WLB<223> T_WLB<222> T_WLB<221> T_WLB<220> T_WLB<219> T_WLB<218> T_WLB<217> T_WLB<216> T_WLB<215> 
+ T_WLB<214> T_WLB<213> T_WLB<212> T_WLB<211> T_WLB<210> T_WLB<209> T_WLB<208> T_WLB<207> T_WLB<206> 
+ T_WLB<205> T_WLB<204> T_WLB<203> T_WLB<202> T_WLB<201> T_WLB<200> T_WLB<199> T_WLB<198> T_WLB<197> 
+ T_WLB<196> T_WLB<195> T_WLB<194> T_WLB<193> T_WLB<192> T_WLB<191> T_WLB<190> T_WLB<189> T_WLB<188> 
+ T_WLB<187> T_WLB<186> T_WLB<185> T_WLB<184> T_WLB<183> T_WLB<182> T_WLB<181> T_WLB<180> T_WLB<179> 
+ T_WLB<178> T_WLB<177> T_WLB<176> T_WLB<175> T_WLB<174> T_WLB<173> T_WLB<172> T_WLB<171> T_WLB<170> 
+ T_WLB<169> T_WLB<168> T_WLB<167> T_WLB<166> T_WLB<165> T_WLB<164> T_WLB<163> T_WLB<162> T_WLB<161> 
+ T_WLB<160> T_WLB<159> T_WLB<158> T_WLB<157> T_WLB<156> T_WLB<155> T_WLB<154> T_WLB<153> T_WLB<152> 
+ T_WLB<151> T_WLB<150> T_WLB<149> T_WLB<148> T_WLB<147> T_WLB<146> T_WLB<145> T_WLB<144> T_WLB<143> 
+ T_WLB<142> T_WLB<141> T_WLB<140> T_WLB<139> T_WLB<138> T_WLB<137> T_WLB<136> T_WLB<135> T_WLB<134> 
+ T_WLB<133> T_WLB<132> T_WLB<131> T_WLB<130> T_WLB<129> T_WLB<128> T_WLB<127> T_WLB<126> T_WLB<125> 
+ T_WLB<124> T_WLB<123> T_WLB<122> T_WLB<121> T_WLB<120> T_WLB<119> T_WLB<118> T_WLB<117> T_WLB<116> 
+ T_WLB<115> T_WLB<114> T_WLB<113> T_WLB<112> T_WLB<111> T_WLB<110> T_WLB<109> T_WLB<108> T_WLB<107> 
+ T_WLB<106> T_WLB<105> T_WLB<104> T_WLB<103> T_WLB<102> T_WLB<101> T_WLB<100> T_WLB<99> T_WLB<98> 
+ T_WLB<97> T_WLB<96> T_WLB<95> T_WLB<94> T_WLB<93> T_WLB<92> T_WLB<91> T_WLB<90> T_WLB<89> 
+ T_WLB<88> T_WLB<87> T_WLB<86> T_WLB<85> T_WLB<84> T_WLB<83> T_WLB<82> T_WLB<81> T_WLB<80> 
+ T_WLB<79> T_WLB<78> T_WLB<77> T_WLB<76> T_WLB<75> T_WLB<74> T_WLB<73> T_WLB<72> T_WLB<71> 
+ T_WLB<70> T_WLB<69> T_WLB<68> T_WLB<67> T_WLB<66> T_WLB<65> T_WLB<64> T_WLB<63> T_WLB<62> 
+ T_WLB<61> T_WLB<60> T_WLB<59> T_WLB<58> T_WLB<57> T_WLB<56> T_WLB<55> T_WLB<54> T_WLB<53> 
+ T_WLB<52> T_WLB<51> T_WLB<50> T_WLB<49> T_WLB<48> T_WLB<47> T_WLB<46> T_WLB<45> T_WLB<44> 
+ T_WLB<43> T_WLB<42> T_WLB<41> T_WLB<40> T_WLB<39> T_WLB<38> T_WLB<37> T_WLB<36> T_WLB<35> 
+ T_WLB<34> T_WLB<33> T_WLB<32> T_WLB<31> T_WLB<30> T_WLB<29> T_WLB<28> T_WLB<27> T_WLB<26> 
+ T_WLB<25> T_WLB<24> T_WLB<23> T_WLB<22> T_WLB<21> T_WLB<20> T_WLB<19> T_WLB<18> T_WLB<17> 
+ T_WLB<16> T_WLB<15> T_WLB<14> T_WLB<13> T_WLB<12> T_WLB<11> T_WLB<10> T_WLB<9> T_WLB<8> 
+ T_WLB<7> T_WLB<6> T_WLB<5> T_WLB<4> T_WLB<3> T_WLB<2> T_WLB<1> T_WLB<0> TIE_VDD 
+ TIE_VSS TM<9> TM<8> TM<7> TM<6> TM<5> TM<4> TM<3> TM<2> 
+ TM<1> TM<0> VDD VSS WENA WENB 
XXDEC_TOP
+ T_PXAA<3> T_PXAA<2> T_PXAA<1> T_PXAA<0> T_PXAB<3> T_PXAB<2> T_PXAB<1> T_PXAB<0> T_PXBA_N<7> 
+ T_PXBA_N<6> T_PXBA_N<5> T_PXBA_N<4> T_PXBA_N<3> T_PXBA_N<2> T_PXBA_N<1> T_PXBA_N<0> T_PXBB_N<7> T_PXBB_N<6> 
+ T_PXBB_N<5> T_PXBB_N<4> T_PXBB_N<3> T_PXBB_N<2> T_PXBB_N<1> T_PXBB_N<0> T_PXCA_N<7> T_PXCA_N<6> T_PXCA_N<5> 
+ T_PXCA_N<4> T_PXCA_N<3> T_PXCA_N<2> T_PXCA_N<1> T_PXCA_N<0> T_PXCB_N<7> T_PXCB_N<6> T_PXCB_N<5> T_PXCB_N<4> 
+ T_PXCB_N<3> T_PXCB_N<2> T_PXCB_N<1> T_PXCB_N<0> VDD VSS T_WLA<255> T_WLA<254> T_WLA<253> 
+ T_WLA<252> T_WLA<251> T_WLA<250> T_WLA<249> T_WLA<248> T_WLA<247> T_WLA<246> T_WLA<245> T_WLA<244> 
+ T_WLA<243> T_WLA<242> T_WLA<241> T_WLA<240> T_WLA<239> T_WLA<238> T_WLA<237> T_WLA<236> T_WLA<235> 
+ T_WLA<234> T_WLA<233> T_WLA<232> T_WLA<231> T_WLA<230> T_WLA<229> T_WLA<228> T_WLA<227> T_WLA<226> 
+ T_WLA<225> T_WLA<224> T_WLA<223> T_WLA<222> T_WLA<221> T_WLA<220> T_WLA<219> T_WLA<218> T_WLA<217> 
+ T_WLA<216> T_WLA<215> T_WLA<214> T_WLA<213> T_WLA<212> T_WLA<211> T_WLA<210> T_WLA<209> T_WLA<208> 
+ T_WLA<207> T_WLA<206> T_WLA<205> T_WLA<204> T_WLA<203> T_WLA<202> T_WLA<201> T_WLA<200> T_WLA<199> 
+ T_WLA<198> T_WLA<197> T_WLA<196> T_WLA<195> T_WLA<194> T_WLA<193> T_WLA<192> T_WLA<191> T_WLA<190> 
+ T_WLA<189> T_WLA<188> T_WLA<187> T_WLA<186> T_WLA<185> T_WLA<184> T_WLA<183> T_WLA<182> T_WLA<181> 
+ T_WLA<180> T_WLA<179> T_WLA<178> T_WLA<177> T_WLA<176> T_WLA<175> T_WLA<174> T_WLA<173> T_WLA<172> 
+ T_WLA<171> T_WLA<170> T_WLA<169> T_WLA<168> T_WLA<167> T_WLA<166> T_WLA<165> T_WLA<164> T_WLA<163> 
+ T_WLA<162> T_WLA<161> T_WLA<160> T_WLA<159> T_WLA<158> T_WLA<157> T_WLA<156> T_WLA<155> T_WLA<154> 
+ T_WLA<153> T_WLA<152> T_WLA<151> T_WLA<150> T_WLA<149> T_WLA<148> T_WLA<147> T_WLA<146> T_WLA<145> 
+ T_WLA<144> T_WLA<143> T_WLA<142> T_WLA<141> T_WLA<140> T_WLA<139> T_WLA<138> T_WLA<137> T_WLA<136> 
+ T_WLA<135> T_WLA<134> T_WLA<133> T_WLA<132> T_WLA<131> T_WLA<130> T_WLA<129> T_WLA<128> T_WLA<127> 
+ T_WLA<126> T_WLA<125> T_WLA<124> T_WLA<123> T_WLA<122> T_WLA<121> T_WLA<120> T_WLA<119> T_WLA<118> 
+ T_WLA<117> T_WLA<116> T_WLA<115> T_WLA<114> T_WLA<113> T_WLA<112> T_WLA<111> T_WLA<110> T_WLA<109> 
+ T_WLA<108> T_WLA<107> T_WLA<106> T_WLA<105> T_WLA<104> T_WLA<103> T_WLA<102> T_WLA<101> T_WLA<100> 
+ T_WLA<99> T_WLA<98> T_WLA<97> T_WLA<96> T_WLA<95> T_WLA<94> T_WLA<93> T_WLA<92> T_WLA<91> 
+ T_WLA<90> T_WLA<89> T_WLA<88> T_WLA<87> T_WLA<86> T_WLA<85> T_WLA<84> T_WLA<83> T_WLA<82> 
+ T_WLA<81> T_WLA<80> T_WLA<79> T_WLA<78> T_WLA<77> T_WLA<76> T_WLA<75> T_WLA<74> T_WLA<73> 
+ T_WLA<72> T_WLA<71> T_WLA<70> T_WLA<69> T_WLA<68> T_WLA<67> T_WLA<66> T_WLA<65> T_WLA<64> 
+ T_WLA<63> T_WLA<62> T_WLA<61> T_WLA<60> T_WLA<59> T_WLA<58> T_WLA<57> T_WLA<56> T_WLA<55> 
+ T_WLA<54> T_WLA<53> T_WLA<52> T_WLA<51> T_WLA<50> T_WLA<49> T_WLA<48> T_WLA<47> T_WLA<46> 
+ T_WLA<45> T_WLA<44> T_WLA<43> T_WLA<42> T_WLA<41> T_WLA<40> T_WLA<39> T_WLA<38> T_WLA<37> 
+ T_WLA<36> T_WLA<35> T_WLA<34> T_WLA<33> T_WLA<32> T_WLA<31> T_WLA<30> T_WLA<29> T_WLA<28> 
+ T_WLA<27> T_WLA<26> T_WLA<25> T_WLA<24> T_WLA<23> T_WLA<22> T_WLA<21> T_WLA<20> T_WLA<19> 
+ T_WLA<18> T_WLA<17> T_WLA<16> T_WLA<15> T_WLA<14> T_WLA<13> T_WLA<12> T_WLA<11> T_WLA<10> 
+ T_WLA<9> T_WLA<8> T_WLA<7> T_WLA<6> T_WLA<5> T_WLA<4> T_WLA<3> T_WLA<2> T_WLA<1> 
+ T_WLA<0> T_WLB<255> T_WLB<254> T_WLB<253> T_WLB<252> T_WLB<251> T_WLB<250> T_WLB<249> T_WLB<248> 
+ T_WLB<247> T_WLB<246> T_WLB<245> T_WLB<244> T_WLB<243> T_WLB<242> T_WLB<241> T_WLB<240> T_WLB<239> 
+ T_WLB<238> T_WLB<237> T_WLB<236> T_WLB<235> T_WLB<234> T_WLB<233> T_WLB<232> T_WLB<231> T_WLB<230> 
+ T_WLB<229> T_WLB<228> T_WLB<227> T_WLB<226> T_WLB<225> T_WLB<224> T_WLB<223> T_WLB<222> T_WLB<221> 
+ T_WLB<220> T_WLB<219> T_WLB<218> T_WLB<217> T_WLB<216> T_WLB<215> T_WLB<214> T_WLB<213> T_WLB<212> 
+ T_WLB<211> T_WLB<210> T_WLB<209> T_WLB<208> T_WLB<207> T_WLB<206> T_WLB<205> T_WLB<204> T_WLB<203> 
+ T_WLB<202> T_WLB<201> T_WLB<200> T_WLB<199> T_WLB<198> T_WLB<197> T_WLB<196> T_WLB<195> T_WLB<194> 
+ T_WLB<193> T_WLB<192> T_WLB<191> T_WLB<190> T_WLB<189> T_WLB<188> T_WLB<187> T_WLB<186> T_WLB<185> 
+ T_WLB<184> T_WLB<183> T_WLB<182> T_WLB<181> T_WLB<180> T_WLB<179> T_WLB<178> T_WLB<177> T_WLB<176> 
+ T_WLB<175> T_WLB<174> T_WLB<173> T_WLB<172> T_WLB<171> T_WLB<170> T_WLB<169> T_WLB<168> T_WLB<167> 
+ T_WLB<166> T_WLB<165> T_WLB<164> T_WLB<163> T_WLB<162> T_WLB<161> T_WLB<160> T_WLB<159> T_WLB<158> 
+ T_WLB<157> T_WLB<156> T_WLB<155> T_WLB<154> T_WLB<153> T_WLB<152> T_WLB<151> T_WLB<150> T_WLB<149> 
+ T_WLB<148> T_WLB<147> T_WLB<146> T_WLB<145> T_WLB<144> T_WLB<143> T_WLB<142> T_WLB<141> T_WLB<140> 
+ T_WLB<139> T_WLB<138> T_WLB<137> T_WLB<136> T_WLB<135> T_WLB<134> T_WLB<133> T_WLB<132> T_WLB<131> 
+ T_WLB<130> T_WLB<129> T_WLB<128> T_WLB<127> T_WLB<126> T_WLB<125> T_WLB<124> T_WLB<123> T_WLB<122> 
+ T_WLB<121> T_WLB<120> T_WLB<119> T_WLB<118> T_WLB<117> T_WLB<116> T_WLB<115> T_WLB<114> T_WLB<113> 
+ T_WLB<112> T_WLB<111> T_WLB<110> T_WLB<109> T_WLB<108> T_WLB<107> T_WLB<106> T_WLB<105> T_WLB<104> 
+ T_WLB<103> T_WLB<102> T_WLB<101> T_WLB<100> T_WLB<99> T_WLB<98> T_WLB<97> T_WLB<96> T_WLB<95> 
+ T_WLB<94> T_WLB<93> T_WLB<92> T_WLB<91> T_WLB<90> T_WLB<89> T_WLB<88> T_WLB<87> T_WLB<86> 
+ T_WLB<85> T_WLB<84> T_WLB<83> T_WLB<82> T_WLB<81> T_WLB<80> T_WLB<79> T_WLB<78> T_WLB<77> 
+ T_WLB<76> T_WLB<75> T_WLB<74> T_WLB<73> T_WLB<72> T_WLB<71> T_WLB<70> T_WLB<69> T_WLB<68> 
+ T_WLB<67> T_WLB<66> T_WLB<65> T_WLB<64> T_WLB<63> T_WLB<62> T_WLB<61> T_WLB<60> T_WLB<59> 
+ T_WLB<58> T_WLB<57> T_WLB<56> T_WLB<55> T_WLB<54> T_WLB<53> T_WLB<52> T_WLB<51> T_WLB<50> 
+ T_WLB<49> T_WLB<48> T_WLB<47> T_WLB<46> T_WLB<45> T_WLB<44> T_WLB<43> T_WLB<42> T_WLB<41> 
+ T_WLB<40> T_WLB<39> T_WLB<38> T_WLB<37> T_WLB<36> T_WLB<35> T_WLB<34> T_WLB<33> T_WLB<32> 
+ T_WLB<31> T_WLB<30> T_WLB<29> T_WLB<28> T_WLB<27> T_WLB<26> T_WLB<25> T_WLB<24> T_WLB<23> 
+ T_WLB<22> T_WLB<21> T_WLB<20> T_WLB<19> T_WLB<18> T_WLB<17> T_WLB<16> T_WLB<15> T_WLB<14> 
+ T_WLB<13> T_WLB<12> T_WLB<11> T_WLB<10> T_WLB<9> T_WLB<8> T_WLB<7> T_WLB<6> T_WLB<5> 
+ T_WLB<4> T_WLB<3> T_WLB<2> T_WLB<1> T_WLB<0>  / dpram16x4096_XDECX256
XCTRL
+ NET133<12> NET133<11> NET133<10> NET133<9> NET133<8> NET133<7> NET133<6> NET133<5> NET133<4> 
+ NET133<3> NET133<2> NET133<1> NET133<0> NET131<12> NET131<11> NET131<10> NET131<9> NET131<8> 
+ NET131<7> NET131<6> NET131<5> NET131<4> NET131<3> NET131<2> NET131<1> NET131<0> B_PXAA<3> 
+ B_PXAA<2> B_PXAA<1> B_PXAA<0> B_PXAB<3> B_PXAB<2> B_PXAB<1> B_PXAB<0> B_PXBA_N<7> B_PXBA_N<6> 
+ B_PXBA_N<5> B_PXBA_N<4> B_PXBA_N<3> B_PXBA_N<2> B_PXBA_N<1> B_PXBA_N<0> B_PXBB_N<7> B_PXBB_N<6> B_PXBB_N<5> 
+ B_PXBB_N<4> B_PXBB_N<3> B_PXBB_N<2> B_PXBB_N<1> B_PXBB_N<0> B_PXCA_N<7> B_PXCA_N<6> B_PXCA_N<5> B_PXCA_N<4> 
+ B_PXCA_N<3> B_PXCA_N<2> B_PXCA_N<1> B_PXCA_N<0> B_PXCB_N<7> B_PXCB_N<6> B_PXCB_N<5> B_PXCB_N<4> B_PXCB_N<3> 
+ B_PXCB_N<2> B_PXCB_N<1> B_PXCB_N<0> NET122 NET121 NET125 NET127 DBL_PD_N<3> DBL_PD_N<2> 
+ DBL_PD_N<1> DBL_PD_N<0> DDQA DDQA_N DDQB DDQB_N DWLA<1> DWLA<0> DWLB<1> 
+ DWLB<0> L_CLK_DQA L_CLK_DQA_N L_CLK_DQB L_CLK_DQB_N L_LWEA L_LWEB L_SA_PREA_N L_SA_PREB_N 
+ L_SAEA_N L_SAEB_N LB_CA<3> LB_CA<2> LB_CA<1> LB_CA<0> LB_CB<3> LB_CB<2> LB_CB<1> 
+ LB_CB<0> LB_MA<3> LB_MA<2> LB_MA<1> LB_MA<0> LB_MB<3> LB_MB<2> LB_MB<1> LB_MB<0> 
+ LB_TM_PREA_N LB_TM_PREB_N LT_CA<3> LT_CA<2> LT_CA<1> LT_CA<0> LT_CB<3> LT_CB<2> LT_CB<1> 
+ LT_CB<0> LT_MA<3> LT_MA<2> LT_MA<1> LT_MA<0> LT_MB<3> LT_MB<2> LT_MB<1> LT_MB<0> 
+ LT_TM_PREA_N LT_TM_PREB_N R_CLK_DQA R_CLK_DQA_N R_CLK_DQB R_CLK_DQB_N R_LWEA R_LWEB R_SA_PREA_N 
+ R_SA_PREB_N R_SAEA_N R_SAEB_N RB_CA<3> RB_CA<2> RB_CA<1> RB_CA<0> RB_CB<3> RB_CB<2> 
+ RB_CB<1> RB_CB<0> RB_MA<3> RB_MA<2> RB_MA<1> RB_MA<0> RB_MB<3> RB_MB<2> RB_MB<1> 
+ RB_MB<0> RB_TM_PREA_N RB_TM_PREB_N RT_CA<3> RT_CA<2> RT_CA<1> RT_CA<0> RT_CB<3> RT_CB<2> 
+ RT_CB<1> RT_CB<0> RT_MA<3> RT_MA<2> RT_MA<1> RT_MA<0> RT_MB<3> RT_MB<2> RT_MB<1> 
+ RT_MB<0> RT_TM_PREA_N RT_TM_PREB_N STCLKA STCLKB T_PXAA<3> T_PXAA<2> T_PXAA<1> T_PXAA<0> 
+ T_PXAB<3> T_PXAB<2> T_PXAB<1> T_PXAB<0> T_PXBA_N<7> T_PXBA_N<6> T_PXBA_N<5> T_PXBA_N<4> T_PXBA_N<3> 
+ T_PXBA_N<2> T_PXBA_N<1> T_PXBA_N<0> T_PXBB_N<7> T_PXBB_N<6> T_PXBB_N<5> T_PXBB_N<4> T_PXBB_N<3> T_PXBB_N<2> 
+ T_PXBB_N<1> T_PXBB_N<0> T_PXCA_N<7> T_PXCA_N<6> T_PXCA_N<5> T_PXCA_N<4> T_PXCA_N<3> T_PXCA_N<2> T_PXCA_N<1> 
+ T_PXCA_N<0> T_PXCB_N<7> T_PXCB_N<6> T_PXCB_N<5> T_PXCB_N<4> T_PXCB_N<3> T_PXCB_N<2> T_PXCB_N<1> T_PXCB_N<0> 
+ NET132<9> NET132<8> NET132<7> NET132<6> NET132<5> NET132<4> NET132<3> NET132<2> NET132<1> 
+ NET132<0> VDD VSS NET123 NET129  / xmc55_dps_local_ctrl8
XXDEC_BOT
+ B_PXAA<3> B_PXAA<2> B_PXAA<1> B_PXAA<0> B_PXAB<3> B_PXAB<2> B_PXAB<1> B_PXAB<0> B_PXBA_N<7> 
+ B_PXBA_N<6> B_PXBA_N<5> B_PXBA_N<4> B_PXBA_N<3> B_PXBA_N<2> B_PXBA_N<1> B_PXBA_N<0> B_PXBB_N<7> B_PXBB_N<6> 
+ B_PXBB_N<5> B_PXBB_N<4> B_PXBB_N<3> B_PXBB_N<2> B_PXBB_N<1> B_PXBB_N<0> B_PXCA_N<7> B_PXCA_N<6> B_PXCA_N<5> 
+ B_PXCA_N<4> B_PXCA_N<3> B_PXCA_N<2> B_PXCA_N<1> B_PXCA_N<0> B_PXCB_N<7> B_PXCB_N<6> B_PXCB_N<5> B_PXCB_N<4> 
+ B_PXCB_N<3> B_PXCB_N<2> B_PXCB_N<1> B_PXCB_N<0> VDD VSS B_WLA<255> B_WLA<254> B_WLA<253> 
+ B_WLA<252> B_WLA<251> B_WLA<250> B_WLA<249> B_WLA<248> B_WLA<247> B_WLA<246> B_WLA<245> B_WLA<244> 
+ B_WLA<243> B_WLA<242> B_WLA<241> B_WLA<240> B_WLA<239> B_WLA<238> B_WLA<237> B_WLA<236> B_WLA<235> 
+ B_WLA<234> B_WLA<233> B_WLA<232> B_WLA<231> B_WLA<230> B_WLA<229> B_WLA<228> B_WLA<227> B_WLA<226> 
+ B_WLA<225> B_WLA<224> B_WLA<223> B_WLA<222> B_WLA<221> B_WLA<220> B_WLA<219> B_WLA<218> B_WLA<217> 
+ B_WLA<216> B_WLA<215> B_WLA<214> B_WLA<213> B_WLA<212> B_WLA<211> B_WLA<210> B_WLA<209> B_WLA<208> 
+ B_WLA<207> B_WLA<206> B_WLA<205> B_WLA<204> B_WLA<203> B_WLA<202> B_WLA<201> B_WLA<200> B_WLA<199> 
+ B_WLA<198> B_WLA<197> B_WLA<196> B_WLA<195> B_WLA<194> B_WLA<193> B_WLA<192> B_WLA<191> B_WLA<190> 
+ B_WLA<189> B_WLA<188> B_WLA<187> B_WLA<186> B_WLA<185> B_WLA<184> B_WLA<183> B_WLA<182> B_WLA<181> 
+ B_WLA<180> B_WLA<179> B_WLA<178> B_WLA<177> B_WLA<176> B_WLA<175> B_WLA<174> B_WLA<173> B_WLA<172> 
+ B_WLA<171> B_WLA<170> B_WLA<169> B_WLA<168> B_WLA<167> B_WLA<166> B_WLA<165> B_WLA<164> B_WLA<163> 
+ B_WLA<162> B_WLA<161> B_WLA<160> B_WLA<159> B_WLA<158> B_WLA<157> B_WLA<156> B_WLA<155> B_WLA<154> 
+ B_WLA<153> B_WLA<152> B_WLA<151> B_WLA<150> B_WLA<149> B_WLA<148> B_WLA<147> B_WLA<146> B_WLA<145> 
+ B_WLA<144> B_WLA<143> B_WLA<142> B_WLA<141> B_WLA<140> B_WLA<139> B_WLA<138> B_WLA<137> B_WLA<136> 
+ B_WLA<135> B_WLA<134> B_WLA<133> B_WLA<132> B_WLA<131> B_WLA<130> B_WLA<129> B_WLA<128> B_WLA<127> 
+ B_WLA<126> B_WLA<125> B_WLA<124> B_WLA<123> B_WLA<122> B_WLA<121> B_WLA<120> B_WLA<119> B_WLA<118> 
+ B_WLA<117> B_WLA<116> B_WLA<115> B_WLA<114> B_WLA<113> B_WLA<112> B_WLA<111> B_WLA<110> B_WLA<109> 
+ B_WLA<108> B_WLA<107> B_WLA<106> B_WLA<105> B_WLA<104> B_WLA<103> B_WLA<102> B_WLA<101> B_WLA<100> 
+ B_WLA<99> B_WLA<98> B_WLA<97> B_WLA<96> B_WLA<95> B_WLA<94> B_WLA<93> B_WLA<92> B_WLA<91> 
+ B_WLA<90> B_WLA<89> B_WLA<88> B_WLA<87> B_WLA<86> B_WLA<85> B_WLA<84> B_WLA<83> B_WLA<82> 
+ B_WLA<81> B_WLA<80> B_WLA<79> B_WLA<78> B_WLA<77> B_WLA<76> B_WLA<75> B_WLA<74> B_WLA<73> 
+ B_WLA<72> B_WLA<71> B_WLA<70> B_WLA<69> B_WLA<68> B_WLA<67> B_WLA<66> B_WLA<65> B_WLA<64> 
+ B_WLA<63> B_WLA<62> B_WLA<61> B_WLA<60> B_WLA<59> B_WLA<58> B_WLA<57> B_WLA<56> B_WLA<55> 
+ B_WLA<54> B_WLA<53> B_WLA<52> B_WLA<51> B_WLA<50> B_WLA<49> B_WLA<48> B_WLA<47> B_WLA<46> 
+ B_WLA<45> B_WLA<44> B_WLA<43> B_WLA<42> B_WLA<41> B_WLA<40> B_WLA<39> B_WLA<38> B_WLA<37> 
+ B_WLA<36> B_WLA<35> B_WLA<34> B_WLA<33> B_WLA<32> B_WLA<31> B_WLA<30> B_WLA<29> B_WLA<28> 
+ B_WLA<27> B_WLA<26> B_WLA<25> B_WLA<24> B_WLA<23> B_WLA<22> B_WLA<21> B_WLA<20> B_WLA<19> 
+ B_WLA<18> B_WLA<17> B_WLA<16> B_WLA<15> B_WLA<14> B_WLA<13> B_WLA<12> B_WLA<11> B_WLA<10> 
+ B_WLA<9> B_WLA<8> B_WLA<7> B_WLA<6> B_WLA<5> B_WLA<4> B_WLA<3> B_WLA<2> B_WLA<1> 
+ B_WLA<0> B_WLB<255> B_WLB<254> B_WLB<253> B_WLB<252> B_WLB<251> B_WLB<250> B_WLB<249> B_WLB<248> 
+ B_WLB<247> B_WLB<246> B_WLB<245> B_WLB<244> B_WLB<243> B_WLB<242> B_WLB<241> B_WLB<240> B_WLB<239> 
+ B_WLB<238> B_WLB<237> B_WLB<236> B_WLB<235> B_WLB<234> B_WLB<233> B_WLB<232> B_WLB<231> B_WLB<230> 
+ B_WLB<229> B_WLB<228> B_WLB<227> B_WLB<226> B_WLB<225> B_WLB<224> B_WLB<223> B_WLB<222> B_WLB<221> 
+ B_WLB<220> B_WLB<219> B_WLB<218> B_WLB<217> B_WLB<216> B_WLB<215> B_WLB<214> B_WLB<213> B_WLB<212> 
+ B_WLB<211> B_WLB<210> B_WLB<209> B_WLB<208> B_WLB<207> B_WLB<206> B_WLB<205> B_WLB<204> B_WLB<203> 
+ B_WLB<202> B_WLB<201> B_WLB<200> B_WLB<199> B_WLB<198> B_WLB<197> B_WLB<196> B_WLB<195> B_WLB<194> 
+ B_WLB<193> B_WLB<192> B_WLB<191> B_WLB<190> B_WLB<189> B_WLB<188> B_WLB<187> B_WLB<186> B_WLB<185> 
+ B_WLB<184> B_WLB<183> B_WLB<182> B_WLB<181> B_WLB<180> B_WLB<179> B_WLB<178> B_WLB<177> B_WLB<176> 
+ B_WLB<175> B_WLB<174> B_WLB<173> B_WLB<172> B_WLB<171> B_WLB<170> B_WLB<169> B_WLB<168> B_WLB<167> 
+ B_WLB<166> B_WLB<165> B_WLB<164> B_WLB<163> B_WLB<162> B_WLB<161> B_WLB<160> B_WLB<159> B_WLB<158> 
+ B_WLB<157> B_WLB<156> B_WLB<155> B_WLB<154> B_WLB<153> B_WLB<152> B_WLB<151> B_WLB<150> B_WLB<149> 
+ B_WLB<148> B_WLB<147> B_WLB<146> B_WLB<145> B_WLB<144> B_WLB<143> B_WLB<142> B_WLB<141> B_WLB<140> 
+ B_WLB<139> B_WLB<138> B_WLB<137> B_WLB<136> B_WLB<135> B_WLB<134> B_WLB<133> B_WLB<132> B_WLB<131> 
+ B_WLB<130> B_WLB<129> B_WLB<128> B_WLB<127> B_WLB<126> B_WLB<125> B_WLB<124> B_WLB<123> B_WLB<122> 
+ B_WLB<121> B_WLB<120> B_WLB<119> B_WLB<118> B_WLB<117> B_WLB<116> B_WLB<115> B_WLB<114> B_WLB<113> 
+ B_WLB<112> B_WLB<111> B_WLB<110> B_WLB<109> B_WLB<108> B_WLB<107> B_WLB<106> B_WLB<105> B_WLB<104> 
+ B_WLB<103> B_WLB<102> B_WLB<101> B_WLB<100> B_WLB<99> B_WLB<98> B_WLB<97> B_WLB<96> B_WLB<95> 
+ B_WLB<94> B_WLB<93> B_WLB<92> B_WLB<91> B_WLB<90> B_WLB<89> B_WLB<88> B_WLB<87> B_WLB<86> 
+ B_WLB<85> B_WLB<84> B_WLB<83> B_WLB<82> B_WLB<81> B_WLB<80> B_WLB<79> B_WLB<78> B_WLB<77> 
+ B_WLB<76> B_WLB<75> B_WLB<74> B_WLB<73> B_WLB<72> B_WLB<71> B_WLB<70> B_WLB<69> B_WLB<68> 
+ B_WLB<67> B_WLB<66> B_WLB<65> B_WLB<64> B_WLB<63> B_WLB<62> B_WLB<61> B_WLB<60> B_WLB<59> 
+ B_WLB<58> B_WLB<57> B_WLB<56> B_WLB<55> B_WLB<54> B_WLB<53> B_WLB<52> B_WLB<51> B_WLB<50> 
+ B_WLB<49> B_WLB<48> B_WLB<47> B_WLB<46> B_WLB<45> B_WLB<44> B_WLB<43> B_WLB<42> B_WLB<41> 
+ B_WLB<40> B_WLB<39> B_WLB<38> B_WLB<37> B_WLB<36> B_WLB<35> B_WLB<34> B_WLB<33> B_WLB<32> 
+ B_WLB<31> B_WLB<30> B_WLB<29> B_WLB<28> B_WLB<27> B_WLB<26> B_WLB<25> B_WLB<24> B_WLB<23> 
+ B_WLB<22> B_WLB<21> B_WLB<20> B_WLB<19> B_WLB<18> B_WLB<17> B_WLB<16> B_WLB<15> B_WLB<14> 
+ B_WLB<13> B_WLB<12> B_WLB<11> B_WLB<10> B_WLB<9> B_WLB<8> B_WLB<7> B_WLB<6> B_WLB<5> 
+ B_WLB<4> B_WLB<3> B_WLB<2> B_WLB<1> B_WLB<0>  / dpram16x4096_XDECX256
XCOLLAR
+ AA<12> AA<11> AA<10> AA<9> AA<8> AA<7> AA<6> AA<5> AA<4> 
+ AA<3> AA<2> AA<1> AA<0> NET133<12> NET133<11> NET133<10> NET133<9> NET133<8> 
+ NET133<7> NET133<6> NET133<5> NET133<4> NET133<3> NET133<2> NET133<1> NET133<0> AB<12> 
+ AB<11> AB<10> AB<9> AB<8> AB<7> AB<6> AB<5> AB<4> AB<3> 
+ AB<2> AB<1> AB<0> NET131<12> NET131<11> NET131<10> NET131<9> NET131<8> NET131<7> 
+ NET131<6> NET131<5> NET131<4> NET131<3> NET131<2> NET131<1> NET131<0> CENA NET122 
+ CENB NET121 CLKA NET125 CLKB NET127 TIE_VDD TIE_VSS TM<9> 
+ TM<8> TM<7> TM<6> TM<5> TM<4> TM<3> TM<2> TM<1> TM<0> 
+ NET132<9> NET132<8> NET132<7> NET132<6> NET132<5> NET132<4> NET132<3> NET132<2> NET132<1> 
+ NET132<0> VDD VSS WENA NET123 WENB NET129  / xmc55_dps_collar_corner
.ENDS

************************************************************************
* Cell Name:    dpram16x4096
* View Name:    schematic
************************************************************************
.SUBCKT dpram16x4096
+ AA<11> AA<10> AA<9> AA<8> AA<7> AA<6> AA<5> AA<4> AA<3> 
+ AA<2> AA<1> AA<0> AB<11> AB<10> AB<9> AB<8> AB<7> AB<6> 
+ AB<5> AB<4> AB<3> AB<2> AB<1> AB<0> BWENA<15> BWENA<14> BWENA<13> 
+ BWENA<12> BWENA<11> BWENA<10> BWENA<9> BWENA<8> BWENA<7> BWENA<6> BWENA<5> BWENA<4> 
+ BWENA<3> BWENA<2> BWENA<1> BWENA<0> BWENB<15> BWENB<14> BWENB<13> BWENB<12> BWENB<11> 
+ BWENB<10> BWENB<9> BWENB<8> BWENB<7> BWENB<6> BWENB<5> BWENB<4> BWENB<3> BWENB<2> 
+ BWENB<1> BWENB<0> CENA CENB CLKA CLKB DA<15> DA<14> DA<13> 
+ DA<12> DA<11> DA<10> DA<9> DA<8> DA<7> DA<6> DA<5> DA<4> 
+ DA<3> DA<2> DA<1> DA<0> DB<15> DB<14> DB<13> DB<12> DB<11> 
+ DB<10> DB<9> DB<8> DB<7> DB<6> DB<5> DB<4> DB<3> DB<2> 
+ DB<1> DB<0> QA<15> QA<14> QA<13> QA<12> QA<11> QA<10> QA<9> 
+ QA<8> QA<7> QA<6> QA<5> QA<4> QA<3> QA<2> QA<1> QA<0> 
+ QB<15> QB<14> QB<13> QB<12> QB<11> QB<10> QB<9> QB<8> QB<7> 
+ QB<6> QB<5> QB<4> QB<3> QB<2> QB<1> QB<0> VDD VSS 
+ WENA WENB 
XDUM_EDGE<0>
+ B_WLB<255> B_WLB<254> B_WLB<253> B_WLB<252> B_WLB<251> B_WLB<250> B_WLB<249> B_WLB<248> B_WLB<247> 
+ B_WLB<246> B_WLB<245> B_WLB<244> B_WLB<243> B_WLB<242> B_WLB<241> B_WLB<240> B_WLB<239> B_WLB<238> 
+ B_WLB<237> B_WLB<236> B_WLB<235> B_WLB<234> B_WLB<233> B_WLB<232> B_WLB<231> B_WLB<230> B_WLB<229> 
+ B_WLB<228> B_WLB<227> B_WLB<226> B_WLB<225> B_WLB<224> B_WLB<223> B_WLB<222> B_WLB<221> B_WLB<220> 
+ B_WLB<219> B_WLB<218> B_WLB<217> B_WLB<216> B_WLB<215> B_WLB<214> B_WLB<213> B_WLB<212> B_WLB<211> 
+ B_WLB<210> B_WLB<209> B_WLB<208> B_WLB<207> B_WLB<206> B_WLB<205> B_WLB<204> B_WLB<203> B_WLB<202> 
+ B_WLB<201> B_WLB<200> B_WLB<199> B_WLB<198> B_WLB<197> B_WLB<196> B_WLB<195> B_WLB<194> B_WLB<193> 
+ B_WLB<192> B_WLB<191> B_WLB<190> B_WLB<189> B_WLB<188> B_WLB<187> B_WLB<186> B_WLB<185> B_WLB<184> 
+ B_WLB<183> B_WLB<182> B_WLB<181> B_WLB<180> B_WLB<179> B_WLB<178> B_WLB<177> B_WLB<176> B_WLB<175> 
+ B_WLB<174> B_WLB<173> B_WLB<172> B_WLB<171> B_WLB<170> B_WLB<169> B_WLB<168> B_WLB<167> B_WLB<166> 
+ B_WLB<165> B_WLB<164> B_WLB<163> B_WLB<162> B_WLB<161> B_WLB<160> B_WLB<159> B_WLB<158> B_WLB<157> 
+ B_WLB<156> B_WLB<155> B_WLB<154> B_WLB<153> B_WLB<152> B_WLB<151> B_WLB<150> B_WLB<149> B_WLB<148> 
+ B_WLB<147> B_WLB<146> B_WLB<145> B_WLB<144> B_WLB<143> B_WLB<142> B_WLB<141> B_WLB<140> B_WLB<139> 
+ B_WLB<138> B_WLB<137> B_WLB<136> B_WLB<135> B_WLB<134> B_WLB<133> B_WLB<132> B_WLB<131> B_WLB<130> 
+ B_WLB<129> B_WLB<128> B_WLB<127> B_WLB<126> B_WLB<125> B_WLB<124> B_WLB<123> B_WLB<122> B_WLB<121> 
+ B_WLB<120> B_WLB<119> B_WLB<118> B_WLB<117> B_WLB<116> B_WLB<115> B_WLB<114> B_WLB<113> B_WLB<112> 
+ B_WLB<111> B_WLB<110> B_WLB<109> B_WLB<108> B_WLB<107> B_WLB<106> B_WLB<105> B_WLB<104> B_WLB<103> 
+ B_WLB<102> B_WLB<101> B_WLB<100> B_WLB<99> B_WLB<98> B_WLB<97> B_WLB<96> B_WLB<95> B_WLB<94> 
+ B_WLB<93> B_WLB<92> B_WLB<91> B_WLB<90> B_WLB<89> B_WLB<88> B_WLB<87> B_WLB<86> B_WLB<85> 
+ B_WLB<84> B_WLB<83> B_WLB<82> B_WLB<81> B_WLB<80> B_WLB<79> B_WLB<78> B_WLB<77> B_WLB<76> 
+ B_WLB<75> B_WLB<74> B_WLB<73> B_WLB<72> B_WLB<71> B_WLB<70> B_WLB<69> B_WLB<68> B_WLB<67> 
+ B_WLB<66> B_WLB<65> B_WLB<64> B_WLB<63> B_WLB<62> B_WLB<61> B_WLB<60> B_WLB<59> B_WLB<58> 
+ B_WLB<57> B_WLB<56> B_WLB<55> B_WLB<54> B_WLB<53> B_WLB<52> B_WLB<51> B_WLB<50> B_WLB<49> 
+ B_WLB<48> B_WLB<47> B_WLB<46> B_WLB<45> B_WLB<44> B_WLB<43> B_WLB<42> B_WLB<41> B_WLB<40> 
+ B_WLB<39> B_WLB<38> B_WLB<37> B_WLB<36> B_WLB<35> B_WLB<34> B_WLB<33> B_WLB<32> B_WLB<31> 
+ B_WLB<30> B_WLB<29> B_WLB<28> B_WLB<27> B_WLB<26> B_WLB<25> B_WLB<24> B_WLB<23> B_WLB<22> 
+ B_WLB<21> B_WLB<20> B_WLB<19> B_WLB<18> B_WLB<17> B_WLB<16> B_WLB<15> B_WLB<14> B_WLB<13> 
+ B_WLB<12> B_WLB<11> B_WLB<10> B_WLB<9> B_WLB<8> B_WLB<7> B_WLB<6> B_WLB<5> B_WLB<4> 
+ B_WLB<3> B_WLB<2> B_WLB<1> B_WLB<0> T_WLB<255> T_WLB<254> T_WLB<253> T_WLB<252> T_WLB<251> 
+ T_WLB<250> T_WLB<249> T_WLB<248> T_WLB<247> T_WLB<246> T_WLB<245> T_WLB<244> T_WLB<243> T_WLB<242> 
+ T_WLB<241> T_WLB<240> T_WLB<239> T_WLB<238> T_WLB<237> T_WLB<236> T_WLB<235> T_WLB<234> T_WLB<233> 
+ T_WLB<232> T_WLB<231> T_WLB<230> T_WLB<229> T_WLB<228> T_WLB<227> T_WLB<226> T_WLB<225> T_WLB<224> 
+ T_WLB<223> T_WLB<222> T_WLB<221> T_WLB<220> T_WLB<219> T_WLB<218> T_WLB<217> T_WLB<216> T_WLB<215> 
+ T_WLB<214> T_WLB<213> T_WLB<212> T_WLB<211> T_WLB<210> T_WLB<209> T_WLB<208> T_WLB<207> T_WLB<206> 
+ T_WLB<205> T_WLB<204> T_WLB<203> T_WLB<202> T_WLB<201> T_WLB<200> T_WLB<199> T_WLB<198> T_WLB<197> 
+ T_WLB<196> T_WLB<195> T_WLB<194> T_WLB<193> T_WLB<192> T_WLB<191> T_WLB<190> T_WLB<189> T_WLB<188> 
+ T_WLB<187> T_WLB<186> T_WLB<185> T_WLB<184> T_WLB<183> T_WLB<182> T_WLB<181> T_WLB<180> T_WLB<179> 
+ T_WLB<178> T_WLB<177> T_WLB<176> T_WLB<175> T_WLB<174> T_WLB<173> T_WLB<172> T_WLB<171> T_WLB<170> 
+ T_WLB<169> T_WLB<168> T_WLB<167> T_WLB<166> T_WLB<165> T_WLB<164> T_WLB<163> T_WLB<162> T_WLB<161> 
+ T_WLB<160> T_WLB<159> T_WLB<158> T_WLB<157> T_WLB<156> T_WLB<155> T_WLB<154> T_WLB<153> T_WLB<152> 
+ T_WLB<151> T_WLB<150> T_WLB<149> T_WLB<148> T_WLB<147> T_WLB<146> T_WLB<145> T_WLB<144> T_WLB<143> 
+ T_WLB<142> T_WLB<141> T_WLB<140> T_WLB<139> T_WLB<138> T_WLB<137> T_WLB<136> T_WLB<135> T_WLB<134> 
+ T_WLB<133> T_WLB<132> T_WLB<131> T_WLB<130> T_WLB<129> T_WLB<128> T_WLB<127> T_WLB<126> T_WLB<125> 
+ T_WLB<124> T_WLB<123> T_WLB<122> T_WLB<121> T_WLB<120> T_WLB<119> T_WLB<118> T_WLB<117> T_WLB<116> 
+ T_WLB<115> T_WLB<114> T_WLB<113> T_WLB<112> T_WLB<111> T_WLB<110> T_WLB<109> T_WLB<108> T_WLB<107> 
+ T_WLB<106> T_WLB<105> T_WLB<104> T_WLB<103> T_WLB<102> T_WLB<101> T_WLB<100> T_WLB<99> T_WLB<98> 
+ T_WLB<97> T_WLB<96> T_WLB<95> T_WLB<94> T_WLB<93> T_WLB<92> T_WLB<91> T_WLB<90> T_WLB<89> 
+ T_WLB<88> T_WLB<87> T_WLB<86> T_WLB<85> T_WLB<84> T_WLB<83> T_WLB<82> T_WLB<81> T_WLB<80> 
+ T_WLB<79> T_WLB<78> T_WLB<77> T_WLB<76> T_WLB<75> T_WLB<74> T_WLB<73> T_WLB<72> T_WLB<71> 
+ T_WLB<70> T_WLB<69> T_WLB<68> T_WLB<67> T_WLB<66> T_WLB<65> T_WLB<64> T_WLB<63> T_WLB<62> 
+ T_WLB<61> T_WLB<60> T_WLB<59> T_WLB<58> T_WLB<57> T_WLB<56> T_WLB<55> T_WLB<54> T_WLB<53> 
+ T_WLB<52> T_WLB<51> T_WLB<50> T_WLB<49> T_WLB<48> T_WLB<47> T_WLB<46> T_WLB<45> T_WLB<44> 
+ T_WLB<43> T_WLB<42> T_WLB<41> T_WLB<40> T_WLB<39> T_WLB<38> T_WLB<37> T_WLB<36> T_WLB<35> 
+ T_WLB<34> T_WLB<33> T_WLB<32> T_WLB<31> T_WLB<30> T_WLB<29> T_WLB<28> T_WLB<27> T_WLB<26> 
+ T_WLB<25> T_WLB<24> T_WLB<23> T_WLB<22> T_WLB<21> T_WLB<20> T_WLB<19> T_WLB<18> T_WLB<17> 
+ T_WLB<16> T_WLB<15> T_WLB<14> T_WLB<13> T_WLB<12> T_WLB<11> T_WLB<10> T_WLB<9> T_WLB<8> 
+ T_WLB<7> T_WLB<6> T_WLB<5> T_WLB<4> T_WLB<3> T_WLB<2> T_WLB<1> T_WLB<0> TIE_VSS 
+ VDD VSS  / dpram16x4096_COL2X8_EDGE_ROWX256
XDUM_EDGE<1>
+ B_WLB<255> B_WLB<254> B_WLB<253> B_WLB<252> B_WLB<251> B_WLB<250> B_WLB<249> B_WLB<248> B_WLB<247> 
+ B_WLB<246> B_WLB<245> B_WLB<244> B_WLB<243> B_WLB<242> B_WLB<241> B_WLB<240> B_WLB<239> B_WLB<238> 
+ B_WLB<237> B_WLB<236> B_WLB<235> B_WLB<234> B_WLB<233> B_WLB<232> B_WLB<231> B_WLB<230> B_WLB<229> 
+ B_WLB<228> B_WLB<227> B_WLB<226> B_WLB<225> B_WLB<224> B_WLB<223> B_WLB<222> B_WLB<221> B_WLB<220> 
+ B_WLB<219> B_WLB<218> B_WLB<217> B_WLB<216> B_WLB<215> B_WLB<214> B_WLB<213> B_WLB<212> B_WLB<211> 
+ B_WLB<210> B_WLB<209> B_WLB<208> B_WLB<207> B_WLB<206> B_WLB<205> B_WLB<204> B_WLB<203> B_WLB<202> 
+ B_WLB<201> B_WLB<200> B_WLB<199> B_WLB<198> B_WLB<197> B_WLB<196> B_WLB<195> B_WLB<194> B_WLB<193> 
+ B_WLB<192> B_WLB<191> B_WLB<190> B_WLB<189> B_WLB<188> B_WLB<187> B_WLB<186> B_WLB<185> B_WLB<184> 
+ B_WLB<183> B_WLB<182> B_WLB<181> B_WLB<180> B_WLB<179> B_WLB<178> B_WLB<177> B_WLB<176> B_WLB<175> 
+ B_WLB<174> B_WLB<173> B_WLB<172> B_WLB<171> B_WLB<170> B_WLB<169> B_WLB<168> B_WLB<167> B_WLB<166> 
+ B_WLB<165> B_WLB<164> B_WLB<163> B_WLB<162> B_WLB<161> B_WLB<160> B_WLB<159> B_WLB<158> B_WLB<157> 
+ B_WLB<156> B_WLB<155> B_WLB<154> B_WLB<153> B_WLB<152> B_WLB<151> B_WLB<150> B_WLB<149> B_WLB<148> 
+ B_WLB<147> B_WLB<146> B_WLB<145> B_WLB<144> B_WLB<143> B_WLB<142> B_WLB<141> B_WLB<140> B_WLB<139> 
+ B_WLB<138> B_WLB<137> B_WLB<136> B_WLB<135> B_WLB<134> B_WLB<133> B_WLB<132> B_WLB<131> B_WLB<130> 
+ B_WLB<129> B_WLB<128> B_WLB<127> B_WLB<126> B_WLB<125> B_WLB<124> B_WLB<123> B_WLB<122> B_WLB<121> 
+ B_WLB<120> B_WLB<119> B_WLB<118> B_WLB<117> B_WLB<116> B_WLB<115> B_WLB<114> B_WLB<113> B_WLB<112> 
+ B_WLB<111> B_WLB<110> B_WLB<109> B_WLB<108> B_WLB<107> B_WLB<106> B_WLB<105> B_WLB<104> B_WLB<103> 
+ B_WLB<102> B_WLB<101> B_WLB<100> B_WLB<99> B_WLB<98> B_WLB<97> B_WLB<96> B_WLB<95> B_WLB<94> 
+ B_WLB<93> B_WLB<92> B_WLB<91> B_WLB<90> B_WLB<89> B_WLB<88> B_WLB<87> B_WLB<86> B_WLB<85> 
+ B_WLB<84> B_WLB<83> B_WLB<82> B_WLB<81> B_WLB<80> B_WLB<79> B_WLB<78> B_WLB<77> B_WLB<76> 
+ B_WLB<75> B_WLB<74> B_WLB<73> B_WLB<72> B_WLB<71> B_WLB<70> B_WLB<69> B_WLB<68> B_WLB<67> 
+ B_WLB<66> B_WLB<65> B_WLB<64> B_WLB<63> B_WLB<62> B_WLB<61> B_WLB<60> B_WLB<59> B_WLB<58> 
+ B_WLB<57> B_WLB<56> B_WLB<55> B_WLB<54> B_WLB<53> B_WLB<52> B_WLB<51> B_WLB<50> B_WLB<49> 
+ B_WLB<48> B_WLB<47> B_WLB<46> B_WLB<45> B_WLB<44> B_WLB<43> B_WLB<42> B_WLB<41> B_WLB<40> 
+ B_WLB<39> B_WLB<38> B_WLB<37> B_WLB<36> B_WLB<35> B_WLB<34> B_WLB<33> B_WLB<32> B_WLB<31> 
+ B_WLB<30> B_WLB<29> B_WLB<28> B_WLB<27> B_WLB<26> B_WLB<25> B_WLB<24> B_WLB<23> B_WLB<22> 
+ B_WLB<21> B_WLB<20> B_WLB<19> B_WLB<18> B_WLB<17> B_WLB<16> B_WLB<15> B_WLB<14> B_WLB<13> 
+ B_WLB<12> B_WLB<11> B_WLB<10> B_WLB<9> B_WLB<8> B_WLB<7> B_WLB<6> B_WLB<5> B_WLB<4> 
+ B_WLB<3> B_WLB<2> B_WLB<1> B_WLB<0> T_WLB<255> T_WLB<254> T_WLB<253> T_WLB<252> T_WLB<251> 
+ T_WLB<250> T_WLB<249> T_WLB<248> T_WLB<247> T_WLB<246> T_WLB<245> T_WLB<244> T_WLB<243> T_WLB<242> 
+ T_WLB<241> T_WLB<240> T_WLB<239> T_WLB<238> T_WLB<237> T_WLB<236> T_WLB<235> T_WLB<234> T_WLB<233> 
+ T_WLB<232> T_WLB<231> T_WLB<230> T_WLB<229> T_WLB<228> T_WLB<227> T_WLB<226> T_WLB<225> T_WLB<224> 
+ T_WLB<223> T_WLB<222> T_WLB<221> T_WLB<220> T_WLB<219> T_WLB<218> T_WLB<217> T_WLB<216> T_WLB<215> 
+ T_WLB<214> T_WLB<213> T_WLB<212> T_WLB<211> T_WLB<210> T_WLB<209> T_WLB<208> T_WLB<207> T_WLB<206> 
+ T_WLB<205> T_WLB<204> T_WLB<203> T_WLB<202> T_WLB<201> T_WLB<200> T_WLB<199> T_WLB<198> T_WLB<197> 
+ T_WLB<196> T_WLB<195> T_WLB<194> T_WLB<193> T_WLB<192> T_WLB<191> T_WLB<190> T_WLB<189> T_WLB<188> 
+ T_WLB<187> T_WLB<186> T_WLB<185> T_WLB<184> T_WLB<183> T_WLB<182> T_WLB<181> T_WLB<180> T_WLB<179> 
+ T_WLB<178> T_WLB<177> T_WLB<176> T_WLB<175> T_WLB<174> T_WLB<173> T_WLB<172> T_WLB<171> T_WLB<170> 
+ T_WLB<169> T_WLB<168> T_WLB<167> T_WLB<166> T_WLB<165> T_WLB<164> T_WLB<163> T_WLB<162> T_WLB<161> 
+ T_WLB<160> T_WLB<159> T_WLB<158> T_WLB<157> T_WLB<156> T_WLB<155> T_WLB<154> T_WLB<153> T_WLB<152> 
+ T_WLB<151> T_WLB<150> T_WLB<149> T_WLB<148> T_WLB<147> T_WLB<146> T_WLB<145> T_WLB<144> T_WLB<143> 
+ T_WLB<142> T_WLB<141> T_WLB<140> T_WLB<139> T_WLB<138> T_WLB<137> T_WLB<136> T_WLB<135> T_WLB<134> 
+ T_WLB<133> T_WLB<132> T_WLB<131> T_WLB<130> T_WLB<129> T_WLB<128> T_WLB<127> T_WLB<126> T_WLB<125> 
+ T_WLB<124> T_WLB<123> T_WLB<122> T_WLB<121> T_WLB<120> T_WLB<119> T_WLB<118> T_WLB<117> T_WLB<116> 
+ T_WLB<115> T_WLB<114> T_WLB<113> T_WLB<112> T_WLB<111> T_WLB<110> T_WLB<109> T_WLB<108> T_WLB<107> 
+ T_WLB<106> T_WLB<105> T_WLB<104> T_WLB<103> T_WLB<102> T_WLB<101> T_WLB<100> T_WLB<99> T_WLB<98> 
+ T_WLB<97> T_WLB<96> T_WLB<95> T_WLB<94> T_WLB<93> T_WLB<92> T_WLB<91> T_WLB<90> T_WLB<89> 
+ T_WLB<88> T_WLB<87> T_WLB<86> T_WLB<85> T_WLB<84> T_WLB<83> T_WLB<82> T_WLB<81> T_WLB<80> 
+ T_WLB<79> T_WLB<78> T_WLB<77> T_WLB<76> T_WLB<75> T_WLB<74> T_WLB<73> T_WLB<72> T_WLB<71> 
+ T_WLB<70> T_WLB<69> T_WLB<68> T_WLB<67> T_WLB<66> T_WLB<65> T_WLB<64> T_WLB<63> T_WLB<62> 
+ T_WLB<61> T_WLB<60> T_WLB<59> T_WLB<58> T_WLB<57> T_WLB<56> T_WLB<55> T_WLB<54> T_WLB<53> 
+ T_WLB<52> T_WLB<51> T_WLB<50> T_WLB<49> T_WLB<48> T_WLB<47> T_WLB<46> T_WLB<45> T_WLB<44> 
+ T_WLB<43> T_WLB<42> T_WLB<41> T_WLB<40> T_WLB<39> T_WLB<38> T_WLB<37> T_WLB<36> T_WLB<35> 
+ T_WLB<34> T_WLB<33> T_WLB<32> T_WLB<31> T_WLB<30> T_WLB<29> T_WLB<28> T_WLB<27> T_WLB<26> 
+ T_WLB<25> T_WLB<24> T_WLB<23> T_WLB<22> T_WLB<21> T_WLB<20> T_WLB<19> T_WLB<18> T_WLB<17> 
+ T_WLB<16> T_WLB<15> T_WLB<14> T_WLB<13> T_WLB<12> T_WLB<11> T_WLB<10> T_WLB<9> T_WLB<8> 
+ T_WLB<7> T_WLB<6> T_WLB<5> T_WLB<4> T_WLB<3> T_WLB<2> T_WLB<1> T_WLB<0> TIE_VSS 
+ VDD VSS  / dpram16x4096_COL2X8_EDGE_ROWX256
XDUM<0>
+ B_WLB<255> B_WLB<254> B_WLB<253> B_WLB<252> B_WLB<251> B_WLB<250> B_WLB<249> B_WLB<248> B_WLB<247> 
+ B_WLB<246> B_WLB<245> B_WLB<244> B_WLB<243> B_WLB<242> B_WLB<241> B_WLB<240> B_WLB<239> B_WLB<238> 
+ B_WLB<237> B_WLB<236> B_WLB<235> B_WLB<234> B_WLB<233> B_WLB<232> B_WLB<231> B_WLB<230> B_WLB<229> 
+ B_WLB<228> B_WLB<227> B_WLB<226> B_WLB<225> B_WLB<224> B_WLB<223> B_WLB<222> B_WLB<221> B_WLB<220> 
+ B_WLB<219> B_WLB<218> B_WLB<217> B_WLB<216> B_WLB<215> B_WLB<214> B_WLB<213> B_WLB<212> B_WLB<211> 
+ B_WLB<210> B_WLB<209> B_WLB<208> B_WLB<207> B_WLB<206> B_WLB<205> B_WLB<204> B_WLB<203> B_WLB<202> 
+ B_WLB<201> B_WLB<200> B_WLB<199> B_WLB<198> B_WLB<197> B_WLB<196> B_WLB<195> B_WLB<194> B_WLB<193> 
+ B_WLB<192> B_WLB<191> B_WLB<190> B_WLB<189> B_WLB<188> B_WLB<187> B_WLB<186> B_WLB<185> B_WLB<184> 
+ B_WLB<183> B_WLB<182> B_WLB<181> B_WLB<180> B_WLB<179> B_WLB<178> B_WLB<177> B_WLB<176> B_WLB<175> 
+ B_WLB<174> B_WLB<173> B_WLB<172> B_WLB<171> B_WLB<170> B_WLB<169> B_WLB<168> B_WLB<167> B_WLB<166> 
+ B_WLB<165> B_WLB<164> B_WLB<163> B_WLB<162> B_WLB<161> B_WLB<160> B_WLB<159> B_WLB<158> B_WLB<157> 
+ B_WLB<156> B_WLB<155> B_WLB<154> B_WLB<153> B_WLB<152> B_WLB<151> B_WLB<150> B_WLB<149> B_WLB<148> 
+ B_WLB<147> B_WLB<146> B_WLB<145> B_WLB<144> B_WLB<143> B_WLB<142> B_WLB<141> B_WLB<140> B_WLB<139> 
+ B_WLB<138> B_WLB<137> B_WLB<136> B_WLB<135> B_WLB<134> B_WLB<133> B_WLB<132> B_WLB<131> B_WLB<130> 
+ B_WLB<129> B_WLB<128> B_WLB<127> B_WLB<126> B_WLB<125> B_WLB<124> B_WLB<123> B_WLB<122> B_WLB<121> 
+ B_WLB<120> B_WLB<119> B_WLB<118> B_WLB<117> B_WLB<116> B_WLB<115> B_WLB<114> B_WLB<113> B_WLB<112> 
+ B_WLB<111> B_WLB<110> B_WLB<109> B_WLB<108> B_WLB<107> B_WLB<106> B_WLB<105> B_WLB<104> B_WLB<103> 
+ B_WLB<102> B_WLB<101> B_WLB<100> B_WLB<99> B_WLB<98> B_WLB<97> B_WLB<96> B_WLB<95> B_WLB<94> 
+ B_WLB<93> B_WLB<92> B_WLB<91> B_WLB<90> B_WLB<89> B_WLB<88> B_WLB<87> B_WLB<86> B_WLB<85> 
+ B_WLB<84> B_WLB<83> B_WLB<82> B_WLB<81> B_WLB<80> B_WLB<79> B_WLB<78> B_WLB<77> B_WLB<76> 
+ B_WLB<75> B_WLB<74> B_WLB<73> B_WLB<72> B_WLB<71> B_WLB<70> B_WLB<69> B_WLB<68> B_WLB<67> 
+ B_WLB<66> B_WLB<65> B_WLB<64> B_WLB<63> B_WLB<62> B_WLB<61> B_WLB<60> B_WLB<59> B_WLB<58> 
+ B_WLB<57> B_WLB<56> B_WLB<55> B_WLB<54> B_WLB<53> B_WLB<52> B_WLB<51> B_WLB<50> B_WLB<49> 
+ B_WLB<48> B_WLB<47> B_WLB<46> B_WLB<45> B_WLB<44> B_WLB<43> B_WLB<42> B_WLB<41> B_WLB<40> 
+ B_WLB<39> B_WLB<38> B_WLB<37> B_WLB<36> B_WLB<35> B_WLB<34> B_WLB<33> B_WLB<32> B_WLB<31> 
+ B_WLB<30> B_WLB<29> B_WLB<28> B_WLB<27> B_WLB<26> B_WLB<25> B_WLB<24> B_WLB<23> B_WLB<22> 
+ B_WLB<21> B_WLB<20> B_WLB<19> B_WLB<18> B_WLB<17> B_WLB<16> B_WLB<15> B_WLB<14> B_WLB<13> 
+ B_WLB<12> B_WLB<11> B_WLB<10> B_WLB<9> B_WLB<8> B_WLB<7> B_WLB<6> B_WLB<5> B_WLB<4> 
+ B_WLB<3> B_WLB<2> B_WLB<1> B_WLB<0> DBL_PD_N<3> DBL_PD_N<2> DBL_PD_N<1> DBL_PD_N<0> DWLA<1> 
+ DWLA<0> STCLKA T_WLB<255> T_WLB<254> T_WLB<253> T_WLB<252> T_WLB<251> T_WLB<250> T_WLB<249> 
+ T_WLB<248> T_WLB<247> T_WLB<246> T_WLB<245> T_WLB<244> T_WLB<243> T_WLB<242> T_WLB<241> T_WLB<240> 
+ T_WLB<239> T_WLB<238> T_WLB<237> T_WLB<236> T_WLB<235> T_WLB<234> T_WLB<233> T_WLB<232> T_WLB<231> 
+ T_WLB<230> T_WLB<229> T_WLB<228> T_WLB<227> T_WLB<226> T_WLB<225> T_WLB<224> T_WLB<223> T_WLB<222> 
+ T_WLB<221> T_WLB<220> T_WLB<219> T_WLB<218> T_WLB<217> T_WLB<216> T_WLB<215> T_WLB<214> T_WLB<213> 
+ T_WLB<212> T_WLB<211> T_WLB<210> T_WLB<209> T_WLB<208> T_WLB<207> T_WLB<206> T_WLB<205> T_WLB<204> 
+ T_WLB<203> T_WLB<202> T_WLB<201> T_WLB<200> T_WLB<199> T_WLB<198> T_WLB<197> T_WLB<196> T_WLB<195> 
+ T_WLB<194> T_WLB<193> T_WLB<192> T_WLB<191> T_WLB<190> T_WLB<189> T_WLB<188> T_WLB<187> T_WLB<186> 
+ T_WLB<185> T_WLB<184> T_WLB<183> T_WLB<182> T_WLB<181> T_WLB<180> T_WLB<179> T_WLB<178> T_WLB<177> 
+ T_WLB<176> T_WLB<175> T_WLB<174> T_WLB<173> T_WLB<172> T_WLB<171> T_WLB<170> T_WLB<169> T_WLB<168> 
+ T_WLB<167> T_WLB<166> T_WLB<165> T_WLB<164> T_WLB<163> T_WLB<162> T_WLB<161> T_WLB<160> T_WLB<159> 
+ T_WLB<158> T_WLB<157> T_WLB<156> T_WLB<155> T_WLB<154> T_WLB<153> T_WLB<152> T_WLB<151> T_WLB<150> 
+ T_WLB<149> T_WLB<148> T_WLB<147> T_WLB<146> T_WLB<145> T_WLB<144> T_WLB<143> T_WLB<142> T_WLB<141> 
+ T_WLB<140> T_WLB<139> T_WLB<138> T_WLB<137> T_WLB<136> T_WLB<135> T_WLB<134> T_WLB<133> T_WLB<132> 
+ T_WLB<131> T_WLB<130> T_WLB<129> T_WLB<128> T_WLB<127> T_WLB<126> T_WLB<125> T_WLB<124> T_WLB<123> 
+ T_WLB<122> T_WLB<121> T_WLB<120> T_WLB<119> T_WLB<118> T_WLB<117> T_WLB<116> T_WLB<115> T_WLB<114> 
+ T_WLB<113> T_WLB<112> T_WLB<111> T_WLB<110> T_WLB<109> T_WLB<108> T_WLB<107> T_WLB<106> T_WLB<105> 
+ T_WLB<104> T_WLB<103> T_WLB<102> T_WLB<101> T_WLB<100> T_WLB<99> T_WLB<98> T_WLB<97> T_WLB<96> 
+ T_WLB<95> T_WLB<94> T_WLB<93> T_WLB<92> T_WLB<91> T_WLB<90> T_WLB<89> T_WLB<88> T_WLB<87> 
+ T_WLB<86> T_WLB<85> T_WLB<84> T_WLB<83> T_WLB<82> T_WLB<81> T_WLB<80> T_WLB<79> T_WLB<78> 
+ T_WLB<77> T_WLB<76> T_WLB<75> T_WLB<74> T_WLB<73> T_WLB<72> T_WLB<71> T_WLB<70> T_WLB<69> 
+ T_WLB<68> T_WLB<67> T_WLB<66> T_WLB<65> T_WLB<64> T_WLB<63> T_WLB<62> T_WLB<61> T_WLB<60> 
+ T_WLB<59> T_WLB<58> T_WLB<57> T_WLB<56> T_WLB<55> T_WLB<54> T_WLB<53> T_WLB<52> T_WLB<51> 
+ T_WLB<50> T_WLB<49> T_WLB<48> T_WLB<47> T_WLB<46> T_WLB<45> T_WLB<44> T_WLB<43> T_WLB<42> 
+ T_WLB<41> T_WLB<40> T_WLB<39> T_WLB<38> T_WLB<37> T_WLB<36> T_WLB<35> T_WLB<34> T_WLB<33> 
+ T_WLB<32> T_WLB<31> T_WLB<30> T_WLB<29> T_WLB<28> T_WLB<27> T_WLB<26> T_WLB<25> T_WLB<24> 
+ T_WLB<23> T_WLB<22> T_WLB<21> T_WLB<20> T_WLB<19> T_WLB<18> T_WLB<17> T_WLB<16> T_WLB<15> 
+ T_WLB<14> T_WLB<13> T_WLB<12> T_WLB<11> T_WLB<10> T_WLB<9> T_WLB<8> T_WLB<7> T_WLB<6> 
+ T_WLB<5> T_WLB<4> T_WLB<3> T_WLB<2> T_WLB<1> T_WLB<0> VDD VSS  / dpram16x4096_COL2X8_DUM_ROWX256
XDUM<1>
+ B_WLB<255> B_WLB<254> B_WLB<253> B_WLB<252> B_WLB<251> B_WLB<250> B_WLB<249> B_WLB<248> B_WLB<247> 
+ B_WLB<246> B_WLB<245> B_WLB<244> B_WLB<243> B_WLB<242> B_WLB<241> B_WLB<240> B_WLB<239> B_WLB<238> 
+ B_WLB<237> B_WLB<236> B_WLB<235> B_WLB<234> B_WLB<233> B_WLB<232> B_WLB<231> B_WLB<230> B_WLB<229> 
+ B_WLB<228> B_WLB<227> B_WLB<226> B_WLB<225> B_WLB<224> B_WLB<223> B_WLB<222> B_WLB<221> B_WLB<220> 
+ B_WLB<219> B_WLB<218> B_WLB<217> B_WLB<216> B_WLB<215> B_WLB<214> B_WLB<213> B_WLB<212> B_WLB<211> 
+ B_WLB<210> B_WLB<209> B_WLB<208> B_WLB<207> B_WLB<206> B_WLB<205> B_WLB<204> B_WLB<203> B_WLB<202> 
+ B_WLB<201> B_WLB<200> B_WLB<199> B_WLB<198> B_WLB<197> B_WLB<196> B_WLB<195> B_WLB<194> B_WLB<193> 
+ B_WLB<192> B_WLB<191> B_WLB<190> B_WLB<189> B_WLB<188> B_WLB<187> B_WLB<186> B_WLB<185> B_WLB<184> 
+ B_WLB<183> B_WLB<182> B_WLB<181> B_WLB<180> B_WLB<179> B_WLB<178> B_WLB<177> B_WLB<176> B_WLB<175> 
+ B_WLB<174> B_WLB<173> B_WLB<172> B_WLB<171> B_WLB<170> B_WLB<169> B_WLB<168> B_WLB<167> B_WLB<166> 
+ B_WLB<165> B_WLB<164> B_WLB<163> B_WLB<162> B_WLB<161> B_WLB<160> B_WLB<159> B_WLB<158> B_WLB<157> 
+ B_WLB<156> B_WLB<155> B_WLB<154> B_WLB<153> B_WLB<152> B_WLB<151> B_WLB<150> B_WLB<149> B_WLB<148> 
+ B_WLB<147> B_WLB<146> B_WLB<145> B_WLB<144> B_WLB<143> B_WLB<142> B_WLB<141> B_WLB<140> B_WLB<139> 
+ B_WLB<138> B_WLB<137> B_WLB<136> B_WLB<135> B_WLB<134> B_WLB<133> B_WLB<132> B_WLB<131> B_WLB<130> 
+ B_WLB<129> B_WLB<128> B_WLB<127> B_WLB<126> B_WLB<125> B_WLB<124> B_WLB<123> B_WLB<122> B_WLB<121> 
+ B_WLB<120> B_WLB<119> B_WLB<118> B_WLB<117> B_WLB<116> B_WLB<115> B_WLB<114> B_WLB<113> B_WLB<112> 
+ B_WLB<111> B_WLB<110> B_WLB<109> B_WLB<108> B_WLB<107> B_WLB<106> B_WLB<105> B_WLB<104> B_WLB<103> 
+ B_WLB<102> B_WLB<101> B_WLB<100> B_WLB<99> B_WLB<98> B_WLB<97> B_WLB<96> B_WLB<95> B_WLB<94> 
+ B_WLB<93> B_WLB<92> B_WLB<91> B_WLB<90> B_WLB<89> B_WLB<88> B_WLB<87> B_WLB<86> B_WLB<85> 
+ B_WLB<84> B_WLB<83> B_WLB<82> B_WLB<81> B_WLB<80> B_WLB<79> B_WLB<78> B_WLB<77> B_WLB<76> 
+ B_WLB<75> B_WLB<74> B_WLB<73> B_WLB<72> B_WLB<71> B_WLB<70> B_WLB<69> B_WLB<68> B_WLB<67> 
+ B_WLB<66> B_WLB<65> B_WLB<64> B_WLB<63> B_WLB<62> B_WLB<61> B_WLB<60> B_WLB<59> B_WLB<58> 
+ B_WLB<57> B_WLB<56> B_WLB<55> B_WLB<54> B_WLB<53> B_WLB<52> B_WLB<51> B_WLB<50> B_WLB<49> 
+ B_WLB<48> B_WLB<47> B_WLB<46> B_WLB<45> B_WLB<44> B_WLB<43> B_WLB<42> B_WLB<41> B_WLB<40> 
+ B_WLB<39> B_WLB<38> B_WLB<37> B_WLB<36> B_WLB<35> B_WLB<34> B_WLB<33> B_WLB<32> B_WLB<31> 
+ B_WLB<30> B_WLB<29> B_WLB<28> B_WLB<27> B_WLB<26> B_WLB<25> B_WLB<24> B_WLB<23> B_WLB<22> 
+ B_WLB<21> B_WLB<20> B_WLB<19> B_WLB<18> B_WLB<17> B_WLB<16> B_WLB<15> B_WLB<14> B_WLB<13> 
+ B_WLB<12> B_WLB<11> B_WLB<10> B_WLB<9> B_WLB<8> B_WLB<7> B_WLB<6> B_WLB<5> B_WLB<4> 
+ B_WLB<3> B_WLB<2> B_WLB<1> B_WLB<0> DBL_PD_N<3> DBL_PD_N<2> DBL_PD_N<1> DBL_PD_N<0> DWLB<1> 
+ DWLB<0> STCLKB T_WLB<255> T_WLB<254> T_WLB<253> T_WLB<252> T_WLB<251> T_WLB<250> T_WLB<249> 
+ T_WLB<248> T_WLB<247> T_WLB<246> T_WLB<245> T_WLB<244> T_WLB<243> T_WLB<242> T_WLB<241> T_WLB<240> 
+ T_WLB<239> T_WLB<238> T_WLB<237> T_WLB<236> T_WLB<235> T_WLB<234> T_WLB<233> T_WLB<232> T_WLB<231> 
+ T_WLB<230> T_WLB<229> T_WLB<228> T_WLB<227> T_WLB<226> T_WLB<225> T_WLB<224> T_WLB<223> T_WLB<222> 
+ T_WLB<221> T_WLB<220> T_WLB<219> T_WLB<218> T_WLB<217> T_WLB<216> T_WLB<215> T_WLB<214> T_WLB<213> 
+ T_WLB<212> T_WLB<211> T_WLB<210> T_WLB<209> T_WLB<208> T_WLB<207> T_WLB<206> T_WLB<205> T_WLB<204> 
+ T_WLB<203> T_WLB<202> T_WLB<201> T_WLB<200> T_WLB<199> T_WLB<198> T_WLB<197> T_WLB<196> T_WLB<195> 
+ T_WLB<194> T_WLB<193> T_WLB<192> T_WLB<191> T_WLB<190> T_WLB<189> T_WLB<188> T_WLB<187> T_WLB<186> 
+ T_WLB<185> T_WLB<184> T_WLB<183> T_WLB<182> T_WLB<181> T_WLB<180> T_WLB<179> T_WLB<178> T_WLB<177> 
+ T_WLB<176> T_WLB<175> T_WLB<174> T_WLB<173> T_WLB<172> T_WLB<171> T_WLB<170> T_WLB<169> T_WLB<168> 
+ T_WLB<167> T_WLB<166> T_WLB<165> T_WLB<164> T_WLB<163> T_WLB<162> T_WLB<161> T_WLB<160> T_WLB<159> 
+ T_WLB<158> T_WLB<157> T_WLB<156> T_WLB<155> T_WLB<154> T_WLB<153> T_WLB<152> T_WLB<151> T_WLB<150> 
+ T_WLB<149> T_WLB<148> T_WLB<147> T_WLB<146> T_WLB<145> T_WLB<144> T_WLB<143> T_WLB<142> T_WLB<141> 
+ T_WLB<140> T_WLB<139> T_WLB<138> T_WLB<137> T_WLB<136> T_WLB<135> T_WLB<134> T_WLB<133> T_WLB<132> 
+ T_WLB<131> T_WLB<130> T_WLB<129> T_WLB<128> T_WLB<127> T_WLB<126> T_WLB<125> T_WLB<124> T_WLB<123> 
+ T_WLB<122> T_WLB<121> T_WLB<120> T_WLB<119> T_WLB<118> T_WLB<117> T_WLB<116> T_WLB<115> T_WLB<114> 
+ T_WLB<113> T_WLB<112> T_WLB<111> T_WLB<110> T_WLB<109> T_WLB<108> T_WLB<107> T_WLB<106> T_WLB<105> 
+ T_WLB<104> T_WLB<103> T_WLB<102> T_WLB<101> T_WLB<100> T_WLB<99> T_WLB<98> T_WLB<97> T_WLB<96> 
+ T_WLB<95> T_WLB<94> T_WLB<93> T_WLB<92> T_WLB<91> T_WLB<90> T_WLB<89> T_WLB<88> T_WLB<87> 
+ T_WLB<86> T_WLB<85> T_WLB<84> T_WLB<83> T_WLB<82> T_WLB<81> T_WLB<80> T_WLB<79> T_WLB<78> 
+ T_WLB<77> T_WLB<76> T_WLB<75> T_WLB<74> T_WLB<73> T_WLB<72> T_WLB<71> T_WLB<70> T_WLB<69> 
+ T_WLB<68> T_WLB<67> T_WLB<66> T_WLB<65> T_WLB<64> T_WLB<63> T_WLB<62> T_WLB<61> T_WLB<60> 
+ T_WLB<59> T_WLB<58> T_WLB<57> T_WLB<56> T_WLB<55> T_WLB<54> T_WLB<53> T_WLB<52> T_WLB<51> 
+ T_WLB<50> T_WLB<49> T_WLB<48> T_WLB<47> T_WLB<46> T_WLB<45> T_WLB<44> T_WLB<43> T_WLB<42> 
+ T_WLB<41> T_WLB<40> T_WLB<39> T_WLB<38> T_WLB<37> T_WLB<36> T_WLB<35> T_WLB<34> T_WLB<33> 
+ T_WLB<32> T_WLB<31> T_WLB<30> T_WLB<29> T_WLB<28> T_WLB<27> T_WLB<26> T_WLB<25> T_WLB<24> 
+ T_WLB<23> T_WLB<22> T_WLB<21> T_WLB<20> T_WLB<19> T_WLB<18> T_WLB<17> T_WLB<16> T_WLB<15> 
+ T_WLB<14> T_WLB<13> T_WLB<12> T_WLB<11> T_WLB<10> T_WLB<9> T_WLB<8> T_WLB<7> T_WLB<6> 
+ T_WLB<5> T_WLB<4> T_WLB<3> T_WLB<2> T_WLB<1> T_WLB<0> VDD VSS  / dpram16x4096_COL2X8_DUM_ROWX256
XCOL2<7>
+ LB_CA<3> LB_CA<2> LB_CA<1> LB_CA<0> LB_CB<3> LB_CB<2> LB_CB<1> LB_CB<0> LB_MA<3> 
+ LB_MA<2> LB_MA<1> LB_MA<0> LB_MB<3> LB_MB<2> LB_MB<1> LB_MB<0> LB_TM_PREA_N LB_TM_PREB_N 
+ B_WLA<255> B_WLA<254> B_WLA<253> B_WLA<252> B_WLA<251> B_WLA<250> B_WLA<249> B_WLA<248> B_WLA<247> 
+ B_WLA<246> B_WLA<245> B_WLA<244> B_WLA<243> B_WLA<242> B_WLA<241> B_WLA<240> B_WLA<239> B_WLA<238> 
+ B_WLA<237> B_WLA<236> B_WLA<235> B_WLA<234> B_WLA<233> B_WLA<232> B_WLA<231> B_WLA<230> B_WLA<229> 
+ B_WLA<228> B_WLA<227> B_WLA<226> B_WLA<225> B_WLA<224> B_WLA<223> B_WLA<222> B_WLA<221> B_WLA<220> 
+ B_WLA<219> B_WLA<218> B_WLA<217> B_WLA<216> B_WLA<215> B_WLA<214> B_WLA<213> B_WLA<212> B_WLA<211> 
+ B_WLA<210> B_WLA<209> B_WLA<208> B_WLA<207> B_WLA<206> B_WLA<205> B_WLA<204> B_WLA<203> B_WLA<202> 
+ B_WLA<201> B_WLA<200> B_WLA<199> B_WLA<198> B_WLA<197> B_WLA<196> B_WLA<195> B_WLA<194> B_WLA<193> 
+ B_WLA<192> B_WLA<191> B_WLA<190> B_WLA<189> B_WLA<188> B_WLA<187> B_WLA<186> B_WLA<185> B_WLA<184> 
+ B_WLA<183> B_WLA<182> B_WLA<181> B_WLA<180> B_WLA<179> B_WLA<178> B_WLA<177> B_WLA<176> B_WLA<175> 
+ B_WLA<174> B_WLA<173> B_WLA<172> B_WLA<171> B_WLA<170> B_WLA<169> B_WLA<168> B_WLA<167> B_WLA<166> 
+ B_WLA<165> B_WLA<164> B_WLA<163> B_WLA<162> B_WLA<161> B_WLA<160> B_WLA<159> B_WLA<158> B_WLA<157> 
+ B_WLA<156> B_WLA<155> B_WLA<154> B_WLA<153> B_WLA<152> B_WLA<151> B_WLA<150> B_WLA<149> B_WLA<148> 
+ B_WLA<147> B_WLA<146> B_WLA<145> B_WLA<144> B_WLA<143> B_WLA<142> B_WLA<141> B_WLA<140> B_WLA<139> 
+ B_WLA<138> B_WLA<137> B_WLA<136> B_WLA<135> B_WLA<134> B_WLA<133> B_WLA<132> B_WLA<131> B_WLA<130> 
+ B_WLA<129> B_WLA<128> B_WLA<127> B_WLA<126> B_WLA<125> B_WLA<124> B_WLA<123> B_WLA<122> B_WLA<121> 
+ B_WLA<120> B_WLA<119> B_WLA<118> B_WLA<117> B_WLA<116> B_WLA<115> B_WLA<114> B_WLA<113> B_WLA<112> 
+ B_WLA<111> B_WLA<110> B_WLA<109> B_WLA<108> B_WLA<107> B_WLA<106> B_WLA<105> B_WLA<104> B_WLA<103> 
+ B_WLA<102> B_WLA<101> B_WLA<100> B_WLA<99> B_WLA<98> B_WLA<97> B_WLA<96> B_WLA<95> B_WLA<94> 
+ B_WLA<93> B_WLA<92> B_WLA<91> B_WLA<90> B_WLA<89> B_WLA<88> B_WLA<87> B_WLA<86> B_WLA<85> 
+ B_WLA<84> B_WLA<83> B_WLA<82> B_WLA<81> B_WLA<80> B_WLA<79> B_WLA<78> B_WLA<77> B_WLA<76> 
+ B_WLA<75> B_WLA<74> B_WLA<73> B_WLA<72> B_WLA<71> B_WLA<70> B_WLA<69> B_WLA<68> B_WLA<67> 
+ B_WLA<66> B_WLA<65> B_WLA<64> B_WLA<63> B_WLA<62> B_WLA<61> B_WLA<60> B_WLA<59> B_WLA<58> 
+ B_WLA<57> B_WLA<56> B_WLA<55> B_WLA<54> B_WLA<53> B_WLA<52> B_WLA<51> B_WLA<50> B_WLA<49> 
+ B_WLA<48> B_WLA<47> B_WLA<46> B_WLA<45> B_WLA<44> B_WLA<43> B_WLA<42> B_WLA<41> B_WLA<40> 
+ B_WLA<39> B_WLA<38> B_WLA<37> B_WLA<36> B_WLA<35> B_WLA<34> B_WLA<33> B_WLA<32> B_WLA<31> 
+ B_WLA<30> B_WLA<29> B_WLA<28> B_WLA<27> B_WLA<26> B_WLA<25> B_WLA<24> B_WLA<23> B_WLA<22> 
+ B_WLA<21> B_WLA<20> B_WLA<19> B_WLA<18> B_WLA<17> B_WLA<16> B_WLA<15> B_WLA<14> B_WLA<13> 
+ B_WLA<12> B_WLA<11> B_WLA<10> B_WLA<9> B_WLA<8> B_WLA<7> B_WLA<6> B_WLA<5> B_WLA<4> 
+ B_WLA<3> B_WLA<2> B_WLA<1> B_WLA<0> B_WLB<255> B_WLB<254> B_WLB<253> B_WLB<252> B_WLB<251> 
+ B_WLB<250> B_WLB<249> B_WLB<248> B_WLB<247> B_WLB<246> B_WLB<245> B_WLB<244> B_WLB<243> B_WLB<242> 
+ B_WLB<241> B_WLB<240> B_WLB<239> B_WLB<238> B_WLB<237> B_WLB<236> B_WLB<235> B_WLB<234> B_WLB<233> 
+ B_WLB<232> B_WLB<231> B_WLB<230> B_WLB<229> B_WLB<228> B_WLB<227> B_WLB<226> B_WLB<225> B_WLB<224> 
+ B_WLB<223> B_WLB<222> B_WLB<221> B_WLB<220> B_WLB<219> B_WLB<218> B_WLB<217> B_WLB<216> B_WLB<215> 
+ B_WLB<214> B_WLB<213> B_WLB<212> B_WLB<211> B_WLB<210> B_WLB<209> B_WLB<208> B_WLB<207> B_WLB<206> 
+ B_WLB<205> B_WLB<204> B_WLB<203> B_WLB<202> B_WLB<201> B_WLB<200> B_WLB<199> B_WLB<198> B_WLB<197> 
+ B_WLB<196> B_WLB<195> B_WLB<194> B_WLB<193> B_WLB<192> B_WLB<191> B_WLB<190> B_WLB<189> B_WLB<188> 
+ B_WLB<187> B_WLB<186> B_WLB<185> B_WLB<184> B_WLB<183> B_WLB<182> B_WLB<181> B_WLB<180> B_WLB<179> 
+ B_WLB<178> B_WLB<177> B_WLB<176> B_WLB<175> B_WLB<174> B_WLB<173> B_WLB<172> B_WLB<171> B_WLB<170> 
+ B_WLB<169> B_WLB<168> B_WLB<167> B_WLB<166> B_WLB<165> B_WLB<164> B_WLB<163> B_WLB<162> B_WLB<161> 
+ B_WLB<160> B_WLB<159> B_WLB<158> B_WLB<157> B_WLB<156> B_WLB<155> B_WLB<154> B_WLB<153> B_WLB<152> 
+ B_WLB<151> B_WLB<150> B_WLB<149> B_WLB<148> B_WLB<147> B_WLB<146> B_WLB<145> B_WLB<144> B_WLB<143> 
+ B_WLB<142> B_WLB<141> B_WLB<140> B_WLB<139> B_WLB<138> B_WLB<137> B_WLB<136> B_WLB<135> B_WLB<134> 
+ B_WLB<133> B_WLB<132> B_WLB<131> B_WLB<130> B_WLB<129> B_WLB<128> B_WLB<127> B_WLB<126> B_WLB<125> 
+ B_WLB<124> B_WLB<123> B_WLB<122> B_WLB<121> B_WLB<120> B_WLB<119> B_WLB<118> B_WLB<117> B_WLB<116> 
+ B_WLB<115> B_WLB<114> B_WLB<113> B_WLB<112> B_WLB<111> B_WLB<110> B_WLB<109> B_WLB<108> B_WLB<107> 
+ B_WLB<106> B_WLB<105> B_WLB<104> B_WLB<103> B_WLB<102> B_WLB<101> B_WLB<100> B_WLB<99> B_WLB<98> 
+ B_WLB<97> B_WLB<96> B_WLB<95> B_WLB<94> B_WLB<93> B_WLB<92> B_WLB<91> B_WLB<90> B_WLB<89> 
+ B_WLB<88> B_WLB<87> B_WLB<86> B_WLB<85> B_WLB<84> B_WLB<83> B_WLB<82> B_WLB<81> B_WLB<80> 
+ B_WLB<79> B_WLB<78> B_WLB<77> B_WLB<76> B_WLB<75> B_WLB<74> B_WLB<73> B_WLB<72> B_WLB<71> 
+ B_WLB<70> B_WLB<69> B_WLB<68> B_WLB<67> B_WLB<66> B_WLB<65> B_WLB<64> B_WLB<63> B_WLB<62> 
+ B_WLB<61> B_WLB<60> B_WLB<59> B_WLB<58> B_WLB<57> B_WLB<56> B_WLB<55> B_WLB<54> B_WLB<53> 
+ B_WLB<52> B_WLB<51> B_WLB<50> B_WLB<49> B_WLB<48> B_WLB<47> B_WLB<46> B_WLB<45> B_WLB<44> 
+ B_WLB<43> B_WLB<42> B_WLB<41> B_WLB<40> B_WLB<39> B_WLB<38> B_WLB<37> B_WLB<36> B_WLB<35> 
+ B_WLB<34> B_WLB<33> B_WLB<32> B_WLB<31> B_WLB<30> B_WLB<29> B_WLB<28> B_WLB<27> B_WLB<26> 
+ B_WLB<25> B_WLB<24> B_WLB<23> B_WLB<22> B_WLB<21> B_WLB<20> B_WLB<19> B_WLB<18> B_WLB<17> 
+ B_WLB<16> B_WLB<15> B_WLB<14> B_WLB<13> B_WLB<12> B_WLB<11> B_WLB<10> B_WLB<9> B_WLB<8> 
+ B_WLB<7> B_WLB<6> B_WLB<5> B_WLB<4> B_WLB<3> B_WLB<2> B_WLB<1> B_WLB<0> BWENA<15> 
+ BWENA<14> BWENB<15> BWENB<14> L_CLK_DQA L_CLK_DQA_N L_CLK_DQB L_CLK_DQB_N DA<15> DA<14> 
+ DB<15> DB<14> DDQA<7> DDQA_N<7> DDQB<7> DDQB_N<7> L_LWEA L_LWEB QA<15> 
+ QA<14> QB<15> QB<14> L_SA_PREA_N L_SA_PREB_N L_SAEA_N L_SAEB_N LT_CA<3> LT_CA<2> 
+ LT_CA<1> LT_CA<0> LT_CB<3> LT_CB<2> LT_CB<1> LT_CB<0> LT_MA<3> LT_MA<2> LT_MA<1> 
+ LT_MA<0> LT_MB<3> LT_MB<2> LT_MB<1> LT_MB<0> LT_TM_PREA_N LT_TM_PREB_N T_WLA<255> T_WLA<254> 
+ T_WLA<253> T_WLA<252> T_WLA<251> T_WLA<250> T_WLA<249> T_WLA<248> T_WLA<247> T_WLA<246> T_WLA<245> 
+ T_WLA<244> T_WLA<243> T_WLA<242> T_WLA<241> T_WLA<240> T_WLA<239> T_WLA<238> T_WLA<237> T_WLA<236> 
+ T_WLA<235> T_WLA<234> T_WLA<233> T_WLA<232> T_WLA<231> T_WLA<230> T_WLA<229> T_WLA<228> T_WLA<227> 
+ T_WLA<226> T_WLA<225> T_WLA<224> T_WLA<223> T_WLA<222> T_WLA<221> T_WLA<220> T_WLA<219> T_WLA<218> 
+ T_WLA<217> T_WLA<216> T_WLA<215> T_WLA<214> T_WLA<213> T_WLA<212> T_WLA<211> T_WLA<210> T_WLA<209> 
+ T_WLA<208> T_WLA<207> T_WLA<206> T_WLA<205> T_WLA<204> T_WLA<203> T_WLA<202> T_WLA<201> T_WLA<200> 
+ T_WLA<199> T_WLA<198> T_WLA<197> T_WLA<196> T_WLA<195> T_WLA<194> T_WLA<193> T_WLA<192> T_WLA<191> 
+ T_WLA<190> T_WLA<189> T_WLA<188> T_WLA<187> T_WLA<186> T_WLA<185> T_WLA<184> T_WLA<183> T_WLA<182> 
+ T_WLA<181> T_WLA<180> T_WLA<179> T_WLA<178> T_WLA<177> T_WLA<176> T_WLA<175> T_WLA<174> T_WLA<173> 
+ T_WLA<172> T_WLA<171> T_WLA<170> T_WLA<169> T_WLA<168> T_WLA<167> T_WLA<166> T_WLA<165> T_WLA<164> 
+ T_WLA<163> T_WLA<162> T_WLA<161> T_WLA<160> T_WLA<159> T_WLA<158> T_WLA<157> T_WLA<156> T_WLA<155> 
+ T_WLA<154> T_WLA<153> T_WLA<152> T_WLA<151> T_WLA<150> T_WLA<149> T_WLA<148> T_WLA<147> T_WLA<146> 
+ T_WLA<145> T_WLA<144> T_WLA<143> T_WLA<142> T_WLA<141> T_WLA<140> T_WLA<139> T_WLA<138> T_WLA<137> 
+ T_WLA<136> T_WLA<135> T_WLA<134> T_WLA<133> T_WLA<132> T_WLA<131> T_WLA<130> T_WLA<129> T_WLA<128> 
+ T_WLA<127> T_WLA<126> T_WLA<125> T_WLA<124> T_WLA<123> T_WLA<122> T_WLA<121> T_WLA<120> T_WLA<119> 
+ T_WLA<118> T_WLA<117> T_WLA<116> T_WLA<115> T_WLA<114> T_WLA<113> T_WLA<112> T_WLA<111> T_WLA<110> 
+ T_WLA<109> T_WLA<108> T_WLA<107> T_WLA<106> T_WLA<105> T_WLA<104> T_WLA<103> T_WLA<102> T_WLA<101> 
+ T_WLA<100> T_WLA<99> T_WLA<98> T_WLA<97> T_WLA<96> T_WLA<95> T_WLA<94> T_WLA<93> T_WLA<92> 
+ T_WLA<91> T_WLA<90> T_WLA<89> T_WLA<88> T_WLA<87> T_WLA<86> T_WLA<85> T_WLA<84> T_WLA<83> 
+ T_WLA<82> T_WLA<81> T_WLA<80> T_WLA<79> T_WLA<78> T_WLA<77> T_WLA<76> T_WLA<75> T_WLA<74> 
+ T_WLA<73> T_WLA<72> T_WLA<71> T_WLA<70> T_WLA<69> T_WLA<68> T_WLA<67> T_WLA<66> T_WLA<65> 
+ T_WLA<64> T_WLA<63> T_WLA<62> T_WLA<61> T_WLA<60> T_WLA<59> T_WLA<58> T_WLA<57> T_WLA<56> 
+ T_WLA<55> T_WLA<54> T_WLA<53> T_WLA<52> T_WLA<51> T_WLA<50> T_WLA<49> T_WLA<48> T_WLA<47> 
+ T_WLA<46> T_WLA<45> T_WLA<44> T_WLA<43> T_WLA<42> T_WLA<41> T_WLA<40> T_WLA<39> T_WLA<38> 
+ T_WLA<37> T_WLA<36> T_WLA<35> T_WLA<34> T_WLA<33> T_WLA<32> T_WLA<31> T_WLA<30> T_WLA<29> 
+ T_WLA<28> T_WLA<27> T_WLA<26> T_WLA<25> T_WLA<24> T_WLA<23> T_WLA<22> T_WLA<21> T_WLA<20> 
+ T_WLA<19> T_WLA<18> T_WLA<17> T_WLA<16> T_WLA<15> T_WLA<14> T_WLA<13> T_WLA<12> T_WLA<11> 
+ T_WLA<10> T_WLA<9> T_WLA<8> T_WLA<7> T_WLA<6> T_WLA<5> T_WLA<4> T_WLA<3> T_WLA<2> 
+ T_WLA<1> T_WLA<0> T_WLB<255> T_WLB<254> T_WLB<253> T_WLB<252> T_WLB<251> T_WLB<250> T_WLB<249> 
+ T_WLB<248> T_WLB<247> T_WLB<246> T_WLB<245> T_WLB<244> T_WLB<243> T_WLB<242> T_WLB<241> T_WLB<240> 
+ T_WLB<239> T_WLB<238> T_WLB<237> T_WLB<236> T_WLB<235> T_WLB<234> T_WLB<233> T_WLB<232> T_WLB<231> 
+ T_WLB<230> T_WLB<229> T_WLB<228> T_WLB<227> T_WLB<226> T_WLB<225> T_WLB<224> T_WLB<223> T_WLB<222> 
+ T_WLB<221> T_WLB<220> T_WLB<219> T_WLB<218> T_WLB<217> T_WLB<216> T_WLB<215> T_WLB<214> T_WLB<213> 
+ T_WLB<212> T_WLB<211> T_WLB<210> T_WLB<209> T_WLB<208> T_WLB<207> T_WLB<206> T_WLB<205> T_WLB<204> 
+ T_WLB<203> T_WLB<202> T_WLB<201> T_WLB<200> T_WLB<199> T_WLB<198> T_WLB<197> T_WLB<196> T_WLB<195> 
+ T_WLB<194> T_WLB<193> T_WLB<192> T_WLB<191> T_WLB<190> T_WLB<189> T_WLB<188> T_WLB<187> T_WLB<186> 
+ T_WLB<185> T_WLB<184> T_WLB<183> T_WLB<182> T_WLB<181> T_WLB<180> T_WLB<179> T_WLB<178> T_WLB<177> 
+ T_WLB<176> T_WLB<175> T_WLB<174> T_WLB<173> T_WLB<172> T_WLB<171> T_WLB<170> T_WLB<169> T_WLB<168> 
+ T_WLB<167> T_WLB<166> T_WLB<165> T_WLB<164> T_WLB<163> T_WLB<162> T_WLB<161> T_WLB<160> T_WLB<159> 
+ T_WLB<158> T_WLB<157> T_WLB<156> T_WLB<155> T_WLB<154> T_WLB<153> T_WLB<152> T_WLB<151> T_WLB<150> 
+ T_WLB<149> T_WLB<148> T_WLB<147> T_WLB<146> T_WLB<145> T_WLB<144> T_WLB<143> T_WLB<142> T_WLB<141> 
+ T_WLB<140> T_WLB<139> T_WLB<138> T_WLB<137> T_WLB<136> T_WLB<135> T_WLB<134> T_WLB<133> T_WLB<132> 
+ T_WLB<131> T_WLB<130> T_WLB<129> T_WLB<128> T_WLB<127> T_WLB<126> T_WLB<125> T_WLB<124> T_WLB<123> 
+ T_WLB<122> T_WLB<121> T_WLB<120> T_WLB<119> T_WLB<118> T_WLB<117> T_WLB<116> T_WLB<115> T_WLB<114> 
+ T_WLB<113> T_WLB<112> T_WLB<111> T_WLB<110> T_WLB<109> T_WLB<108> T_WLB<107> T_WLB<106> T_WLB<105> 
+ T_WLB<104> T_WLB<103> T_WLB<102> T_WLB<101> T_WLB<100> T_WLB<99> T_WLB<98> T_WLB<97> T_WLB<96> 
+ T_WLB<95> T_WLB<94> T_WLB<93> T_WLB<92> T_WLB<91> T_WLB<90> T_WLB<89> T_WLB<88> T_WLB<87> 
+ T_WLB<86> T_WLB<85> T_WLB<84> T_WLB<83> T_WLB<82> T_WLB<81> T_WLB<80> T_WLB<79> T_WLB<78> 
+ T_WLB<77> T_WLB<76> T_WLB<75> T_WLB<74> T_WLB<73> T_WLB<72> T_WLB<71> T_WLB<70> T_WLB<69> 
+ T_WLB<68> T_WLB<67> T_WLB<66> T_WLB<65> T_WLB<64> T_WLB<63> T_WLB<62> T_WLB<61> T_WLB<60> 
+ T_WLB<59> T_WLB<58> T_WLB<57> T_WLB<56> T_WLB<55> T_WLB<54> T_WLB<53> T_WLB<52> T_WLB<51> 
+ T_WLB<50> T_WLB<49> T_WLB<48> T_WLB<47> T_WLB<46> T_WLB<45> T_WLB<44> T_WLB<43> T_WLB<42> 
+ T_WLB<41> T_WLB<40> T_WLB<39> T_WLB<38> T_WLB<37> T_WLB<36> T_WLB<35> T_WLB<34> T_WLB<33> 
+ T_WLB<32> T_WLB<31> T_WLB<30> T_WLB<29> T_WLB<28> T_WLB<27> T_WLB<26> T_WLB<25> T_WLB<24> 
+ T_WLB<23> T_WLB<22> T_WLB<21> T_WLB<20> T_WLB<19> T_WLB<18> T_WLB<17> T_WLB<16> T_WLB<15> 
+ T_WLB<14> T_WLB<13> T_WLB<12> T_WLB<11> T_WLB<10> T_WLB<9> T_WLB<8> T_WLB<7> T_WLB<6> 
+ T_WLB<5> T_WLB<4> T_WLB<3> T_WLB<2> T_WLB<1> T_WLB<0> VDD VSS  / dpram16x4096_SingleCOL2X8_ROWX256
XCOL2<6>
+ LB_CA<3> LB_CA<2> LB_CA<1> LB_CA<0> LB_CB<3> LB_CB<2> LB_CB<1> LB_CB<0> LB_MA<3> 
+ LB_MA<2> LB_MA<1> LB_MA<0> LB_MB<3> LB_MB<2> LB_MB<1> LB_MB<0> LB_TM_PREA_N LB_TM_PREB_N 
+ B_WLA<255> B_WLA<254> B_WLA<253> B_WLA<252> B_WLA<251> B_WLA<250> B_WLA<249> B_WLA<248> B_WLA<247> 
+ B_WLA<246> B_WLA<245> B_WLA<244> B_WLA<243> B_WLA<242> B_WLA<241> B_WLA<240> B_WLA<239> B_WLA<238> 
+ B_WLA<237> B_WLA<236> B_WLA<235> B_WLA<234> B_WLA<233> B_WLA<232> B_WLA<231> B_WLA<230> B_WLA<229> 
+ B_WLA<228> B_WLA<227> B_WLA<226> B_WLA<225> B_WLA<224> B_WLA<223> B_WLA<222> B_WLA<221> B_WLA<220> 
+ B_WLA<219> B_WLA<218> B_WLA<217> B_WLA<216> B_WLA<215> B_WLA<214> B_WLA<213> B_WLA<212> B_WLA<211> 
+ B_WLA<210> B_WLA<209> B_WLA<208> B_WLA<207> B_WLA<206> B_WLA<205> B_WLA<204> B_WLA<203> B_WLA<202> 
+ B_WLA<201> B_WLA<200> B_WLA<199> B_WLA<198> B_WLA<197> B_WLA<196> B_WLA<195> B_WLA<194> B_WLA<193> 
+ B_WLA<192> B_WLA<191> B_WLA<190> B_WLA<189> B_WLA<188> B_WLA<187> B_WLA<186> B_WLA<185> B_WLA<184> 
+ B_WLA<183> B_WLA<182> B_WLA<181> B_WLA<180> B_WLA<179> B_WLA<178> B_WLA<177> B_WLA<176> B_WLA<175> 
+ B_WLA<174> B_WLA<173> B_WLA<172> B_WLA<171> B_WLA<170> B_WLA<169> B_WLA<168> B_WLA<167> B_WLA<166> 
+ B_WLA<165> B_WLA<164> B_WLA<163> B_WLA<162> B_WLA<161> B_WLA<160> B_WLA<159> B_WLA<158> B_WLA<157> 
+ B_WLA<156> B_WLA<155> B_WLA<154> B_WLA<153> B_WLA<152> B_WLA<151> B_WLA<150> B_WLA<149> B_WLA<148> 
+ B_WLA<147> B_WLA<146> B_WLA<145> B_WLA<144> B_WLA<143> B_WLA<142> B_WLA<141> B_WLA<140> B_WLA<139> 
+ B_WLA<138> B_WLA<137> B_WLA<136> B_WLA<135> B_WLA<134> B_WLA<133> B_WLA<132> B_WLA<131> B_WLA<130> 
+ B_WLA<129> B_WLA<128> B_WLA<127> B_WLA<126> B_WLA<125> B_WLA<124> B_WLA<123> B_WLA<122> B_WLA<121> 
+ B_WLA<120> B_WLA<119> B_WLA<118> B_WLA<117> B_WLA<116> B_WLA<115> B_WLA<114> B_WLA<113> B_WLA<112> 
+ B_WLA<111> B_WLA<110> B_WLA<109> B_WLA<108> B_WLA<107> B_WLA<106> B_WLA<105> B_WLA<104> B_WLA<103> 
+ B_WLA<102> B_WLA<101> B_WLA<100> B_WLA<99> B_WLA<98> B_WLA<97> B_WLA<96> B_WLA<95> B_WLA<94> 
+ B_WLA<93> B_WLA<92> B_WLA<91> B_WLA<90> B_WLA<89> B_WLA<88> B_WLA<87> B_WLA<86> B_WLA<85> 
+ B_WLA<84> B_WLA<83> B_WLA<82> B_WLA<81> B_WLA<80> B_WLA<79> B_WLA<78> B_WLA<77> B_WLA<76> 
+ B_WLA<75> B_WLA<74> B_WLA<73> B_WLA<72> B_WLA<71> B_WLA<70> B_WLA<69> B_WLA<68> B_WLA<67> 
+ B_WLA<66> B_WLA<65> B_WLA<64> B_WLA<63> B_WLA<62> B_WLA<61> B_WLA<60> B_WLA<59> B_WLA<58> 
+ B_WLA<57> B_WLA<56> B_WLA<55> B_WLA<54> B_WLA<53> B_WLA<52> B_WLA<51> B_WLA<50> B_WLA<49> 
+ B_WLA<48> B_WLA<47> B_WLA<46> B_WLA<45> B_WLA<44> B_WLA<43> B_WLA<42> B_WLA<41> B_WLA<40> 
+ B_WLA<39> B_WLA<38> B_WLA<37> B_WLA<36> B_WLA<35> B_WLA<34> B_WLA<33> B_WLA<32> B_WLA<31> 
+ B_WLA<30> B_WLA<29> B_WLA<28> B_WLA<27> B_WLA<26> B_WLA<25> B_WLA<24> B_WLA<23> B_WLA<22> 
+ B_WLA<21> B_WLA<20> B_WLA<19> B_WLA<18> B_WLA<17> B_WLA<16> B_WLA<15> B_WLA<14> B_WLA<13> 
+ B_WLA<12> B_WLA<11> B_WLA<10> B_WLA<9> B_WLA<8> B_WLA<7> B_WLA<6> B_WLA<5> B_WLA<4> 
+ B_WLA<3> B_WLA<2> B_WLA<1> B_WLA<0> B_WLB<255> B_WLB<254> B_WLB<253> B_WLB<252> B_WLB<251> 
+ B_WLB<250> B_WLB<249> B_WLB<248> B_WLB<247> B_WLB<246> B_WLB<245> B_WLB<244> B_WLB<243> B_WLB<242> 
+ B_WLB<241> B_WLB<240> B_WLB<239> B_WLB<238> B_WLB<237> B_WLB<236> B_WLB<235> B_WLB<234> B_WLB<233> 
+ B_WLB<232> B_WLB<231> B_WLB<230> B_WLB<229> B_WLB<228> B_WLB<227> B_WLB<226> B_WLB<225> B_WLB<224> 
+ B_WLB<223> B_WLB<222> B_WLB<221> B_WLB<220> B_WLB<219> B_WLB<218> B_WLB<217> B_WLB<216> B_WLB<215> 
+ B_WLB<214> B_WLB<213> B_WLB<212> B_WLB<211> B_WLB<210> B_WLB<209> B_WLB<208> B_WLB<207> B_WLB<206> 
+ B_WLB<205> B_WLB<204> B_WLB<203> B_WLB<202> B_WLB<201> B_WLB<200> B_WLB<199> B_WLB<198> B_WLB<197> 
+ B_WLB<196> B_WLB<195> B_WLB<194> B_WLB<193> B_WLB<192> B_WLB<191> B_WLB<190> B_WLB<189> B_WLB<188> 
+ B_WLB<187> B_WLB<186> B_WLB<185> B_WLB<184> B_WLB<183> B_WLB<182> B_WLB<181> B_WLB<180> B_WLB<179> 
+ B_WLB<178> B_WLB<177> B_WLB<176> B_WLB<175> B_WLB<174> B_WLB<173> B_WLB<172> B_WLB<171> B_WLB<170> 
+ B_WLB<169> B_WLB<168> B_WLB<167> B_WLB<166> B_WLB<165> B_WLB<164> B_WLB<163> B_WLB<162> B_WLB<161> 
+ B_WLB<160> B_WLB<159> B_WLB<158> B_WLB<157> B_WLB<156> B_WLB<155> B_WLB<154> B_WLB<153> B_WLB<152> 
+ B_WLB<151> B_WLB<150> B_WLB<149> B_WLB<148> B_WLB<147> B_WLB<146> B_WLB<145> B_WLB<144> B_WLB<143> 
+ B_WLB<142> B_WLB<141> B_WLB<140> B_WLB<139> B_WLB<138> B_WLB<137> B_WLB<136> B_WLB<135> B_WLB<134> 
+ B_WLB<133> B_WLB<132> B_WLB<131> B_WLB<130> B_WLB<129> B_WLB<128> B_WLB<127> B_WLB<126> B_WLB<125> 
+ B_WLB<124> B_WLB<123> B_WLB<122> B_WLB<121> B_WLB<120> B_WLB<119> B_WLB<118> B_WLB<117> B_WLB<116> 
+ B_WLB<115> B_WLB<114> B_WLB<113> B_WLB<112> B_WLB<111> B_WLB<110> B_WLB<109> B_WLB<108> B_WLB<107> 
+ B_WLB<106> B_WLB<105> B_WLB<104> B_WLB<103> B_WLB<102> B_WLB<101> B_WLB<100> B_WLB<99> B_WLB<98> 
+ B_WLB<97> B_WLB<96> B_WLB<95> B_WLB<94> B_WLB<93> B_WLB<92> B_WLB<91> B_WLB<90> B_WLB<89> 
+ B_WLB<88> B_WLB<87> B_WLB<86> B_WLB<85> B_WLB<84> B_WLB<83> B_WLB<82> B_WLB<81> B_WLB<80> 
+ B_WLB<79> B_WLB<78> B_WLB<77> B_WLB<76> B_WLB<75> B_WLB<74> B_WLB<73> B_WLB<72> B_WLB<71> 
+ B_WLB<70> B_WLB<69> B_WLB<68> B_WLB<67> B_WLB<66> B_WLB<65> B_WLB<64> B_WLB<63> B_WLB<62> 
+ B_WLB<61> B_WLB<60> B_WLB<59> B_WLB<58> B_WLB<57> B_WLB<56> B_WLB<55> B_WLB<54> B_WLB<53> 
+ B_WLB<52> B_WLB<51> B_WLB<50> B_WLB<49> B_WLB<48> B_WLB<47> B_WLB<46> B_WLB<45> B_WLB<44> 
+ B_WLB<43> B_WLB<42> B_WLB<41> B_WLB<40> B_WLB<39> B_WLB<38> B_WLB<37> B_WLB<36> B_WLB<35> 
+ B_WLB<34> B_WLB<33> B_WLB<32> B_WLB<31> B_WLB<30> B_WLB<29> B_WLB<28> B_WLB<27> B_WLB<26> 
+ B_WLB<25> B_WLB<24> B_WLB<23> B_WLB<22> B_WLB<21> B_WLB<20> B_WLB<19> B_WLB<18> B_WLB<17> 
+ B_WLB<16> B_WLB<15> B_WLB<14> B_WLB<13> B_WLB<12> B_WLB<11> B_WLB<10> B_WLB<9> B_WLB<8> 
+ B_WLB<7> B_WLB<6> B_WLB<5> B_WLB<4> B_WLB<3> B_WLB<2> B_WLB<1> B_WLB<0> BWENA<13> 
+ BWENA<12> BWENB<13> BWENB<12> L_CLK_DQA L_CLK_DQA_N L_CLK_DQB L_CLK_DQB_N DA<13> DA<12> 
+ DB<13> DB<12> DDQA<6> DDQA_N<6> DDQB<6> DDQB_N<6> L_LWEA L_LWEB QA<13> 
+ QA<12> QB<13> QB<12> L_SA_PREA_N L_SA_PREB_N L_SAEA_N L_SAEB_N LT_CA<3> LT_CA<2> 
+ LT_CA<1> LT_CA<0> LT_CB<3> LT_CB<2> LT_CB<1> LT_CB<0> LT_MA<3> LT_MA<2> LT_MA<1> 
+ LT_MA<0> LT_MB<3> LT_MB<2> LT_MB<1> LT_MB<0> LT_TM_PREA_N LT_TM_PREB_N T_WLA<255> T_WLA<254> 
+ T_WLA<253> T_WLA<252> T_WLA<251> T_WLA<250> T_WLA<249> T_WLA<248> T_WLA<247> T_WLA<246> T_WLA<245> 
+ T_WLA<244> T_WLA<243> T_WLA<242> T_WLA<241> T_WLA<240> T_WLA<239> T_WLA<238> T_WLA<237> T_WLA<236> 
+ T_WLA<235> T_WLA<234> T_WLA<233> T_WLA<232> T_WLA<231> T_WLA<230> T_WLA<229> T_WLA<228> T_WLA<227> 
+ T_WLA<226> T_WLA<225> T_WLA<224> T_WLA<223> T_WLA<222> T_WLA<221> T_WLA<220> T_WLA<219> T_WLA<218> 
+ T_WLA<217> T_WLA<216> T_WLA<215> T_WLA<214> T_WLA<213> T_WLA<212> T_WLA<211> T_WLA<210> T_WLA<209> 
+ T_WLA<208> T_WLA<207> T_WLA<206> T_WLA<205> T_WLA<204> T_WLA<203> T_WLA<202> T_WLA<201> T_WLA<200> 
+ T_WLA<199> T_WLA<198> T_WLA<197> T_WLA<196> T_WLA<195> T_WLA<194> T_WLA<193> T_WLA<192> T_WLA<191> 
+ T_WLA<190> T_WLA<189> T_WLA<188> T_WLA<187> T_WLA<186> T_WLA<185> T_WLA<184> T_WLA<183> T_WLA<182> 
+ T_WLA<181> T_WLA<180> T_WLA<179> T_WLA<178> T_WLA<177> T_WLA<176> T_WLA<175> T_WLA<174> T_WLA<173> 
+ T_WLA<172> T_WLA<171> T_WLA<170> T_WLA<169> T_WLA<168> T_WLA<167> T_WLA<166> T_WLA<165> T_WLA<164> 
+ T_WLA<163> T_WLA<162> T_WLA<161> T_WLA<160> T_WLA<159> T_WLA<158> T_WLA<157> T_WLA<156> T_WLA<155> 
+ T_WLA<154> T_WLA<153> T_WLA<152> T_WLA<151> T_WLA<150> T_WLA<149> T_WLA<148> T_WLA<147> T_WLA<146> 
+ T_WLA<145> T_WLA<144> T_WLA<143> T_WLA<142> T_WLA<141> T_WLA<140> T_WLA<139> T_WLA<138> T_WLA<137> 
+ T_WLA<136> T_WLA<135> T_WLA<134> T_WLA<133> T_WLA<132> T_WLA<131> T_WLA<130> T_WLA<129> T_WLA<128> 
+ T_WLA<127> T_WLA<126> T_WLA<125> T_WLA<124> T_WLA<123> T_WLA<122> T_WLA<121> T_WLA<120> T_WLA<119> 
+ T_WLA<118> T_WLA<117> T_WLA<116> T_WLA<115> T_WLA<114> T_WLA<113> T_WLA<112> T_WLA<111> T_WLA<110> 
+ T_WLA<109> T_WLA<108> T_WLA<107> T_WLA<106> T_WLA<105> T_WLA<104> T_WLA<103> T_WLA<102> T_WLA<101> 
+ T_WLA<100> T_WLA<99> T_WLA<98> T_WLA<97> T_WLA<96> T_WLA<95> T_WLA<94> T_WLA<93> T_WLA<92> 
+ T_WLA<91> T_WLA<90> T_WLA<89> T_WLA<88> T_WLA<87> T_WLA<86> T_WLA<85> T_WLA<84> T_WLA<83> 
+ T_WLA<82> T_WLA<81> T_WLA<80> T_WLA<79> T_WLA<78> T_WLA<77> T_WLA<76> T_WLA<75> T_WLA<74> 
+ T_WLA<73> T_WLA<72> T_WLA<71> T_WLA<70> T_WLA<69> T_WLA<68> T_WLA<67> T_WLA<66> T_WLA<65> 
+ T_WLA<64> T_WLA<63> T_WLA<62> T_WLA<61> T_WLA<60> T_WLA<59> T_WLA<58> T_WLA<57> T_WLA<56> 
+ T_WLA<55> T_WLA<54> T_WLA<53> T_WLA<52> T_WLA<51> T_WLA<50> T_WLA<49> T_WLA<48> T_WLA<47> 
+ T_WLA<46> T_WLA<45> T_WLA<44> T_WLA<43> T_WLA<42> T_WLA<41> T_WLA<40> T_WLA<39> T_WLA<38> 
+ T_WLA<37> T_WLA<36> T_WLA<35> T_WLA<34> T_WLA<33> T_WLA<32> T_WLA<31> T_WLA<30> T_WLA<29> 
+ T_WLA<28> T_WLA<27> T_WLA<26> T_WLA<25> T_WLA<24> T_WLA<23> T_WLA<22> T_WLA<21> T_WLA<20> 
+ T_WLA<19> T_WLA<18> T_WLA<17> T_WLA<16> T_WLA<15> T_WLA<14> T_WLA<13> T_WLA<12> T_WLA<11> 
+ T_WLA<10> T_WLA<9> T_WLA<8> T_WLA<7> T_WLA<6> T_WLA<5> T_WLA<4> T_WLA<3> T_WLA<2> 
+ T_WLA<1> T_WLA<0> T_WLB<255> T_WLB<254> T_WLB<253> T_WLB<252> T_WLB<251> T_WLB<250> T_WLB<249> 
+ T_WLB<248> T_WLB<247> T_WLB<246> T_WLB<245> T_WLB<244> T_WLB<243> T_WLB<242> T_WLB<241> T_WLB<240> 
+ T_WLB<239> T_WLB<238> T_WLB<237> T_WLB<236> T_WLB<235> T_WLB<234> T_WLB<233> T_WLB<232> T_WLB<231> 
+ T_WLB<230> T_WLB<229> T_WLB<228> T_WLB<227> T_WLB<226> T_WLB<225> T_WLB<224> T_WLB<223> T_WLB<222> 
+ T_WLB<221> T_WLB<220> T_WLB<219> T_WLB<218> T_WLB<217> T_WLB<216> T_WLB<215> T_WLB<214> T_WLB<213> 
+ T_WLB<212> T_WLB<211> T_WLB<210> T_WLB<209> T_WLB<208> T_WLB<207> T_WLB<206> T_WLB<205> T_WLB<204> 
+ T_WLB<203> T_WLB<202> T_WLB<201> T_WLB<200> T_WLB<199> T_WLB<198> T_WLB<197> T_WLB<196> T_WLB<195> 
+ T_WLB<194> T_WLB<193> T_WLB<192> T_WLB<191> T_WLB<190> T_WLB<189> T_WLB<188> T_WLB<187> T_WLB<186> 
+ T_WLB<185> T_WLB<184> T_WLB<183> T_WLB<182> T_WLB<181> T_WLB<180> T_WLB<179> T_WLB<178> T_WLB<177> 
+ T_WLB<176> T_WLB<175> T_WLB<174> T_WLB<173> T_WLB<172> T_WLB<171> T_WLB<170> T_WLB<169> T_WLB<168> 
+ T_WLB<167> T_WLB<166> T_WLB<165> T_WLB<164> T_WLB<163> T_WLB<162> T_WLB<161> T_WLB<160> T_WLB<159> 
+ T_WLB<158> T_WLB<157> T_WLB<156> T_WLB<155> T_WLB<154> T_WLB<153> T_WLB<152> T_WLB<151> T_WLB<150> 
+ T_WLB<149> T_WLB<148> T_WLB<147> T_WLB<146> T_WLB<145> T_WLB<144> T_WLB<143> T_WLB<142> T_WLB<141> 
+ T_WLB<140> T_WLB<139> T_WLB<138> T_WLB<137> T_WLB<136> T_WLB<135> T_WLB<134> T_WLB<133> T_WLB<132> 
+ T_WLB<131> T_WLB<130> T_WLB<129> T_WLB<128> T_WLB<127> T_WLB<126> T_WLB<125> T_WLB<124> T_WLB<123> 
+ T_WLB<122> T_WLB<121> T_WLB<120> T_WLB<119> T_WLB<118> T_WLB<117> T_WLB<116> T_WLB<115> T_WLB<114> 
+ T_WLB<113> T_WLB<112> T_WLB<111> T_WLB<110> T_WLB<109> T_WLB<108> T_WLB<107> T_WLB<106> T_WLB<105> 
+ T_WLB<104> T_WLB<103> T_WLB<102> T_WLB<101> T_WLB<100> T_WLB<99> T_WLB<98> T_WLB<97> T_WLB<96> 
+ T_WLB<95> T_WLB<94> T_WLB<93> T_WLB<92> T_WLB<91> T_WLB<90> T_WLB<89> T_WLB<88> T_WLB<87> 
+ T_WLB<86> T_WLB<85> T_WLB<84> T_WLB<83> T_WLB<82> T_WLB<81> T_WLB<80> T_WLB<79> T_WLB<78> 
+ T_WLB<77> T_WLB<76> T_WLB<75> T_WLB<74> T_WLB<73> T_WLB<72> T_WLB<71> T_WLB<70> T_WLB<69> 
+ T_WLB<68> T_WLB<67> T_WLB<66> T_WLB<65> T_WLB<64> T_WLB<63> T_WLB<62> T_WLB<61> T_WLB<60> 
+ T_WLB<59> T_WLB<58> T_WLB<57> T_WLB<56> T_WLB<55> T_WLB<54> T_WLB<53> T_WLB<52> T_WLB<51> 
+ T_WLB<50> T_WLB<49> T_WLB<48> T_WLB<47> T_WLB<46> T_WLB<45> T_WLB<44> T_WLB<43> T_WLB<42> 
+ T_WLB<41> T_WLB<40> T_WLB<39> T_WLB<38> T_WLB<37> T_WLB<36> T_WLB<35> T_WLB<34> T_WLB<33> 
+ T_WLB<32> T_WLB<31> T_WLB<30> T_WLB<29> T_WLB<28> T_WLB<27> T_WLB<26> T_WLB<25> T_WLB<24> 
+ T_WLB<23> T_WLB<22> T_WLB<21> T_WLB<20> T_WLB<19> T_WLB<18> T_WLB<17> T_WLB<16> T_WLB<15> 
+ T_WLB<14> T_WLB<13> T_WLB<12> T_WLB<11> T_WLB<10> T_WLB<9> T_WLB<8> T_WLB<7> T_WLB<6> 
+ T_WLB<5> T_WLB<4> T_WLB<3> T_WLB<2> T_WLB<1> T_WLB<0> VDD VSS  / dpram16x4096_SingleCOL2X8_ROWX256
XCOL2<5>
+ LB_CA<3> LB_CA<2> LB_CA<1> LB_CA<0> LB_CB<3> LB_CB<2> LB_CB<1> LB_CB<0> LB_MA<3> 
+ LB_MA<2> LB_MA<1> LB_MA<0> LB_MB<3> LB_MB<2> LB_MB<1> LB_MB<0> LB_TM_PREA_N LB_TM_PREB_N 
+ B_WLA<255> B_WLA<254> B_WLA<253> B_WLA<252> B_WLA<251> B_WLA<250> B_WLA<249> B_WLA<248> B_WLA<247> 
+ B_WLA<246> B_WLA<245> B_WLA<244> B_WLA<243> B_WLA<242> B_WLA<241> B_WLA<240> B_WLA<239> B_WLA<238> 
+ B_WLA<237> B_WLA<236> B_WLA<235> B_WLA<234> B_WLA<233> B_WLA<232> B_WLA<231> B_WLA<230> B_WLA<229> 
+ B_WLA<228> B_WLA<227> B_WLA<226> B_WLA<225> B_WLA<224> B_WLA<223> B_WLA<222> B_WLA<221> B_WLA<220> 
+ B_WLA<219> B_WLA<218> B_WLA<217> B_WLA<216> B_WLA<215> B_WLA<214> B_WLA<213> B_WLA<212> B_WLA<211> 
+ B_WLA<210> B_WLA<209> B_WLA<208> B_WLA<207> B_WLA<206> B_WLA<205> B_WLA<204> B_WLA<203> B_WLA<202> 
+ B_WLA<201> B_WLA<200> B_WLA<199> B_WLA<198> B_WLA<197> B_WLA<196> B_WLA<195> B_WLA<194> B_WLA<193> 
+ B_WLA<192> B_WLA<191> B_WLA<190> B_WLA<189> B_WLA<188> B_WLA<187> B_WLA<186> B_WLA<185> B_WLA<184> 
+ B_WLA<183> B_WLA<182> B_WLA<181> B_WLA<180> B_WLA<179> B_WLA<178> B_WLA<177> B_WLA<176> B_WLA<175> 
+ B_WLA<174> B_WLA<173> B_WLA<172> B_WLA<171> B_WLA<170> B_WLA<169> B_WLA<168> B_WLA<167> B_WLA<166> 
+ B_WLA<165> B_WLA<164> B_WLA<163> B_WLA<162> B_WLA<161> B_WLA<160> B_WLA<159> B_WLA<158> B_WLA<157> 
+ B_WLA<156> B_WLA<155> B_WLA<154> B_WLA<153> B_WLA<152> B_WLA<151> B_WLA<150> B_WLA<149> B_WLA<148> 
+ B_WLA<147> B_WLA<146> B_WLA<145> B_WLA<144> B_WLA<143> B_WLA<142> B_WLA<141> B_WLA<140> B_WLA<139> 
+ B_WLA<138> B_WLA<137> B_WLA<136> B_WLA<135> B_WLA<134> B_WLA<133> B_WLA<132> B_WLA<131> B_WLA<130> 
+ B_WLA<129> B_WLA<128> B_WLA<127> B_WLA<126> B_WLA<125> B_WLA<124> B_WLA<123> B_WLA<122> B_WLA<121> 
+ B_WLA<120> B_WLA<119> B_WLA<118> B_WLA<117> B_WLA<116> B_WLA<115> B_WLA<114> B_WLA<113> B_WLA<112> 
+ B_WLA<111> B_WLA<110> B_WLA<109> B_WLA<108> B_WLA<107> B_WLA<106> B_WLA<105> B_WLA<104> B_WLA<103> 
+ B_WLA<102> B_WLA<101> B_WLA<100> B_WLA<99> B_WLA<98> B_WLA<97> B_WLA<96> B_WLA<95> B_WLA<94> 
+ B_WLA<93> B_WLA<92> B_WLA<91> B_WLA<90> B_WLA<89> B_WLA<88> B_WLA<87> B_WLA<86> B_WLA<85> 
+ B_WLA<84> B_WLA<83> B_WLA<82> B_WLA<81> B_WLA<80> B_WLA<79> B_WLA<78> B_WLA<77> B_WLA<76> 
+ B_WLA<75> B_WLA<74> B_WLA<73> B_WLA<72> B_WLA<71> B_WLA<70> B_WLA<69> B_WLA<68> B_WLA<67> 
+ B_WLA<66> B_WLA<65> B_WLA<64> B_WLA<63> B_WLA<62> B_WLA<61> B_WLA<60> B_WLA<59> B_WLA<58> 
+ B_WLA<57> B_WLA<56> B_WLA<55> B_WLA<54> B_WLA<53> B_WLA<52> B_WLA<51> B_WLA<50> B_WLA<49> 
+ B_WLA<48> B_WLA<47> B_WLA<46> B_WLA<45> B_WLA<44> B_WLA<43> B_WLA<42> B_WLA<41> B_WLA<40> 
+ B_WLA<39> B_WLA<38> B_WLA<37> B_WLA<36> B_WLA<35> B_WLA<34> B_WLA<33> B_WLA<32> B_WLA<31> 
+ B_WLA<30> B_WLA<29> B_WLA<28> B_WLA<27> B_WLA<26> B_WLA<25> B_WLA<24> B_WLA<23> B_WLA<22> 
+ B_WLA<21> B_WLA<20> B_WLA<19> B_WLA<18> B_WLA<17> B_WLA<16> B_WLA<15> B_WLA<14> B_WLA<13> 
+ B_WLA<12> B_WLA<11> B_WLA<10> B_WLA<9> B_WLA<8> B_WLA<7> B_WLA<6> B_WLA<5> B_WLA<4> 
+ B_WLA<3> B_WLA<2> B_WLA<1> B_WLA<0> B_WLB<255> B_WLB<254> B_WLB<253> B_WLB<252> B_WLB<251> 
+ B_WLB<250> B_WLB<249> B_WLB<248> B_WLB<247> B_WLB<246> B_WLB<245> B_WLB<244> B_WLB<243> B_WLB<242> 
+ B_WLB<241> B_WLB<240> B_WLB<239> B_WLB<238> B_WLB<237> B_WLB<236> B_WLB<235> B_WLB<234> B_WLB<233> 
+ B_WLB<232> B_WLB<231> B_WLB<230> B_WLB<229> B_WLB<228> B_WLB<227> B_WLB<226> B_WLB<225> B_WLB<224> 
+ B_WLB<223> B_WLB<222> B_WLB<221> B_WLB<220> B_WLB<219> B_WLB<218> B_WLB<217> B_WLB<216> B_WLB<215> 
+ B_WLB<214> B_WLB<213> B_WLB<212> B_WLB<211> B_WLB<210> B_WLB<209> B_WLB<208> B_WLB<207> B_WLB<206> 
+ B_WLB<205> B_WLB<204> B_WLB<203> B_WLB<202> B_WLB<201> B_WLB<200> B_WLB<199> B_WLB<198> B_WLB<197> 
+ B_WLB<196> B_WLB<195> B_WLB<194> B_WLB<193> B_WLB<192> B_WLB<191> B_WLB<190> B_WLB<189> B_WLB<188> 
+ B_WLB<187> B_WLB<186> B_WLB<185> B_WLB<184> B_WLB<183> B_WLB<182> B_WLB<181> B_WLB<180> B_WLB<179> 
+ B_WLB<178> B_WLB<177> B_WLB<176> B_WLB<175> B_WLB<174> B_WLB<173> B_WLB<172> B_WLB<171> B_WLB<170> 
+ B_WLB<169> B_WLB<168> B_WLB<167> B_WLB<166> B_WLB<165> B_WLB<164> B_WLB<163> B_WLB<162> B_WLB<161> 
+ B_WLB<160> B_WLB<159> B_WLB<158> B_WLB<157> B_WLB<156> B_WLB<155> B_WLB<154> B_WLB<153> B_WLB<152> 
+ B_WLB<151> B_WLB<150> B_WLB<149> B_WLB<148> B_WLB<147> B_WLB<146> B_WLB<145> B_WLB<144> B_WLB<143> 
+ B_WLB<142> B_WLB<141> B_WLB<140> B_WLB<139> B_WLB<138> B_WLB<137> B_WLB<136> B_WLB<135> B_WLB<134> 
+ B_WLB<133> B_WLB<132> B_WLB<131> B_WLB<130> B_WLB<129> B_WLB<128> B_WLB<127> B_WLB<126> B_WLB<125> 
+ B_WLB<124> B_WLB<123> B_WLB<122> B_WLB<121> B_WLB<120> B_WLB<119> B_WLB<118> B_WLB<117> B_WLB<116> 
+ B_WLB<115> B_WLB<114> B_WLB<113> B_WLB<112> B_WLB<111> B_WLB<110> B_WLB<109> B_WLB<108> B_WLB<107> 
+ B_WLB<106> B_WLB<105> B_WLB<104> B_WLB<103> B_WLB<102> B_WLB<101> B_WLB<100> B_WLB<99> B_WLB<98> 
+ B_WLB<97> B_WLB<96> B_WLB<95> B_WLB<94> B_WLB<93> B_WLB<92> B_WLB<91> B_WLB<90> B_WLB<89> 
+ B_WLB<88> B_WLB<87> B_WLB<86> B_WLB<85> B_WLB<84> B_WLB<83> B_WLB<82> B_WLB<81> B_WLB<80> 
+ B_WLB<79> B_WLB<78> B_WLB<77> B_WLB<76> B_WLB<75> B_WLB<74> B_WLB<73> B_WLB<72> B_WLB<71> 
+ B_WLB<70> B_WLB<69> B_WLB<68> B_WLB<67> B_WLB<66> B_WLB<65> B_WLB<64> B_WLB<63> B_WLB<62> 
+ B_WLB<61> B_WLB<60> B_WLB<59> B_WLB<58> B_WLB<57> B_WLB<56> B_WLB<55> B_WLB<54> B_WLB<53> 
+ B_WLB<52> B_WLB<51> B_WLB<50> B_WLB<49> B_WLB<48> B_WLB<47> B_WLB<46> B_WLB<45> B_WLB<44> 
+ B_WLB<43> B_WLB<42> B_WLB<41> B_WLB<40> B_WLB<39> B_WLB<38> B_WLB<37> B_WLB<36> B_WLB<35> 
+ B_WLB<34> B_WLB<33> B_WLB<32> B_WLB<31> B_WLB<30> B_WLB<29> B_WLB<28> B_WLB<27> B_WLB<26> 
+ B_WLB<25> B_WLB<24> B_WLB<23> B_WLB<22> B_WLB<21> B_WLB<20> B_WLB<19> B_WLB<18> B_WLB<17> 
+ B_WLB<16> B_WLB<15> B_WLB<14> B_WLB<13> B_WLB<12> B_WLB<11> B_WLB<10> B_WLB<9> B_WLB<8> 
+ B_WLB<7> B_WLB<6> B_WLB<5> B_WLB<4> B_WLB<3> B_WLB<2> B_WLB<1> B_WLB<0> BWENA<11> 
+ BWENA<10> BWENB<11> BWENB<10> L_CLK_DQA L_CLK_DQA_N L_CLK_DQB L_CLK_DQB_N DA<11> DA<10> 
+ DB<11> DB<10> DDQA<5> DDQA_N<5> DDQB<5> DDQB_N<5> L_LWEA L_LWEB QA<11> 
+ QA<10> QB<11> QB<10> L_SA_PREA_N L_SA_PREB_N L_SAEA_N L_SAEB_N LT_CA<3> LT_CA<2> 
+ LT_CA<1> LT_CA<0> LT_CB<3> LT_CB<2> LT_CB<1> LT_CB<0> LT_MA<3> LT_MA<2> LT_MA<1> 
+ LT_MA<0> LT_MB<3> LT_MB<2> LT_MB<1> LT_MB<0> LT_TM_PREA_N LT_TM_PREB_N T_WLA<255> T_WLA<254> 
+ T_WLA<253> T_WLA<252> T_WLA<251> T_WLA<250> T_WLA<249> T_WLA<248> T_WLA<247> T_WLA<246> T_WLA<245> 
+ T_WLA<244> T_WLA<243> T_WLA<242> T_WLA<241> T_WLA<240> T_WLA<239> T_WLA<238> T_WLA<237> T_WLA<236> 
+ T_WLA<235> T_WLA<234> T_WLA<233> T_WLA<232> T_WLA<231> T_WLA<230> T_WLA<229> T_WLA<228> T_WLA<227> 
+ T_WLA<226> T_WLA<225> T_WLA<224> T_WLA<223> T_WLA<222> T_WLA<221> T_WLA<220> T_WLA<219> T_WLA<218> 
+ T_WLA<217> T_WLA<216> T_WLA<215> T_WLA<214> T_WLA<213> T_WLA<212> T_WLA<211> T_WLA<210> T_WLA<209> 
+ T_WLA<208> T_WLA<207> T_WLA<206> T_WLA<205> T_WLA<204> T_WLA<203> T_WLA<202> T_WLA<201> T_WLA<200> 
+ T_WLA<199> T_WLA<198> T_WLA<197> T_WLA<196> T_WLA<195> T_WLA<194> T_WLA<193> T_WLA<192> T_WLA<191> 
+ T_WLA<190> T_WLA<189> T_WLA<188> T_WLA<187> T_WLA<186> T_WLA<185> T_WLA<184> T_WLA<183> T_WLA<182> 
+ T_WLA<181> T_WLA<180> T_WLA<179> T_WLA<178> T_WLA<177> T_WLA<176> T_WLA<175> T_WLA<174> T_WLA<173> 
+ T_WLA<172> T_WLA<171> T_WLA<170> T_WLA<169> T_WLA<168> T_WLA<167> T_WLA<166> T_WLA<165> T_WLA<164> 
+ T_WLA<163> T_WLA<162> T_WLA<161> T_WLA<160> T_WLA<159> T_WLA<158> T_WLA<157> T_WLA<156> T_WLA<155> 
+ T_WLA<154> T_WLA<153> T_WLA<152> T_WLA<151> T_WLA<150> T_WLA<149> T_WLA<148> T_WLA<147> T_WLA<146> 
+ T_WLA<145> T_WLA<144> T_WLA<143> T_WLA<142> T_WLA<141> T_WLA<140> T_WLA<139> T_WLA<138> T_WLA<137> 
+ T_WLA<136> T_WLA<135> T_WLA<134> T_WLA<133> T_WLA<132> T_WLA<131> T_WLA<130> T_WLA<129> T_WLA<128> 
+ T_WLA<127> T_WLA<126> T_WLA<125> T_WLA<124> T_WLA<123> T_WLA<122> T_WLA<121> T_WLA<120> T_WLA<119> 
+ T_WLA<118> T_WLA<117> T_WLA<116> T_WLA<115> T_WLA<114> T_WLA<113> T_WLA<112> T_WLA<111> T_WLA<110> 
+ T_WLA<109> T_WLA<108> T_WLA<107> T_WLA<106> T_WLA<105> T_WLA<104> T_WLA<103> T_WLA<102> T_WLA<101> 
+ T_WLA<100> T_WLA<99> T_WLA<98> T_WLA<97> T_WLA<96> T_WLA<95> T_WLA<94> T_WLA<93> T_WLA<92> 
+ T_WLA<91> T_WLA<90> T_WLA<89> T_WLA<88> T_WLA<87> T_WLA<86> T_WLA<85> T_WLA<84> T_WLA<83> 
+ T_WLA<82> T_WLA<81> T_WLA<80> T_WLA<79> T_WLA<78> T_WLA<77> T_WLA<76> T_WLA<75> T_WLA<74> 
+ T_WLA<73> T_WLA<72> T_WLA<71> T_WLA<70> T_WLA<69> T_WLA<68> T_WLA<67> T_WLA<66> T_WLA<65> 
+ T_WLA<64> T_WLA<63> T_WLA<62> T_WLA<61> T_WLA<60> T_WLA<59> T_WLA<58> T_WLA<57> T_WLA<56> 
+ T_WLA<55> T_WLA<54> T_WLA<53> T_WLA<52> T_WLA<51> T_WLA<50> T_WLA<49> T_WLA<48> T_WLA<47> 
+ T_WLA<46> T_WLA<45> T_WLA<44> T_WLA<43> T_WLA<42> T_WLA<41> T_WLA<40> T_WLA<39> T_WLA<38> 
+ T_WLA<37> T_WLA<36> T_WLA<35> T_WLA<34> T_WLA<33> T_WLA<32> T_WLA<31> T_WLA<30> T_WLA<29> 
+ T_WLA<28> T_WLA<27> T_WLA<26> T_WLA<25> T_WLA<24> T_WLA<23> T_WLA<22> T_WLA<21> T_WLA<20> 
+ T_WLA<19> T_WLA<18> T_WLA<17> T_WLA<16> T_WLA<15> T_WLA<14> T_WLA<13> T_WLA<12> T_WLA<11> 
+ T_WLA<10> T_WLA<9> T_WLA<8> T_WLA<7> T_WLA<6> T_WLA<5> T_WLA<4> T_WLA<3> T_WLA<2> 
+ T_WLA<1> T_WLA<0> T_WLB<255> T_WLB<254> T_WLB<253> T_WLB<252> T_WLB<251> T_WLB<250> T_WLB<249> 
+ T_WLB<248> T_WLB<247> T_WLB<246> T_WLB<245> T_WLB<244> T_WLB<243> T_WLB<242> T_WLB<241> T_WLB<240> 
+ T_WLB<239> T_WLB<238> T_WLB<237> T_WLB<236> T_WLB<235> T_WLB<234> T_WLB<233> T_WLB<232> T_WLB<231> 
+ T_WLB<230> T_WLB<229> T_WLB<228> T_WLB<227> T_WLB<226> T_WLB<225> T_WLB<224> T_WLB<223> T_WLB<222> 
+ T_WLB<221> T_WLB<220> T_WLB<219> T_WLB<218> T_WLB<217> T_WLB<216> T_WLB<215> T_WLB<214> T_WLB<213> 
+ T_WLB<212> T_WLB<211> T_WLB<210> T_WLB<209> T_WLB<208> T_WLB<207> T_WLB<206> T_WLB<205> T_WLB<204> 
+ T_WLB<203> T_WLB<202> T_WLB<201> T_WLB<200> T_WLB<199> T_WLB<198> T_WLB<197> T_WLB<196> T_WLB<195> 
+ T_WLB<194> T_WLB<193> T_WLB<192> T_WLB<191> T_WLB<190> T_WLB<189> T_WLB<188> T_WLB<187> T_WLB<186> 
+ T_WLB<185> T_WLB<184> T_WLB<183> T_WLB<182> T_WLB<181> T_WLB<180> T_WLB<179> T_WLB<178> T_WLB<177> 
+ T_WLB<176> T_WLB<175> T_WLB<174> T_WLB<173> T_WLB<172> T_WLB<171> T_WLB<170> T_WLB<169> T_WLB<168> 
+ T_WLB<167> T_WLB<166> T_WLB<165> T_WLB<164> T_WLB<163> T_WLB<162> T_WLB<161> T_WLB<160> T_WLB<159> 
+ T_WLB<158> T_WLB<157> T_WLB<156> T_WLB<155> T_WLB<154> T_WLB<153> T_WLB<152> T_WLB<151> T_WLB<150> 
+ T_WLB<149> T_WLB<148> T_WLB<147> T_WLB<146> T_WLB<145> T_WLB<144> T_WLB<143> T_WLB<142> T_WLB<141> 
+ T_WLB<140> T_WLB<139> T_WLB<138> T_WLB<137> T_WLB<136> T_WLB<135> T_WLB<134> T_WLB<133> T_WLB<132> 
+ T_WLB<131> T_WLB<130> T_WLB<129> T_WLB<128> T_WLB<127> T_WLB<126> T_WLB<125> T_WLB<124> T_WLB<123> 
+ T_WLB<122> T_WLB<121> T_WLB<120> T_WLB<119> T_WLB<118> T_WLB<117> T_WLB<116> T_WLB<115> T_WLB<114> 
+ T_WLB<113> T_WLB<112> T_WLB<111> T_WLB<110> T_WLB<109> T_WLB<108> T_WLB<107> T_WLB<106> T_WLB<105> 
+ T_WLB<104> T_WLB<103> T_WLB<102> T_WLB<101> T_WLB<100> T_WLB<99> T_WLB<98> T_WLB<97> T_WLB<96> 
+ T_WLB<95> T_WLB<94> T_WLB<93> T_WLB<92> T_WLB<91> T_WLB<90> T_WLB<89> T_WLB<88> T_WLB<87> 
+ T_WLB<86> T_WLB<85> T_WLB<84> T_WLB<83> T_WLB<82> T_WLB<81> T_WLB<80> T_WLB<79> T_WLB<78> 
+ T_WLB<77> T_WLB<76> T_WLB<75> T_WLB<74> T_WLB<73> T_WLB<72> T_WLB<71> T_WLB<70> T_WLB<69> 
+ T_WLB<68> T_WLB<67> T_WLB<66> T_WLB<65> T_WLB<64> T_WLB<63> T_WLB<62> T_WLB<61> T_WLB<60> 
+ T_WLB<59> T_WLB<58> T_WLB<57> T_WLB<56> T_WLB<55> T_WLB<54> T_WLB<53> T_WLB<52> T_WLB<51> 
+ T_WLB<50> T_WLB<49> T_WLB<48> T_WLB<47> T_WLB<46> T_WLB<45> T_WLB<44> T_WLB<43> T_WLB<42> 
+ T_WLB<41> T_WLB<40> T_WLB<39> T_WLB<38> T_WLB<37> T_WLB<36> T_WLB<35> T_WLB<34> T_WLB<33> 
+ T_WLB<32> T_WLB<31> T_WLB<30> T_WLB<29> T_WLB<28> T_WLB<27> T_WLB<26> T_WLB<25> T_WLB<24> 
+ T_WLB<23> T_WLB<22> T_WLB<21> T_WLB<20> T_WLB<19> T_WLB<18> T_WLB<17> T_WLB<16> T_WLB<15> 
+ T_WLB<14> T_WLB<13> T_WLB<12> T_WLB<11> T_WLB<10> T_WLB<9> T_WLB<8> T_WLB<7> T_WLB<6> 
+ T_WLB<5> T_WLB<4> T_WLB<3> T_WLB<2> T_WLB<1> T_WLB<0> VDD VSS  / dpram16x4096_SingleCOL2X8_ROWX256
XCOL2<4>
+ LB_CA<3> LB_CA<2> LB_CA<1> LB_CA<0> LB_CB<3> LB_CB<2> LB_CB<1> LB_CB<0> LB_MA<3> 
+ LB_MA<2> LB_MA<1> LB_MA<0> LB_MB<3> LB_MB<2> LB_MB<1> LB_MB<0> LB_TM_PREA_N LB_TM_PREB_N 
+ B_WLA<255> B_WLA<254> B_WLA<253> B_WLA<252> B_WLA<251> B_WLA<250> B_WLA<249> B_WLA<248> B_WLA<247> 
+ B_WLA<246> B_WLA<245> B_WLA<244> B_WLA<243> B_WLA<242> B_WLA<241> B_WLA<240> B_WLA<239> B_WLA<238> 
+ B_WLA<237> B_WLA<236> B_WLA<235> B_WLA<234> B_WLA<233> B_WLA<232> B_WLA<231> B_WLA<230> B_WLA<229> 
+ B_WLA<228> B_WLA<227> B_WLA<226> B_WLA<225> B_WLA<224> B_WLA<223> B_WLA<222> B_WLA<221> B_WLA<220> 
+ B_WLA<219> B_WLA<218> B_WLA<217> B_WLA<216> B_WLA<215> B_WLA<214> B_WLA<213> B_WLA<212> B_WLA<211> 
+ B_WLA<210> B_WLA<209> B_WLA<208> B_WLA<207> B_WLA<206> B_WLA<205> B_WLA<204> B_WLA<203> B_WLA<202> 
+ B_WLA<201> B_WLA<200> B_WLA<199> B_WLA<198> B_WLA<197> B_WLA<196> B_WLA<195> B_WLA<194> B_WLA<193> 
+ B_WLA<192> B_WLA<191> B_WLA<190> B_WLA<189> B_WLA<188> B_WLA<187> B_WLA<186> B_WLA<185> B_WLA<184> 
+ B_WLA<183> B_WLA<182> B_WLA<181> B_WLA<180> B_WLA<179> B_WLA<178> B_WLA<177> B_WLA<176> B_WLA<175> 
+ B_WLA<174> B_WLA<173> B_WLA<172> B_WLA<171> B_WLA<170> B_WLA<169> B_WLA<168> B_WLA<167> B_WLA<166> 
+ B_WLA<165> B_WLA<164> B_WLA<163> B_WLA<162> B_WLA<161> B_WLA<160> B_WLA<159> B_WLA<158> B_WLA<157> 
+ B_WLA<156> B_WLA<155> B_WLA<154> B_WLA<153> B_WLA<152> B_WLA<151> B_WLA<150> B_WLA<149> B_WLA<148> 
+ B_WLA<147> B_WLA<146> B_WLA<145> B_WLA<144> B_WLA<143> B_WLA<142> B_WLA<141> B_WLA<140> B_WLA<139> 
+ B_WLA<138> B_WLA<137> B_WLA<136> B_WLA<135> B_WLA<134> B_WLA<133> B_WLA<132> B_WLA<131> B_WLA<130> 
+ B_WLA<129> B_WLA<128> B_WLA<127> B_WLA<126> B_WLA<125> B_WLA<124> B_WLA<123> B_WLA<122> B_WLA<121> 
+ B_WLA<120> B_WLA<119> B_WLA<118> B_WLA<117> B_WLA<116> B_WLA<115> B_WLA<114> B_WLA<113> B_WLA<112> 
+ B_WLA<111> B_WLA<110> B_WLA<109> B_WLA<108> B_WLA<107> B_WLA<106> B_WLA<105> B_WLA<104> B_WLA<103> 
+ B_WLA<102> B_WLA<101> B_WLA<100> B_WLA<99> B_WLA<98> B_WLA<97> B_WLA<96> B_WLA<95> B_WLA<94> 
+ B_WLA<93> B_WLA<92> B_WLA<91> B_WLA<90> B_WLA<89> B_WLA<88> B_WLA<87> B_WLA<86> B_WLA<85> 
+ B_WLA<84> B_WLA<83> B_WLA<82> B_WLA<81> B_WLA<80> B_WLA<79> B_WLA<78> B_WLA<77> B_WLA<76> 
+ B_WLA<75> B_WLA<74> B_WLA<73> B_WLA<72> B_WLA<71> B_WLA<70> B_WLA<69> B_WLA<68> B_WLA<67> 
+ B_WLA<66> B_WLA<65> B_WLA<64> B_WLA<63> B_WLA<62> B_WLA<61> B_WLA<60> B_WLA<59> B_WLA<58> 
+ B_WLA<57> B_WLA<56> B_WLA<55> B_WLA<54> B_WLA<53> B_WLA<52> B_WLA<51> B_WLA<50> B_WLA<49> 
+ B_WLA<48> B_WLA<47> B_WLA<46> B_WLA<45> B_WLA<44> B_WLA<43> B_WLA<42> B_WLA<41> B_WLA<40> 
+ B_WLA<39> B_WLA<38> B_WLA<37> B_WLA<36> B_WLA<35> B_WLA<34> B_WLA<33> B_WLA<32> B_WLA<31> 
+ B_WLA<30> B_WLA<29> B_WLA<28> B_WLA<27> B_WLA<26> B_WLA<25> B_WLA<24> B_WLA<23> B_WLA<22> 
+ B_WLA<21> B_WLA<20> B_WLA<19> B_WLA<18> B_WLA<17> B_WLA<16> B_WLA<15> B_WLA<14> B_WLA<13> 
+ B_WLA<12> B_WLA<11> B_WLA<10> B_WLA<9> B_WLA<8> B_WLA<7> B_WLA<6> B_WLA<5> B_WLA<4> 
+ B_WLA<3> B_WLA<2> B_WLA<1> B_WLA<0> B_WLB<255> B_WLB<254> B_WLB<253> B_WLB<252> B_WLB<251> 
+ B_WLB<250> B_WLB<249> B_WLB<248> B_WLB<247> B_WLB<246> B_WLB<245> B_WLB<244> B_WLB<243> B_WLB<242> 
+ B_WLB<241> B_WLB<240> B_WLB<239> B_WLB<238> B_WLB<237> B_WLB<236> B_WLB<235> B_WLB<234> B_WLB<233> 
+ B_WLB<232> B_WLB<231> B_WLB<230> B_WLB<229> B_WLB<228> B_WLB<227> B_WLB<226> B_WLB<225> B_WLB<224> 
+ B_WLB<223> B_WLB<222> B_WLB<221> B_WLB<220> B_WLB<219> B_WLB<218> B_WLB<217> B_WLB<216> B_WLB<215> 
+ B_WLB<214> B_WLB<213> B_WLB<212> B_WLB<211> B_WLB<210> B_WLB<209> B_WLB<208> B_WLB<207> B_WLB<206> 
+ B_WLB<205> B_WLB<204> B_WLB<203> B_WLB<202> B_WLB<201> B_WLB<200> B_WLB<199> B_WLB<198> B_WLB<197> 
+ B_WLB<196> B_WLB<195> B_WLB<194> B_WLB<193> B_WLB<192> B_WLB<191> B_WLB<190> B_WLB<189> B_WLB<188> 
+ B_WLB<187> B_WLB<186> B_WLB<185> B_WLB<184> B_WLB<183> B_WLB<182> B_WLB<181> B_WLB<180> B_WLB<179> 
+ B_WLB<178> B_WLB<177> B_WLB<176> B_WLB<175> B_WLB<174> B_WLB<173> B_WLB<172> B_WLB<171> B_WLB<170> 
+ B_WLB<169> B_WLB<168> B_WLB<167> B_WLB<166> B_WLB<165> B_WLB<164> B_WLB<163> B_WLB<162> B_WLB<161> 
+ B_WLB<160> B_WLB<159> B_WLB<158> B_WLB<157> B_WLB<156> B_WLB<155> B_WLB<154> B_WLB<153> B_WLB<152> 
+ B_WLB<151> B_WLB<150> B_WLB<149> B_WLB<148> B_WLB<147> B_WLB<146> B_WLB<145> B_WLB<144> B_WLB<143> 
+ B_WLB<142> B_WLB<141> B_WLB<140> B_WLB<139> B_WLB<138> B_WLB<137> B_WLB<136> B_WLB<135> B_WLB<134> 
+ B_WLB<133> B_WLB<132> B_WLB<131> B_WLB<130> B_WLB<129> B_WLB<128> B_WLB<127> B_WLB<126> B_WLB<125> 
+ B_WLB<124> B_WLB<123> B_WLB<122> B_WLB<121> B_WLB<120> B_WLB<119> B_WLB<118> B_WLB<117> B_WLB<116> 
+ B_WLB<115> B_WLB<114> B_WLB<113> B_WLB<112> B_WLB<111> B_WLB<110> B_WLB<109> B_WLB<108> B_WLB<107> 
+ B_WLB<106> B_WLB<105> B_WLB<104> B_WLB<103> B_WLB<102> B_WLB<101> B_WLB<100> B_WLB<99> B_WLB<98> 
+ B_WLB<97> B_WLB<96> B_WLB<95> B_WLB<94> B_WLB<93> B_WLB<92> B_WLB<91> B_WLB<90> B_WLB<89> 
+ B_WLB<88> B_WLB<87> B_WLB<86> B_WLB<85> B_WLB<84> B_WLB<83> B_WLB<82> B_WLB<81> B_WLB<80> 
+ B_WLB<79> B_WLB<78> B_WLB<77> B_WLB<76> B_WLB<75> B_WLB<74> B_WLB<73> B_WLB<72> B_WLB<71> 
+ B_WLB<70> B_WLB<69> B_WLB<68> B_WLB<67> B_WLB<66> B_WLB<65> B_WLB<64> B_WLB<63> B_WLB<62> 
+ B_WLB<61> B_WLB<60> B_WLB<59> B_WLB<58> B_WLB<57> B_WLB<56> B_WLB<55> B_WLB<54> B_WLB<53> 
+ B_WLB<52> B_WLB<51> B_WLB<50> B_WLB<49> B_WLB<48> B_WLB<47> B_WLB<46> B_WLB<45> B_WLB<44> 
+ B_WLB<43> B_WLB<42> B_WLB<41> B_WLB<40> B_WLB<39> B_WLB<38> B_WLB<37> B_WLB<36> B_WLB<35> 
+ B_WLB<34> B_WLB<33> B_WLB<32> B_WLB<31> B_WLB<30> B_WLB<29> B_WLB<28> B_WLB<27> B_WLB<26> 
+ B_WLB<25> B_WLB<24> B_WLB<23> B_WLB<22> B_WLB<21> B_WLB<20> B_WLB<19> B_WLB<18> B_WLB<17> 
+ B_WLB<16> B_WLB<15> B_WLB<14> B_WLB<13> B_WLB<12> B_WLB<11> B_WLB<10> B_WLB<9> B_WLB<8> 
+ B_WLB<7> B_WLB<6> B_WLB<5> B_WLB<4> B_WLB<3> B_WLB<2> B_WLB<1> B_WLB<0> BWENA<9> 
+ BWENA<8> BWENB<9> BWENB<8> L_CLK_DQA L_CLK_DQA_N L_CLK_DQB L_CLK_DQB_N DA<9> DA<8> 
+ DB<9> DB<8> DDQA<4> DDQA_N<4> DDQB<4> DDQB_N<4> L_LWEA L_LWEB QA<9> 
+ QA<8> QB<9> QB<8> L_SA_PREA_N L_SA_PREB_N L_SAEA_N L_SAEB_N LT_CA<3> LT_CA<2> 
+ LT_CA<1> LT_CA<0> LT_CB<3> LT_CB<2> LT_CB<1> LT_CB<0> LT_MA<3> LT_MA<2> LT_MA<1> 
+ LT_MA<0> LT_MB<3> LT_MB<2> LT_MB<1> LT_MB<0> LT_TM_PREA_N LT_TM_PREB_N T_WLA<255> T_WLA<254> 
+ T_WLA<253> T_WLA<252> T_WLA<251> T_WLA<250> T_WLA<249> T_WLA<248> T_WLA<247> T_WLA<246> T_WLA<245> 
+ T_WLA<244> T_WLA<243> T_WLA<242> T_WLA<241> T_WLA<240> T_WLA<239> T_WLA<238> T_WLA<237> T_WLA<236> 
+ T_WLA<235> T_WLA<234> T_WLA<233> T_WLA<232> T_WLA<231> T_WLA<230> T_WLA<229> T_WLA<228> T_WLA<227> 
+ T_WLA<226> T_WLA<225> T_WLA<224> T_WLA<223> T_WLA<222> T_WLA<221> T_WLA<220> T_WLA<219> T_WLA<218> 
+ T_WLA<217> T_WLA<216> T_WLA<215> T_WLA<214> T_WLA<213> T_WLA<212> T_WLA<211> T_WLA<210> T_WLA<209> 
+ T_WLA<208> T_WLA<207> T_WLA<206> T_WLA<205> T_WLA<204> T_WLA<203> T_WLA<202> T_WLA<201> T_WLA<200> 
+ T_WLA<199> T_WLA<198> T_WLA<197> T_WLA<196> T_WLA<195> T_WLA<194> T_WLA<193> T_WLA<192> T_WLA<191> 
+ T_WLA<190> T_WLA<189> T_WLA<188> T_WLA<187> T_WLA<186> T_WLA<185> T_WLA<184> T_WLA<183> T_WLA<182> 
+ T_WLA<181> T_WLA<180> T_WLA<179> T_WLA<178> T_WLA<177> T_WLA<176> T_WLA<175> T_WLA<174> T_WLA<173> 
+ T_WLA<172> T_WLA<171> T_WLA<170> T_WLA<169> T_WLA<168> T_WLA<167> T_WLA<166> T_WLA<165> T_WLA<164> 
+ T_WLA<163> T_WLA<162> T_WLA<161> T_WLA<160> T_WLA<159> T_WLA<158> T_WLA<157> T_WLA<156> T_WLA<155> 
+ T_WLA<154> T_WLA<153> T_WLA<152> T_WLA<151> T_WLA<150> T_WLA<149> T_WLA<148> T_WLA<147> T_WLA<146> 
+ T_WLA<145> T_WLA<144> T_WLA<143> T_WLA<142> T_WLA<141> T_WLA<140> T_WLA<139> T_WLA<138> T_WLA<137> 
+ T_WLA<136> T_WLA<135> T_WLA<134> T_WLA<133> T_WLA<132> T_WLA<131> T_WLA<130> T_WLA<129> T_WLA<128> 
+ T_WLA<127> T_WLA<126> T_WLA<125> T_WLA<124> T_WLA<123> T_WLA<122> T_WLA<121> T_WLA<120> T_WLA<119> 
+ T_WLA<118> T_WLA<117> T_WLA<116> T_WLA<115> T_WLA<114> T_WLA<113> T_WLA<112> T_WLA<111> T_WLA<110> 
+ T_WLA<109> T_WLA<108> T_WLA<107> T_WLA<106> T_WLA<105> T_WLA<104> T_WLA<103> T_WLA<102> T_WLA<101> 
+ T_WLA<100> T_WLA<99> T_WLA<98> T_WLA<97> T_WLA<96> T_WLA<95> T_WLA<94> T_WLA<93> T_WLA<92> 
+ T_WLA<91> T_WLA<90> T_WLA<89> T_WLA<88> T_WLA<87> T_WLA<86> T_WLA<85> T_WLA<84> T_WLA<83> 
+ T_WLA<82> T_WLA<81> T_WLA<80> T_WLA<79> T_WLA<78> T_WLA<77> T_WLA<76> T_WLA<75> T_WLA<74> 
+ T_WLA<73> T_WLA<72> T_WLA<71> T_WLA<70> T_WLA<69> T_WLA<68> T_WLA<67> T_WLA<66> T_WLA<65> 
+ T_WLA<64> T_WLA<63> T_WLA<62> T_WLA<61> T_WLA<60> T_WLA<59> T_WLA<58> T_WLA<57> T_WLA<56> 
+ T_WLA<55> T_WLA<54> T_WLA<53> T_WLA<52> T_WLA<51> T_WLA<50> T_WLA<49> T_WLA<48> T_WLA<47> 
+ T_WLA<46> T_WLA<45> T_WLA<44> T_WLA<43> T_WLA<42> T_WLA<41> T_WLA<40> T_WLA<39> T_WLA<38> 
+ T_WLA<37> T_WLA<36> T_WLA<35> T_WLA<34> T_WLA<33> T_WLA<32> T_WLA<31> T_WLA<30> T_WLA<29> 
+ T_WLA<28> T_WLA<27> T_WLA<26> T_WLA<25> T_WLA<24> T_WLA<23> T_WLA<22> T_WLA<21> T_WLA<20> 
+ T_WLA<19> T_WLA<18> T_WLA<17> T_WLA<16> T_WLA<15> T_WLA<14> T_WLA<13> T_WLA<12> T_WLA<11> 
+ T_WLA<10> T_WLA<9> T_WLA<8> T_WLA<7> T_WLA<6> T_WLA<5> T_WLA<4> T_WLA<3> T_WLA<2> 
+ T_WLA<1> T_WLA<0> T_WLB<255> T_WLB<254> T_WLB<253> T_WLB<252> T_WLB<251> T_WLB<250> T_WLB<249> 
+ T_WLB<248> T_WLB<247> T_WLB<246> T_WLB<245> T_WLB<244> T_WLB<243> T_WLB<242> T_WLB<241> T_WLB<240> 
+ T_WLB<239> T_WLB<238> T_WLB<237> T_WLB<236> T_WLB<235> T_WLB<234> T_WLB<233> T_WLB<232> T_WLB<231> 
+ T_WLB<230> T_WLB<229> T_WLB<228> T_WLB<227> T_WLB<226> T_WLB<225> T_WLB<224> T_WLB<223> T_WLB<222> 
+ T_WLB<221> T_WLB<220> T_WLB<219> T_WLB<218> T_WLB<217> T_WLB<216> T_WLB<215> T_WLB<214> T_WLB<213> 
+ T_WLB<212> T_WLB<211> T_WLB<210> T_WLB<209> T_WLB<208> T_WLB<207> T_WLB<206> T_WLB<205> T_WLB<204> 
+ T_WLB<203> T_WLB<202> T_WLB<201> T_WLB<200> T_WLB<199> T_WLB<198> T_WLB<197> T_WLB<196> T_WLB<195> 
+ T_WLB<194> T_WLB<193> T_WLB<192> T_WLB<191> T_WLB<190> T_WLB<189> T_WLB<188> T_WLB<187> T_WLB<186> 
+ T_WLB<185> T_WLB<184> T_WLB<183> T_WLB<182> T_WLB<181> T_WLB<180> T_WLB<179> T_WLB<178> T_WLB<177> 
+ T_WLB<176> T_WLB<175> T_WLB<174> T_WLB<173> T_WLB<172> T_WLB<171> T_WLB<170> T_WLB<169> T_WLB<168> 
+ T_WLB<167> T_WLB<166> T_WLB<165> T_WLB<164> T_WLB<163> T_WLB<162> T_WLB<161> T_WLB<160> T_WLB<159> 
+ T_WLB<158> T_WLB<157> T_WLB<156> T_WLB<155> T_WLB<154> T_WLB<153> T_WLB<152> T_WLB<151> T_WLB<150> 
+ T_WLB<149> T_WLB<148> T_WLB<147> T_WLB<146> T_WLB<145> T_WLB<144> T_WLB<143> T_WLB<142> T_WLB<141> 
+ T_WLB<140> T_WLB<139> T_WLB<138> T_WLB<137> T_WLB<136> T_WLB<135> T_WLB<134> T_WLB<133> T_WLB<132> 
+ T_WLB<131> T_WLB<130> T_WLB<129> T_WLB<128> T_WLB<127> T_WLB<126> T_WLB<125> T_WLB<124> T_WLB<123> 
+ T_WLB<122> T_WLB<121> T_WLB<120> T_WLB<119> T_WLB<118> T_WLB<117> T_WLB<116> T_WLB<115> T_WLB<114> 
+ T_WLB<113> T_WLB<112> T_WLB<111> T_WLB<110> T_WLB<109> T_WLB<108> T_WLB<107> T_WLB<106> T_WLB<105> 
+ T_WLB<104> T_WLB<103> T_WLB<102> T_WLB<101> T_WLB<100> T_WLB<99> T_WLB<98> T_WLB<97> T_WLB<96> 
+ T_WLB<95> T_WLB<94> T_WLB<93> T_WLB<92> T_WLB<91> T_WLB<90> T_WLB<89> T_WLB<88> T_WLB<87> 
+ T_WLB<86> T_WLB<85> T_WLB<84> T_WLB<83> T_WLB<82> T_WLB<81> T_WLB<80> T_WLB<79> T_WLB<78> 
+ T_WLB<77> T_WLB<76> T_WLB<75> T_WLB<74> T_WLB<73> T_WLB<72> T_WLB<71> T_WLB<70> T_WLB<69> 
+ T_WLB<68> T_WLB<67> T_WLB<66> T_WLB<65> T_WLB<64> T_WLB<63> T_WLB<62> T_WLB<61> T_WLB<60> 
+ T_WLB<59> T_WLB<58> T_WLB<57> T_WLB<56> T_WLB<55> T_WLB<54> T_WLB<53> T_WLB<52> T_WLB<51> 
+ T_WLB<50> T_WLB<49> T_WLB<48> T_WLB<47> T_WLB<46> T_WLB<45> T_WLB<44> T_WLB<43> T_WLB<42> 
+ T_WLB<41> T_WLB<40> T_WLB<39> T_WLB<38> T_WLB<37> T_WLB<36> T_WLB<35> T_WLB<34> T_WLB<33> 
+ T_WLB<32> T_WLB<31> T_WLB<30> T_WLB<29> T_WLB<28> T_WLB<27> T_WLB<26> T_WLB<25> T_WLB<24> 
+ T_WLB<23> T_WLB<22> T_WLB<21> T_WLB<20> T_WLB<19> T_WLB<18> T_WLB<17> T_WLB<16> T_WLB<15> 
+ T_WLB<14> T_WLB<13> T_WLB<12> T_WLB<11> T_WLB<10> T_WLB<9> T_WLB<8> T_WLB<7> T_WLB<6> 
+ T_WLB<5> T_WLB<4> T_WLB<3> T_WLB<2> T_WLB<1> T_WLB<0> VDD VSS  / dpram16x4096_SingleCOL2X8_ROWX256
XCOL2<3>
+ RB_CA<3> RB_CA<2> RB_CA<1> RB_CA<0> RB_CB<3> RB_CB<2> RB_CB<1> RB_CB<0> RB_MA<3> 
+ RB_MA<2> RB_MA<1> RB_MA<0> RB_MB<3> RB_MB<2> RB_MB<1> RB_MB<0> RB_TM_PREB_N RB_TM_PREA_N 
+ B_WLA<255> B_WLA<254> B_WLA<253> B_WLA<252> B_WLA<251> B_WLA<250> B_WLA<249> B_WLA<248> B_WLA<247> 
+ B_WLA<246> B_WLA<245> B_WLA<244> B_WLA<243> B_WLA<242> B_WLA<241> B_WLA<240> B_WLA<239> B_WLA<238> 
+ B_WLA<237> B_WLA<236> B_WLA<235> B_WLA<234> B_WLA<233> B_WLA<232> B_WLA<231> B_WLA<230> B_WLA<229> 
+ B_WLA<228> B_WLA<227> B_WLA<226> B_WLA<225> B_WLA<224> B_WLA<223> B_WLA<222> B_WLA<221> B_WLA<220> 
+ B_WLA<219> B_WLA<218> B_WLA<217> B_WLA<216> B_WLA<215> B_WLA<214> B_WLA<213> B_WLA<212> B_WLA<211> 
+ B_WLA<210> B_WLA<209> B_WLA<208> B_WLA<207> B_WLA<206> B_WLA<205> B_WLA<204> B_WLA<203> B_WLA<202> 
+ B_WLA<201> B_WLA<200> B_WLA<199> B_WLA<198> B_WLA<197> B_WLA<196> B_WLA<195> B_WLA<194> B_WLA<193> 
+ B_WLA<192> B_WLA<191> B_WLA<190> B_WLA<189> B_WLA<188> B_WLA<187> B_WLA<186> B_WLA<185> B_WLA<184> 
+ B_WLA<183> B_WLA<182> B_WLA<181> B_WLA<180> B_WLA<179> B_WLA<178> B_WLA<177> B_WLA<176> B_WLA<175> 
+ B_WLA<174> B_WLA<173> B_WLA<172> B_WLA<171> B_WLA<170> B_WLA<169> B_WLA<168> B_WLA<167> B_WLA<166> 
+ B_WLA<165> B_WLA<164> B_WLA<163> B_WLA<162> B_WLA<161> B_WLA<160> B_WLA<159> B_WLA<158> B_WLA<157> 
+ B_WLA<156> B_WLA<155> B_WLA<154> B_WLA<153> B_WLA<152> B_WLA<151> B_WLA<150> B_WLA<149> B_WLA<148> 
+ B_WLA<147> B_WLA<146> B_WLA<145> B_WLA<144> B_WLA<143> B_WLA<142> B_WLA<141> B_WLA<140> B_WLA<139> 
+ B_WLA<138> B_WLA<137> B_WLA<136> B_WLA<135> B_WLA<134> B_WLA<133> B_WLA<132> B_WLA<131> B_WLA<130> 
+ B_WLA<129> B_WLA<128> B_WLA<127> B_WLA<126> B_WLA<125> B_WLA<124> B_WLA<123> B_WLA<122> B_WLA<121> 
+ B_WLA<120> B_WLA<119> B_WLA<118> B_WLA<117> B_WLA<116> B_WLA<115> B_WLA<114> B_WLA<113> B_WLA<112> 
+ B_WLA<111> B_WLA<110> B_WLA<109> B_WLA<108> B_WLA<107> B_WLA<106> B_WLA<105> B_WLA<104> B_WLA<103> 
+ B_WLA<102> B_WLA<101> B_WLA<100> B_WLA<99> B_WLA<98> B_WLA<97> B_WLA<96> B_WLA<95> B_WLA<94> 
+ B_WLA<93> B_WLA<92> B_WLA<91> B_WLA<90> B_WLA<89> B_WLA<88> B_WLA<87> B_WLA<86> B_WLA<85> 
+ B_WLA<84> B_WLA<83> B_WLA<82> B_WLA<81> B_WLA<80> B_WLA<79> B_WLA<78> B_WLA<77> B_WLA<76> 
+ B_WLA<75> B_WLA<74> B_WLA<73> B_WLA<72> B_WLA<71> B_WLA<70> B_WLA<69> B_WLA<68> B_WLA<67> 
+ B_WLA<66> B_WLA<65> B_WLA<64> B_WLA<63> B_WLA<62> B_WLA<61> B_WLA<60> B_WLA<59> B_WLA<58> 
+ B_WLA<57> B_WLA<56> B_WLA<55> B_WLA<54> B_WLA<53> B_WLA<52> B_WLA<51> B_WLA<50> B_WLA<49> 
+ B_WLA<48> B_WLA<47> B_WLA<46> B_WLA<45> B_WLA<44> B_WLA<43> B_WLA<42> B_WLA<41> B_WLA<40> 
+ B_WLA<39> B_WLA<38> B_WLA<37> B_WLA<36> B_WLA<35> B_WLA<34> B_WLA<33> B_WLA<32> B_WLA<31> 
+ B_WLA<30> B_WLA<29> B_WLA<28> B_WLA<27> B_WLA<26> B_WLA<25> B_WLA<24> B_WLA<23> B_WLA<22> 
+ B_WLA<21> B_WLA<20> B_WLA<19> B_WLA<18> B_WLA<17> B_WLA<16> B_WLA<15> B_WLA<14> B_WLA<13> 
+ B_WLA<12> B_WLA<11> B_WLA<10> B_WLA<9> B_WLA<8> B_WLA<7> B_WLA<6> B_WLA<5> B_WLA<4> 
+ B_WLA<3> B_WLA<2> B_WLA<1> B_WLA<0> B_WLB<255> B_WLB<254> B_WLB<253> B_WLB<252> B_WLB<251> 
+ B_WLB<250> B_WLB<249> B_WLB<248> B_WLB<247> B_WLB<246> B_WLB<245> B_WLB<244> B_WLB<243> B_WLB<242> 
+ B_WLB<241> B_WLB<240> B_WLB<239> B_WLB<238> B_WLB<237> B_WLB<236> B_WLB<235> B_WLB<234> B_WLB<233> 
+ B_WLB<232> B_WLB<231> B_WLB<230> B_WLB<229> B_WLB<228> B_WLB<227> B_WLB<226> B_WLB<225> B_WLB<224> 
+ B_WLB<223> B_WLB<222> B_WLB<221> B_WLB<220> B_WLB<219> B_WLB<218> B_WLB<217> B_WLB<216> B_WLB<215> 
+ B_WLB<214> B_WLB<213> B_WLB<212> B_WLB<211> B_WLB<210> B_WLB<209> B_WLB<208> B_WLB<207> B_WLB<206> 
+ B_WLB<205> B_WLB<204> B_WLB<203> B_WLB<202> B_WLB<201> B_WLB<200> B_WLB<199> B_WLB<198> B_WLB<197> 
+ B_WLB<196> B_WLB<195> B_WLB<194> B_WLB<193> B_WLB<192> B_WLB<191> B_WLB<190> B_WLB<189> B_WLB<188> 
+ B_WLB<187> B_WLB<186> B_WLB<185> B_WLB<184> B_WLB<183> B_WLB<182> B_WLB<181> B_WLB<180> B_WLB<179> 
+ B_WLB<178> B_WLB<177> B_WLB<176> B_WLB<175> B_WLB<174> B_WLB<173> B_WLB<172> B_WLB<171> B_WLB<170> 
+ B_WLB<169> B_WLB<168> B_WLB<167> B_WLB<166> B_WLB<165> B_WLB<164> B_WLB<163> B_WLB<162> B_WLB<161> 
+ B_WLB<160> B_WLB<159> B_WLB<158> B_WLB<157> B_WLB<156> B_WLB<155> B_WLB<154> B_WLB<153> B_WLB<152> 
+ B_WLB<151> B_WLB<150> B_WLB<149> B_WLB<148> B_WLB<147> B_WLB<146> B_WLB<145> B_WLB<144> B_WLB<143> 
+ B_WLB<142> B_WLB<141> B_WLB<140> B_WLB<139> B_WLB<138> B_WLB<137> B_WLB<136> B_WLB<135> B_WLB<134> 
+ B_WLB<133> B_WLB<132> B_WLB<131> B_WLB<130> B_WLB<129> B_WLB<128> B_WLB<127> B_WLB<126> B_WLB<125> 
+ B_WLB<124> B_WLB<123> B_WLB<122> B_WLB<121> B_WLB<120> B_WLB<119> B_WLB<118> B_WLB<117> B_WLB<116> 
+ B_WLB<115> B_WLB<114> B_WLB<113> B_WLB<112> B_WLB<111> B_WLB<110> B_WLB<109> B_WLB<108> B_WLB<107> 
+ B_WLB<106> B_WLB<105> B_WLB<104> B_WLB<103> B_WLB<102> B_WLB<101> B_WLB<100> B_WLB<99> B_WLB<98> 
+ B_WLB<97> B_WLB<96> B_WLB<95> B_WLB<94> B_WLB<93> B_WLB<92> B_WLB<91> B_WLB<90> B_WLB<89> 
+ B_WLB<88> B_WLB<87> B_WLB<86> B_WLB<85> B_WLB<84> B_WLB<83> B_WLB<82> B_WLB<81> B_WLB<80> 
+ B_WLB<79> B_WLB<78> B_WLB<77> B_WLB<76> B_WLB<75> B_WLB<74> B_WLB<73> B_WLB<72> B_WLB<71> 
+ B_WLB<70> B_WLB<69> B_WLB<68> B_WLB<67> B_WLB<66> B_WLB<65> B_WLB<64> B_WLB<63> B_WLB<62> 
+ B_WLB<61> B_WLB<60> B_WLB<59> B_WLB<58> B_WLB<57> B_WLB<56> B_WLB<55> B_WLB<54> B_WLB<53> 
+ B_WLB<52> B_WLB<51> B_WLB<50> B_WLB<49> B_WLB<48> B_WLB<47> B_WLB<46> B_WLB<45> B_WLB<44> 
+ B_WLB<43> B_WLB<42> B_WLB<41> B_WLB<40> B_WLB<39> B_WLB<38> B_WLB<37> B_WLB<36> B_WLB<35> 
+ B_WLB<34> B_WLB<33> B_WLB<32> B_WLB<31> B_WLB<30> B_WLB<29> B_WLB<28> B_WLB<27> B_WLB<26> 
+ B_WLB<25> B_WLB<24> B_WLB<23> B_WLB<22> B_WLB<21> B_WLB<20> B_WLB<19> B_WLB<18> B_WLB<17> 
+ B_WLB<16> B_WLB<15> B_WLB<14> B_WLB<13> B_WLB<12> B_WLB<11> B_WLB<10> B_WLB<9> B_WLB<8> 
+ B_WLB<7> B_WLB<6> B_WLB<5> B_WLB<4> B_WLB<3> B_WLB<2> B_WLB<1> B_WLB<0> BWENA<7> 
+ BWENA<6> BWENB<7> BWENB<6> R_CLK_DQA R_CLK_DQA_N R_CLK_DQB R_CLK_DQB_N DA<7> DA<6> 
+ DB<7> DB<6> DDQA<3> DDQA_N<3> DDQB<3> DDQB_N<3> R_LWEA R_LWEB QA<7> 
+ QA<6> QB<7> QB<6> R_SA_PREA_N R_SA_PREB_N R_SAEA_N R_SAEB_N RT_CA<3> RT_CA<2> 
+ RT_CA<1> RT_CA<0> RT_CB<3> RT_CB<2> RT_CB<1> RT_CB<0> RT_MA<3> RT_MA<2> RT_MA<1> 
+ RT_MA<0> RT_MB<3> RT_MB<2> RT_MB<1> RT_MB<0> R_TM_PREA_N R_TM_PREB_N T_WLA<255> T_WLA<254> 
+ T_WLA<253> T_WLA<252> T_WLA<251> T_WLA<250> T_WLA<249> T_WLA<248> T_WLA<247> T_WLA<246> T_WLA<245> 
+ T_WLA<244> T_WLA<243> T_WLA<242> T_WLA<241> T_WLA<240> T_WLA<239> T_WLA<238> T_WLA<237> T_WLA<236> 
+ T_WLA<235> T_WLA<234> T_WLA<233> T_WLA<232> T_WLA<231> T_WLA<230> T_WLA<229> T_WLA<228> T_WLA<227> 
+ T_WLA<226> T_WLA<225> T_WLA<224> T_WLA<223> T_WLA<222> T_WLA<221> T_WLA<220> T_WLA<219> T_WLA<218> 
+ T_WLA<217> T_WLA<216> T_WLA<215> T_WLA<214> T_WLA<213> T_WLA<212> T_WLA<211> T_WLA<210> T_WLA<209> 
+ T_WLA<208> T_WLA<207> T_WLA<206> T_WLA<205> T_WLA<204> T_WLA<203> T_WLA<202> T_WLA<201> T_WLA<200> 
+ T_WLA<199> T_WLA<198> T_WLA<197> T_WLA<196> T_WLA<195> T_WLA<194> T_WLA<193> T_WLA<192> T_WLA<191> 
+ T_WLA<190> T_WLA<189> T_WLA<188> T_WLA<187> T_WLA<186> T_WLA<185> T_WLA<184> T_WLA<183> T_WLA<182> 
+ T_WLA<181> T_WLA<180> T_WLA<179> T_WLA<178> T_WLA<177> T_WLA<176> T_WLA<175> T_WLA<174> T_WLA<173> 
+ T_WLA<172> T_WLA<171> T_WLA<170> T_WLA<169> T_WLA<168> T_WLA<167> T_WLA<166> T_WLA<165> T_WLA<164> 
+ T_WLA<163> T_WLA<162> T_WLA<161> T_WLA<160> T_WLA<159> T_WLA<158> T_WLA<157> T_WLA<156> T_WLA<155> 
+ T_WLA<154> T_WLA<153> T_WLA<152> T_WLA<151> T_WLA<150> T_WLA<149> T_WLA<148> T_WLA<147> T_WLA<146> 
+ T_WLA<145> T_WLA<144> T_WLA<143> T_WLA<142> T_WLA<141> T_WLA<140> T_WLA<139> T_WLA<138> T_WLA<137> 
+ T_WLA<136> T_WLA<135> T_WLA<134> T_WLA<133> T_WLA<132> T_WLA<131> T_WLA<130> T_WLA<129> T_WLA<128> 
+ T_WLA<127> T_WLA<126> T_WLA<125> T_WLA<124> T_WLA<123> T_WLA<122> T_WLA<121> T_WLA<120> T_WLA<119> 
+ T_WLA<118> T_WLA<117> T_WLA<116> T_WLA<115> T_WLA<114> T_WLA<113> T_WLA<112> T_WLA<111> T_WLA<110> 
+ T_WLA<109> T_WLA<108> T_WLA<107> T_WLA<106> T_WLA<105> T_WLA<104> T_WLA<103> T_WLA<102> T_WLA<101> 
+ T_WLA<100> T_WLA<99> T_WLA<98> T_WLA<97> T_WLA<96> T_WLA<95> T_WLA<94> T_WLA<93> T_WLA<92> 
+ T_WLA<91> T_WLA<90> T_WLA<89> T_WLA<88> T_WLA<87> T_WLA<86> T_WLA<85> T_WLA<84> T_WLA<83> 
+ T_WLA<82> T_WLA<81> T_WLA<80> T_WLA<79> T_WLA<78> T_WLA<77> T_WLA<76> T_WLA<75> T_WLA<74> 
+ T_WLA<73> T_WLA<72> T_WLA<71> T_WLA<70> T_WLA<69> T_WLA<68> T_WLA<67> T_WLA<66> T_WLA<65> 
+ T_WLA<64> T_WLA<63> T_WLA<62> T_WLA<61> T_WLA<60> T_WLA<59> T_WLA<58> T_WLA<57> T_WLA<56> 
+ T_WLA<55> T_WLA<54> T_WLA<53> T_WLA<52> T_WLA<51> T_WLA<50> T_WLA<49> T_WLA<48> T_WLA<47> 
+ T_WLA<46> T_WLA<45> T_WLA<44> T_WLA<43> T_WLA<42> T_WLA<41> T_WLA<40> T_WLA<39> T_WLA<38> 
+ T_WLA<37> T_WLA<36> T_WLA<35> T_WLA<34> T_WLA<33> T_WLA<32> T_WLA<31> T_WLA<30> T_WLA<29> 
+ T_WLA<28> T_WLA<27> T_WLA<26> T_WLA<25> T_WLA<24> T_WLA<23> T_WLA<22> T_WLA<21> T_WLA<20> 
+ T_WLA<19> T_WLA<18> T_WLA<17> T_WLA<16> T_WLA<15> T_WLA<14> T_WLA<13> T_WLA<12> T_WLA<11> 
+ T_WLA<10> T_WLA<9> T_WLA<8> T_WLA<7> T_WLA<6> T_WLA<5> T_WLA<4> T_WLA<3> T_WLA<2> 
+ T_WLA<1> T_WLA<0> T_WLB<255> T_WLB<254> T_WLB<253> T_WLB<252> T_WLB<251> T_WLB<250> T_WLB<249> 
+ T_WLB<248> T_WLB<247> T_WLB<246> T_WLB<245> T_WLB<244> T_WLB<243> T_WLB<242> T_WLB<241> T_WLB<240> 
+ T_WLB<239> T_WLB<238> T_WLB<237> T_WLB<236> T_WLB<235> T_WLB<234> T_WLB<233> T_WLB<232> T_WLB<231> 
+ T_WLB<230> T_WLB<229> T_WLB<228> T_WLB<227> T_WLB<226> T_WLB<225> T_WLB<224> T_WLB<223> T_WLB<222> 
+ T_WLB<221> T_WLB<220> T_WLB<219> T_WLB<218> T_WLB<217> T_WLB<216> T_WLB<215> T_WLB<214> T_WLB<213> 
+ T_WLB<212> T_WLB<211> T_WLB<210> T_WLB<209> T_WLB<208> T_WLB<207> T_WLB<206> T_WLB<205> T_WLB<204> 
+ T_WLB<203> T_WLB<202> T_WLB<201> T_WLB<200> T_WLB<199> T_WLB<198> T_WLB<197> T_WLB<196> T_WLB<195> 
+ T_WLB<194> T_WLB<193> T_WLB<192> T_WLB<191> T_WLB<190> T_WLB<189> T_WLB<188> T_WLB<187> T_WLB<186> 
+ T_WLB<185> T_WLB<184> T_WLB<183> T_WLB<182> T_WLB<181> T_WLB<180> T_WLB<179> T_WLB<178> T_WLB<177> 
+ T_WLB<176> T_WLB<175> T_WLB<174> T_WLB<173> T_WLB<172> T_WLB<171> T_WLB<170> T_WLB<169> T_WLB<168> 
+ T_WLB<167> T_WLB<166> T_WLB<165> T_WLB<164> T_WLB<163> T_WLB<162> T_WLB<161> T_WLB<160> T_WLB<159> 
+ T_WLB<158> T_WLB<157> T_WLB<156> T_WLB<155> T_WLB<154> T_WLB<153> T_WLB<152> T_WLB<151> T_WLB<150> 
+ T_WLB<149> T_WLB<148> T_WLB<147> T_WLB<146> T_WLB<145> T_WLB<144> T_WLB<143> T_WLB<142> T_WLB<141> 
+ T_WLB<140> T_WLB<139> T_WLB<138> T_WLB<137> T_WLB<136> T_WLB<135> T_WLB<134> T_WLB<133> T_WLB<132> 
+ T_WLB<131> T_WLB<130> T_WLB<129> T_WLB<128> T_WLB<127> T_WLB<126> T_WLB<125> T_WLB<124> T_WLB<123> 
+ T_WLB<122> T_WLB<121> T_WLB<120> T_WLB<119> T_WLB<118> T_WLB<117> T_WLB<116> T_WLB<115> T_WLB<114> 
+ T_WLB<113> T_WLB<112> T_WLB<111> T_WLB<110> T_WLB<109> T_WLB<108> T_WLB<107> T_WLB<106> T_WLB<105> 
+ T_WLB<104> T_WLB<103> T_WLB<102> T_WLB<101> T_WLB<100> T_WLB<99> T_WLB<98> T_WLB<97> T_WLB<96> 
+ T_WLB<95> T_WLB<94> T_WLB<93> T_WLB<92> T_WLB<91> T_WLB<90> T_WLB<89> T_WLB<88> T_WLB<87> 
+ T_WLB<86> T_WLB<85> T_WLB<84> T_WLB<83> T_WLB<82> T_WLB<81> T_WLB<80> T_WLB<79> T_WLB<78> 
+ T_WLB<77> T_WLB<76> T_WLB<75> T_WLB<74> T_WLB<73> T_WLB<72> T_WLB<71> T_WLB<70> T_WLB<69> 
+ T_WLB<68> T_WLB<67> T_WLB<66> T_WLB<65> T_WLB<64> T_WLB<63> T_WLB<62> T_WLB<61> T_WLB<60> 
+ T_WLB<59> T_WLB<58> T_WLB<57> T_WLB<56> T_WLB<55> T_WLB<54> T_WLB<53> T_WLB<52> T_WLB<51> 
+ T_WLB<50> T_WLB<49> T_WLB<48> T_WLB<47> T_WLB<46> T_WLB<45> T_WLB<44> T_WLB<43> T_WLB<42> 
+ T_WLB<41> T_WLB<40> T_WLB<39> T_WLB<38> T_WLB<37> T_WLB<36> T_WLB<35> T_WLB<34> T_WLB<33> 
+ T_WLB<32> T_WLB<31> T_WLB<30> T_WLB<29> T_WLB<28> T_WLB<27> T_WLB<26> T_WLB<25> T_WLB<24> 
+ T_WLB<23> T_WLB<22> T_WLB<21> T_WLB<20> T_WLB<19> T_WLB<18> T_WLB<17> T_WLB<16> T_WLB<15> 
+ T_WLB<14> T_WLB<13> T_WLB<12> T_WLB<11> T_WLB<10> T_WLB<9> T_WLB<8> T_WLB<7> T_WLB<6> 
+ T_WLB<5> T_WLB<4> T_WLB<3> T_WLB<2> T_WLB<1> T_WLB<0> VDD VSS  / dpram16x4096_SingleCOL2X8_ROWX256
XCOL2<2>
+ RB_CA<3> RB_CA<2> RB_CA<1> RB_CA<0> RB_CB<3> RB_CB<2> RB_CB<1> RB_CB<0> RB_MA<3> 
+ RB_MA<2> RB_MA<1> RB_MA<0> RB_MB<3> RB_MB<2> RB_MB<1> RB_MB<0> RB_TM_PREB_N RB_TM_PREA_N 
+ B_WLA<255> B_WLA<254> B_WLA<253> B_WLA<252> B_WLA<251> B_WLA<250> B_WLA<249> B_WLA<248> B_WLA<247> 
+ B_WLA<246> B_WLA<245> B_WLA<244> B_WLA<243> B_WLA<242> B_WLA<241> B_WLA<240> B_WLA<239> B_WLA<238> 
+ B_WLA<237> B_WLA<236> B_WLA<235> B_WLA<234> B_WLA<233> B_WLA<232> B_WLA<231> B_WLA<230> B_WLA<229> 
+ B_WLA<228> B_WLA<227> B_WLA<226> B_WLA<225> B_WLA<224> B_WLA<223> B_WLA<222> B_WLA<221> B_WLA<220> 
+ B_WLA<219> B_WLA<218> B_WLA<217> B_WLA<216> B_WLA<215> B_WLA<214> B_WLA<213> B_WLA<212> B_WLA<211> 
+ B_WLA<210> B_WLA<209> B_WLA<208> B_WLA<207> B_WLA<206> B_WLA<205> B_WLA<204> B_WLA<203> B_WLA<202> 
+ B_WLA<201> B_WLA<200> B_WLA<199> B_WLA<198> B_WLA<197> B_WLA<196> B_WLA<195> B_WLA<194> B_WLA<193> 
+ B_WLA<192> B_WLA<191> B_WLA<190> B_WLA<189> B_WLA<188> B_WLA<187> B_WLA<186> B_WLA<185> B_WLA<184> 
+ B_WLA<183> B_WLA<182> B_WLA<181> B_WLA<180> B_WLA<179> B_WLA<178> B_WLA<177> B_WLA<176> B_WLA<175> 
+ B_WLA<174> B_WLA<173> B_WLA<172> B_WLA<171> B_WLA<170> B_WLA<169> B_WLA<168> B_WLA<167> B_WLA<166> 
+ B_WLA<165> B_WLA<164> B_WLA<163> B_WLA<162> B_WLA<161> B_WLA<160> B_WLA<159> B_WLA<158> B_WLA<157> 
+ B_WLA<156> B_WLA<155> B_WLA<154> B_WLA<153> B_WLA<152> B_WLA<151> B_WLA<150> B_WLA<149> B_WLA<148> 
+ B_WLA<147> B_WLA<146> B_WLA<145> B_WLA<144> B_WLA<143> B_WLA<142> B_WLA<141> B_WLA<140> B_WLA<139> 
+ B_WLA<138> B_WLA<137> B_WLA<136> B_WLA<135> B_WLA<134> B_WLA<133> B_WLA<132> B_WLA<131> B_WLA<130> 
+ B_WLA<129> B_WLA<128> B_WLA<127> B_WLA<126> B_WLA<125> B_WLA<124> B_WLA<123> B_WLA<122> B_WLA<121> 
+ B_WLA<120> B_WLA<119> B_WLA<118> B_WLA<117> B_WLA<116> B_WLA<115> B_WLA<114> B_WLA<113> B_WLA<112> 
+ B_WLA<111> B_WLA<110> B_WLA<109> B_WLA<108> B_WLA<107> B_WLA<106> B_WLA<105> B_WLA<104> B_WLA<103> 
+ B_WLA<102> B_WLA<101> B_WLA<100> B_WLA<99> B_WLA<98> B_WLA<97> B_WLA<96> B_WLA<95> B_WLA<94> 
+ B_WLA<93> B_WLA<92> B_WLA<91> B_WLA<90> B_WLA<89> B_WLA<88> B_WLA<87> B_WLA<86> B_WLA<85> 
+ B_WLA<84> B_WLA<83> B_WLA<82> B_WLA<81> B_WLA<80> B_WLA<79> B_WLA<78> B_WLA<77> B_WLA<76> 
+ B_WLA<75> B_WLA<74> B_WLA<73> B_WLA<72> B_WLA<71> B_WLA<70> B_WLA<69> B_WLA<68> B_WLA<67> 
+ B_WLA<66> B_WLA<65> B_WLA<64> B_WLA<63> B_WLA<62> B_WLA<61> B_WLA<60> B_WLA<59> B_WLA<58> 
+ B_WLA<57> B_WLA<56> B_WLA<55> B_WLA<54> B_WLA<53> B_WLA<52> B_WLA<51> B_WLA<50> B_WLA<49> 
+ B_WLA<48> B_WLA<47> B_WLA<46> B_WLA<45> B_WLA<44> B_WLA<43> B_WLA<42> B_WLA<41> B_WLA<40> 
+ B_WLA<39> B_WLA<38> B_WLA<37> B_WLA<36> B_WLA<35> B_WLA<34> B_WLA<33> B_WLA<32> B_WLA<31> 
+ B_WLA<30> B_WLA<29> B_WLA<28> B_WLA<27> B_WLA<26> B_WLA<25> B_WLA<24> B_WLA<23> B_WLA<22> 
+ B_WLA<21> B_WLA<20> B_WLA<19> B_WLA<18> B_WLA<17> B_WLA<16> B_WLA<15> B_WLA<14> B_WLA<13> 
+ B_WLA<12> B_WLA<11> B_WLA<10> B_WLA<9> B_WLA<8> B_WLA<7> B_WLA<6> B_WLA<5> B_WLA<4> 
+ B_WLA<3> B_WLA<2> B_WLA<1> B_WLA<0> B_WLB<255> B_WLB<254> B_WLB<253> B_WLB<252> B_WLB<251> 
+ B_WLB<250> B_WLB<249> B_WLB<248> B_WLB<247> B_WLB<246> B_WLB<245> B_WLB<244> B_WLB<243> B_WLB<242> 
+ B_WLB<241> B_WLB<240> B_WLB<239> B_WLB<238> B_WLB<237> B_WLB<236> B_WLB<235> B_WLB<234> B_WLB<233> 
+ B_WLB<232> B_WLB<231> B_WLB<230> B_WLB<229> B_WLB<228> B_WLB<227> B_WLB<226> B_WLB<225> B_WLB<224> 
+ B_WLB<223> B_WLB<222> B_WLB<221> B_WLB<220> B_WLB<219> B_WLB<218> B_WLB<217> B_WLB<216> B_WLB<215> 
+ B_WLB<214> B_WLB<213> B_WLB<212> B_WLB<211> B_WLB<210> B_WLB<209> B_WLB<208> B_WLB<207> B_WLB<206> 
+ B_WLB<205> B_WLB<204> B_WLB<203> B_WLB<202> B_WLB<201> B_WLB<200> B_WLB<199> B_WLB<198> B_WLB<197> 
+ B_WLB<196> B_WLB<195> B_WLB<194> B_WLB<193> B_WLB<192> B_WLB<191> B_WLB<190> B_WLB<189> B_WLB<188> 
+ B_WLB<187> B_WLB<186> B_WLB<185> B_WLB<184> B_WLB<183> B_WLB<182> B_WLB<181> B_WLB<180> B_WLB<179> 
+ B_WLB<178> B_WLB<177> B_WLB<176> B_WLB<175> B_WLB<174> B_WLB<173> B_WLB<172> B_WLB<171> B_WLB<170> 
+ B_WLB<169> B_WLB<168> B_WLB<167> B_WLB<166> B_WLB<165> B_WLB<164> B_WLB<163> B_WLB<162> B_WLB<161> 
+ B_WLB<160> B_WLB<159> B_WLB<158> B_WLB<157> B_WLB<156> B_WLB<155> B_WLB<154> B_WLB<153> B_WLB<152> 
+ B_WLB<151> B_WLB<150> B_WLB<149> B_WLB<148> B_WLB<147> B_WLB<146> B_WLB<145> B_WLB<144> B_WLB<143> 
+ B_WLB<142> B_WLB<141> B_WLB<140> B_WLB<139> B_WLB<138> B_WLB<137> B_WLB<136> B_WLB<135> B_WLB<134> 
+ B_WLB<133> B_WLB<132> B_WLB<131> B_WLB<130> B_WLB<129> B_WLB<128> B_WLB<127> B_WLB<126> B_WLB<125> 
+ B_WLB<124> B_WLB<123> B_WLB<122> B_WLB<121> B_WLB<120> B_WLB<119> B_WLB<118> B_WLB<117> B_WLB<116> 
+ B_WLB<115> B_WLB<114> B_WLB<113> B_WLB<112> B_WLB<111> B_WLB<110> B_WLB<109> B_WLB<108> B_WLB<107> 
+ B_WLB<106> B_WLB<105> B_WLB<104> B_WLB<103> B_WLB<102> B_WLB<101> B_WLB<100> B_WLB<99> B_WLB<98> 
+ B_WLB<97> B_WLB<96> B_WLB<95> B_WLB<94> B_WLB<93> B_WLB<92> B_WLB<91> B_WLB<90> B_WLB<89> 
+ B_WLB<88> B_WLB<87> B_WLB<86> B_WLB<85> B_WLB<84> B_WLB<83> B_WLB<82> B_WLB<81> B_WLB<80> 
+ B_WLB<79> B_WLB<78> B_WLB<77> B_WLB<76> B_WLB<75> B_WLB<74> B_WLB<73> B_WLB<72> B_WLB<71> 
+ B_WLB<70> B_WLB<69> B_WLB<68> B_WLB<67> B_WLB<66> B_WLB<65> B_WLB<64> B_WLB<63> B_WLB<62> 
+ B_WLB<61> B_WLB<60> B_WLB<59> B_WLB<58> B_WLB<57> B_WLB<56> B_WLB<55> B_WLB<54> B_WLB<53> 
+ B_WLB<52> B_WLB<51> B_WLB<50> B_WLB<49> B_WLB<48> B_WLB<47> B_WLB<46> B_WLB<45> B_WLB<44> 
+ B_WLB<43> B_WLB<42> B_WLB<41> B_WLB<40> B_WLB<39> B_WLB<38> B_WLB<37> B_WLB<36> B_WLB<35> 
+ B_WLB<34> B_WLB<33> B_WLB<32> B_WLB<31> B_WLB<30> B_WLB<29> B_WLB<28> B_WLB<27> B_WLB<26> 
+ B_WLB<25> B_WLB<24> B_WLB<23> B_WLB<22> B_WLB<21> B_WLB<20> B_WLB<19> B_WLB<18> B_WLB<17> 
+ B_WLB<16> B_WLB<15> B_WLB<14> B_WLB<13> B_WLB<12> B_WLB<11> B_WLB<10> B_WLB<9> B_WLB<8> 
+ B_WLB<7> B_WLB<6> B_WLB<5> B_WLB<4> B_WLB<3> B_WLB<2> B_WLB<1> B_WLB<0> BWENA<5> 
+ BWENA<4> BWENB<5> BWENB<4> R_CLK_DQA R_CLK_DQA_N R_CLK_DQB R_CLK_DQB_N DA<5> DA<4> 
+ DB<5> DB<4> DDQA<2> DDQA_N<2> DDQB<2> DDQB_N<2> R_LWEA R_LWEB QA<5> 
+ QA<4> QB<5> QB<4> R_SA_PREA_N R_SA_PREB_N R_SAEA_N R_SAEB_N RT_CA<3> RT_CA<2> 
+ RT_CA<1> RT_CA<0> RT_CB<3> RT_CB<2> RT_CB<1> RT_CB<0> RT_MA<3> RT_MA<2> RT_MA<1> 
+ RT_MA<0> RT_MB<3> RT_MB<2> RT_MB<1> RT_MB<0> R_TM_PREA_N R_TM_PREB_N T_WLA<255> T_WLA<254> 
+ T_WLA<253> T_WLA<252> T_WLA<251> T_WLA<250> T_WLA<249> T_WLA<248> T_WLA<247> T_WLA<246> T_WLA<245> 
+ T_WLA<244> T_WLA<243> T_WLA<242> T_WLA<241> T_WLA<240> T_WLA<239> T_WLA<238> T_WLA<237> T_WLA<236> 
+ T_WLA<235> T_WLA<234> T_WLA<233> T_WLA<232> T_WLA<231> T_WLA<230> T_WLA<229> T_WLA<228> T_WLA<227> 
+ T_WLA<226> T_WLA<225> T_WLA<224> T_WLA<223> T_WLA<222> T_WLA<221> T_WLA<220> T_WLA<219> T_WLA<218> 
+ T_WLA<217> T_WLA<216> T_WLA<215> T_WLA<214> T_WLA<213> T_WLA<212> T_WLA<211> T_WLA<210> T_WLA<209> 
+ T_WLA<208> T_WLA<207> T_WLA<206> T_WLA<205> T_WLA<204> T_WLA<203> T_WLA<202> T_WLA<201> T_WLA<200> 
+ T_WLA<199> T_WLA<198> T_WLA<197> T_WLA<196> T_WLA<195> T_WLA<194> T_WLA<193> T_WLA<192> T_WLA<191> 
+ T_WLA<190> T_WLA<189> T_WLA<188> T_WLA<187> T_WLA<186> T_WLA<185> T_WLA<184> T_WLA<183> T_WLA<182> 
+ T_WLA<181> T_WLA<180> T_WLA<179> T_WLA<178> T_WLA<177> T_WLA<176> T_WLA<175> T_WLA<174> T_WLA<173> 
+ T_WLA<172> T_WLA<171> T_WLA<170> T_WLA<169> T_WLA<168> T_WLA<167> T_WLA<166> T_WLA<165> T_WLA<164> 
+ T_WLA<163> T_WLA<162> T_WLA<161> T_WLA<160> T_WLA<159> T_WLA<158> T_WLA<157> T_WLA<156> T_WLA<155> 
+ T_WLA<154> T_WLA<153> T_WLA<152> T_WLA<151> T_WLA<150> T_WLA<149> T_WLA<148> T_WLA<147> T_WLA<146> 
+ T_WLA<145> T_WLA<144> T_WLA<143> T_WLA<142> T_WLA<141> T_WLA<140> T_WLA<139> T_WLA<138> T_WLA<137> 
+ T_WLA<136> T_WLA<135> T_WLA<134> T_WLA<133> T_WLA<132> T_WLA<131> T_WLA<130> T_WLA<129> T_WLA<128> 
+ T_WLA<127> T_WLA<126> T_WLA<125> T_WLA<124> T_WLA<123> T_WLA<122> T_WLA<121> T_WLA<120> T_WLA<119> 
+ T_WLA<118> T_WLA<117> T_WLA<116> T_WLA<115> T_WLA<114> T_WLA<113> T_WLA<112> T_WLA<111> T_WLA<110> 
+ T_WLA<109> T_WLA<108> T_WLA<107> T_WLA<106> T_WLA<105> T_WLA<104> T_WLA<103> T_WLA<102> T_WLA<101> 
+ T_WLA<100> T_WLA<99> T_WLA<98> T_WLA<97> T_WLA<96> T_WLA<95> T_WLA<94> T_WLA<93> T_WLA<92> 
+ T_WLA<91> T_WLA<90> T_WLA<89> T_WLA<88> T_WLA<87> T_WLA<86> T_WLA<85> T_WLA<84> T_WLA<83> 
+ T_WLA<82> T_WLA<81> T_WLA<80> T_WLA<79> T_WLA<78> T_WLA<77> T_WLA<76> T_WLA<75> T_WLA<74> 
+ T_WLA<73> T_WLA<72> T_WLA<71> T_WLA<70> T_WLA<69> T_WLA<68> T_WLA<67> T_WLA<66> T_WLA<65> 
+ T_WLA<64> T_WLA<63> T_WLA<62> T_WLA<61> T_WLA<60> T_WLA<59> T_WLA<58> T_WLA<57> T_WLA<56> 
+ T_WLA<55> T_WLA<54> T_WLA<53> T_WLA<52> T_WLA<51> T_WLA<50> T_WLA<49> T_WLA<48> T_WLA<47> 
+ T_WLA<46> T_WLA<45> T_WLA<44> T_WLA<43> T_WLA<42> T_WLA<41> T_WLA<40> T_WLA<39> T_WLA<38> 
+ T_WLA<37> T_WLA<36> T_WLA<35> T_WLA<34> T_WLA<33> T_WLA<32> T_WLA<31> T_WLA<30> T_WLA<29> 
+ T_WLA<28> T_WLA<27> T_WLA<26> T_WLA<25> T_WLA<24> T_WLA<23> T_WLA<22> T_WLA<21> T_WLA<20> 
+ T_WLA<19> T_WLA<18> T_WLA<17> T_WLA<16> T_WLA<15> T_WLA<14> T_WLA<13> T_WLA<12> T_WLA<11> 
+ T_WLA<10> T_WLA<9> T_WLA<8> T_WLA<7> T_WLA<6> T_WLA<5> T_WLA<4> T_WLA<3> T_WLA<2> 
+ T_WLA<1> T_WLA<0> T_WLB<255> T_WLB<254> T_WLB<253> T_WLB<252> T_WLB<251> T_WLB<250> T_WLB<249> 
+ T_WLB<248> T_WLB<247> T_WLB<246> T_WLB<245> T_WLB<244> T_WLB<243> T_WLB<242> T_WLB<241> T_WLB<240> 
+ T_WLB<239> T_WLB<238> T_WLB<237> T_WLB<236> T_WLB<235> T_WLB<234> T_WLB<233> T_WLB<232> T_WLB<231> 
+ T_WLB<230> T_WLB<229> T_WLB<228> T_WLB<227> T_WLB<226> T_WLB<225> T_WLB<224> T_WLB<223> T_WLB<222> 
+ T_WLB<221> T_WLB<220> T_WLB<219> T_WLB<218> T_WLB<217> T_WLB<216> T_WLB<215> T_WLB<214> T_WLB<213> 
+ T_WLB<212> T_WLB<211> T_WLB<210> T_WLB<209> T_WLB<208> T_WLB<207> T_WLB<206> T_WLB<205> T_WLB<204> 
+ T_WLB<203> T_WLB<202> T_WLB<201> T_WLB<200> T_WLB<199> T_WLB<198> T_WLB<197> T_WLB<196> T_WLB<195> 
+ T_WLB<194> T_WLB<193> T_WLB<192> T_WLB<191> T_WLB<190> T_WLB<189> T_WLB<188> T_WLB<187> T_WLB<186> 
+ T_WLB<185> T_WLB<184> T_WLB<183> T_WLB<182> T_WLB<181> T_WLB<180> T_WLB<179> T_WLB<178> T_WLB<177> 
+ T_WLB<176> T_WLB<175> T_WLB<174> T_WLB<173> T_WLB<172> T_WLB<171> T_WLB<170> T_WLB<169> T_WLB<168> 
+ T_WLB<167> T_WLB<166> T_WLB<165> T_WLB<164> T_WLB<163> T_WLB<162> T_WLB<161> T_WLB<160> T_WLB<159> 
+ T_WLB<158> T_WLB<157> T_WLB<156> T_WLB<155> T_WLB<154> T_WLB<153> T_WLB<152> T_WLB<151> T_WLB<150> 
+ T_WLB<149> T_WLB<148> T_WLB<147> T_WLB<146> T_WLB<145> T_WLB<144> T_WLB<143> T_WLB<142> T_WLB<141> 
+ T_WLB<140> T_WLB<139> T_WLB<138> T_WLB<137> T_WLB<136> T_WLB<135> T_WLB<134> T_WLB<133> T_WLB<132> 
+ T_WLB<131> T_WLB<130> T_WLB<129> T_WLB<128> T_WLB<127> T_WLB<126> T_WLB<125> T_WLB<124> T_WLB<123> 
+ T_WLB<122> T_WLB<121> T_WLB<120> T_WLB<119> T_WLB<118> T_WLB<117> T_WLB<116> T_WLB<115> T_WLB<114> 
+ T_WLB<113> T_WLB<112> T_WLB<111> T_WLB<110> T_WLB<109> T_WLB<108> T_WLB<107> T_WLB<106> T_WLB<105> 
+ T_WLB<104> T_WLB<103> T_WLB<102> T_WLB<101> T_WLB<100> T_WLB<99> T_WLB<98> T_WLB<97> T_WLB<96> 
+ T_WLB<95> T_WLB<94> T_WLB<93> T_WLB<92> T_WLB<91> T_WLB<90> T_WLB<89> T_WLB<88> T_WLB<87> 
+ T_WLB<86> T_WLB<85> T_WLB<84> T_WLB<83> T_WLB<82> T_WLB<81> T_WLB<80> T_WLB<79> T_WLB<78> 
+ T_WLB<77> T_WLB<76> T_WLB<75> T_WLB<74> T_WLB<73> T_WLB<72> T_WLB<71> T_WLB<70> T_WLB<69> 
+ T_WLB<68> T_WLB<67> T_WLB<66> T_WLB<65> T_WLB<64> T_WLB<63> T_WLB<62> T_WLB<61> T_WLB<60> 
+ T_WLB<59> T_WLB<58> T_WLB<57> T_WLB<56> T_WLB<55> T_WLB<54> T_WLB<53> T_WLB<52> T_WLB<51> 
+ T_WLB<50> T_WLB<49> T_WLB<48> T_WLB<47> T_WLB<46> T_WLB<45> T_WLB<44> T_WLB<43> T_WLB<42> 
+ T_WLB<41> T_WLB<40> T_WLB<39> T_WLB<38> T_WLB<37> T_WLB<36> T_WLB<35> T_WLB<34> T_WLB<33> 
+ T_WLB<32> T_WLB<31> T_WLB<30> T_WLB<29> T_WLB<28> T_WLB<27> T_WLB<26> T_WLB<25> T_WLB<24> 
+ T_WLB<23> T_WLB<22> T_WLB<21> T_WLB<20> T_WLB<19> T_WLB<18> T_WLB<17> T_WLB<16> T_WLB<15> 
+ T_WLB<14> T_WLB<13> T_WLB<12> T_WLB<11> T_WLB<10> T_WLB<9> T_WLB<8> T_WLB<7> T_WLB<6> 
+ T_WLB<5> T_WLB<4> T_WLB<3> T_WLB<2> T_WLB<1> T_WLB<0> VDD VSS  / dpram16x4096_SingleCOL2X8_ROWX256
XCOL2<1>
+ RB_CA<3> RB_CA<2> RB_CA<1> RB_CA<0> RB_CB<3> RB_CB<2> RB_CB<1> RB_CB<0> RB_MA<3> 
+ RB_MA<2> RB_MA<1> RB_MA<0> RB_MB<3> RB_MB<2> RB_MB<1> RB_MB<0> RB_TM_PREB_N RB_TM_PREA_N 
+ B_WLA<255> B_WLA<254> B_WLA<253> B_WLA<252> B_WLA<251> B_WLA<250> B_WLA<249> B_WLA<248> B_WLA<247> 
+ B_WLA<246> B_WLA<245> B_WLA<244> B_WLA<243> B_WLA<242> B_WLA<241> B_WLA<240> B_WLA<239> B_WLA<238> 
+ B_WLA<237> B_WLA<236> B_WLA<235> B_WLA<234> B_WLA<233> B_WLA<232> B_WLA<231> B_WLA<230> B_WLA<229> 
+ B_WLA<228> B_WLA<227> B_WLA<226> B_WLA<225> B_WLA<224> B_WLA<223> B_WLA<222> B_WLA<221> B_WLA<220> 
+ B_WLA<219> B_WLA<218> B_WLA<217> B_WLA<216> B_WLA<215> B_WLA<214> B_WLA<213> B_WLA<212> B_WLA<211> 
+ B_WLA<210> B_WLA<209> B_WLA<208> B_WLA<207> B_WLA<206> B_WLA<205> B_WLA<204> B_WLA<203> B_WLA<202> 
+ B_WLA<201> B_WLA<200> B_WLA<199> B_WLA<198> B_WLA<197> B_WLA<196> B_WLA<195> B_WLA<194> B_WLA<193> 
+ B_WLA<192> B_WLA<191> B_WLA<190> B_WLA<189> B_WLA<188> B_WLA<187> B_WLA<186> B_WLA<185> B_WLA<184> 
+ B_WLA<183> B_WLA<182> B_WLA<181> B_WLA<180> B_WLA<179> B_WLA<178> B_WLA<177> B_WLA<176> B_WLA<175> 
+ B_WLA<174> B_WLA<173> B_WLA<172> B_WLA<171> B_WLA<170> B_WLA<169> B_WLA<168> B_WLA<167> B_WLA<166> 
+ B_WLA<165> B_WLA<164> B_WLA<163> B_WLA<162> B_WLA<161> B_WLA<160> B_WLA<159> B_WLA<158> B_WLA<157> 
+ B_WLA<156> B_WLA<155> B_WLA<154> B_WLA<153> B_WLA<152> B_WLA<151> B_WLA<150> B_WLA<149> B_WLA<148> 
+ B_WLA<147> B_WLA<146> B_WLA<145> B_WLA<144> B_WLA<143> B_WLA<142> B_WLA<141> B_WLA<140> B_WLA<139> 
+ B_WLA<138> B_WLA<137> B_WLA<136> B_WLA<135> B_WLA<134> B_WLA<133> B_WLA<132> B_WLA<131> B_WLA<130> 
+ B_WLA<129> B_WLA<128> B_WLA<127> B_WLA<126> B_WLA<125> B_WLA<124> B_WLA<123> B_WLA<122> B_WLA<121> 
+ B_WLA<120> B_WLA<119> B_WLA<118> B_WLA<117> B_WLA<116> B_WLA<115> B_WLA<114> B_WLA<113> B_WLA<112> 
+ B_WLA<111> B_WLA<110> B_WLA<109> B_WLA<108> B_WLA<107> B_WLA<106> B_WLA<105> B_WLA<104> B_WLA<103> 
+ B_WLA<102> B_WLA<101> B_WLA<100> B_WLA<99> B_WLA<98> B_WLA<97> B_WLA<96> B_WLA<95> B_WLA<94> 
+ B_WLA<93> B_WLA<92> B_WLA<91> B_WLA<90> B_WLA<89> B_WLA<88> B_WLA<87> B_WLA<86> B_WLA<85> 
+ B_WLA<84> B_WLA<83> B_WLA<82> B_WLA<81> B_WLA<80> B_WLA<79> B_WLA<78> B_WLA<77> B_WLA<76> 
+ B_WLA<75> B_WLA<74> B_WLA<73> B_WLA<72> B_WLA<71> B_WLA<70> B_WLA<69> B_WLA<68> B_WLA<67> 
+ B_WLA<66> B_WLA<65> B_WLA<64> B_WLA<63> B_WLA<62> B_WLA<61> B_WLA<60> B_WLA<59> B_WLA<58> 
+ B_WLA<57> B_WLA<56> B_WLA<55> B_WLA<54> B_WLA<53> B_WLA<52> B_WLA<51> B_WLA<50> B_WLA<49> 
+ B_WLA<48> B_WLA<47> B_WLA<46> B_WLA<45> B_WLA<44> B_WLA<43> B_WLA<42> B_WLA<41> B_WLA<40> 
+ B_WLA<39> B_WLA<38> B_WLA<37> B_WLA<36> B_WLA<35> B_WLA<34> B_WLA<33> B_WLA<32> B_WLA<31> 
+ B_WLA<30> B_WLA<29> B_WLA<28> B_WLA<27> B_WLA<26> B_WLA<25> B_WLA<24> B_WLA<23> B_WLA<22> 
+ B_WLA<21> B_WLA<20> B_WLA<19> B_WLA<18> B_WLA<17> B_WLA<16> B_WLA<15> B_WLA<14> B_WLA<13> 
+ B_WLA<12> B_WLA<11> B_WLA<10> B_WLA<9> B_WLA<8> B_WLA<7> B_WLA<6> B_WLA<5> B_WLA<4> 
+ B_WLA<3> B_WLA<2> B_WLA<1> B_WLA<0> B_WLB<255> B_WLB<254> B_WLB<253> B_WLB<252> B_WLB<251> 
+ B_WLB<250> B_WLB<249> B_WLB<248> B_WLB<247> B_WLB<246> B_WLB<245> B_WLB<244> B_WLB<243> B_WLB<242> 
+ B_WLB<241> B_WLB<240> B_WLB<239> B_WLB<238> B_WLB<237> B_WLB<236> B_WLB<235> B_WLB<234> B_WLB<233> 
+ B_WLB<232> B_WLB<231> B_WLB<230> B_WLB<229> B_WLB<228> B_WLB<227> B_WLB<226> B_WLB<225> B_WLB<224> 
+ B_WLB<223> B_WLB<222> B_WLB<221> B_WLB<220> B_WLB<219> B_WLB<218> B_WLB<217> B_WLB<216> B_WLB<215> 
+ B_WLB<214> B_WLB<213> B_WLB<212> B_WLB<211> B_WLB<210> B_WLB<209> B_WLB<208> B_WLB<207> B_WLB<206> 
+ B_WLB<205> B_WLB<204> B_WLB<203> B_WLB<202> B_WLB<201> B_WLB<200> B_WLB<199> B_WLB<198> B_WLB<197> 
+ B_WLB<196> B_WLB<195> B_WLB<194> B_WLB<193> B_WLB<192> B_WLB<191> B_WLB<190> B_WLB<189> B_WLB<188> 
+ B_WLB<187> B_WLB<186> B_WLB<185> B_WLB<184> B_WLB<183> B_WLB<182> B_WLB<181> B_WLB<180> B_WLB<179> 
+ B_WLB<178> B_WLB<177> B_WLB<176> B_WLB<175> B_WLB<174> B_WLB<173> B_WLB<172> B_WLB<171> B_WLB<170> 
+ B_WLB<169> B_WLB<168> B_WLB<167> B_WLB<166> B_WLB<165> B_WLB<164> B_WLB<163> B_WLB<162> B_WLB<161> 
+ B_WLB<160> B_WLB<159> B_WLB<158> B_WLB<157> B_WLB<156> B_WLB<155> B_WLB<154> B_WLB<153> B_WLB<152> 
+ B_WLB<151> B_WLB<150> B_WLB<149> B_WLB<148> B_WLB<147> B_WLB<146> B_WLB<145> B_WLB<144> B_WLB<143> 
+ B_WLB<142> B_WLB<141> B_WLB<140> B_WLB<139> B_WLB<138> B_WLB<137> B_WLB<136> B_WLB<135> B_WLB<134> 
+ B_WLB<133> B_WLB<132> B_WLB<131> B_WLB<130> B_WLB<129> B_WLB<128> B_WLB<127> B_WLB<126> B_WLB<125> 
+ B_WLB<124> B_WLB<123> B_WLB<122> B_WLB<121> B_WLB<120> B_WLB<119> B_WLB<118> B_WLB<117> B_WLB<116> 
+ B_WLB<115> B_WLB<114> B_WLB<113> B_WLB<112> B_WLB<111> B_WLB<110> B_WLB<109> B_WLB<108> B_WLB<107> 
+ B_WLB<106> B_WLB<105> B_WLB<104> B_WLB<103> B_WLB<102> B_WLB<101> B_WLB<100> B_WLB<99> B_WLB<98> 
+ B_WLB<97> B_WLB<96> B_WLB<95> B_WLB<94> B_WLB<93> B_WLB<92> B_WLB<91> B_WLB<90> B_WLB<89> 
+ B_WLB<88> B_WLB<87> B_WLB<86> B_WLB<85> B_WLB<84> B_WLB<83> B_WLB<82> B_WLB<81> B_WLB<80> 
+ B_WLB<79> B_WLB<78> B_WLB<77> B_WLB<76> B_WLB<75> B_WLB<74> B_WLB<73> B_WLB<72> B_WLB<71> 
+ B_WLB<70> B_WLB<69> B_WLB<68> B_WLB<67> B_WLB<66> B_WLB<65> B_WLB<64> B_WLB<63> B_WLB<62> 
+ B_WLB<61> B_WLB<60> B_WLB<59> B_WLB<58> B_WLB<57> B_WLB<56> B_WLB<55> B_WLB<54> B_WLB<53> 
+ B_WLB<52> B_WLB<51> B_WLB<50> B_WLB<49> B_WLB<48> B_WLB<47> B_WLB<46> B_WLB<45> B_WLB<44> 
+ B_WLB<43> B_WLB<42> B_WLB<41> B_WLB<40> B_WLB<39> B_WLB<38> B_WLB<37> B_WLB<36> B_WLB<35> 
+ B_WLB<34> B_WLB<33> B_WLB<32> B_WLB<31> B_WLB<30> B_WLB<29> B_WLB<28> B_WLB<27> B_WLB<26> 
+ B_WLB<25> B_WLB<24> B_WLB<23> B_WLB<22> B_WLB<21> B_WLB<20> B_WLB<19> B_WLB<18> B_WLB<17> 
+ B_WLB<16> B_WLB<15> B_WLB<14> B_WLB<13> B_WLB<12> B_WLB<11> B_WLB<10> B_WLB<9> B_WLB<8> 
+ B_WLB<7> B_WLB<6> B_WLB<5> B_WLB<4> B_WLB<3> B_WLB<2> B_WLB<1> B_WLB<0> BWENA<3> 
+ BWENA<2> BWENB<3> BWENB<2> R_CLK_DQA R_CLK_DQA_N R_CLK_DQB R_CLK_DQB_N DA<3> DA<2> 
+ DB<3> DB<2> DDQA<1> DDQA_N<1> DDQB<1> DDQB_N<1> R_LWEA R_LWEB QA<3> 
+ QA<2> QB<3> QB<2> R_SA_PREA_N R_SA_PREB_N R_SAEA_N R_SAEB_N RT_CA<3> RT_CA<2> 
+ RT_CA<1> RT_CA<0> RT_CB<3> RT_CB<2> RT_CB<1> RT_CB<0> RT_MA<3> RT_MA<2> RT_MA<1> 
+ RT_MA<0> RT_MB<3> RT_MB<2> RT_MB<1> RT_MB<0> R_TM_PREA_N R_TM_PREB_N T_WLA<255> T_WLA<254> 
+ T_WLA<253> T_WLA<252> T_WLA<251> T_WLA<250> T_WLA<249> T_WLA<248> T_WLA<247> T_WLA<246> T_WLA<245> 
+ T_WLA<244> T_WLA<243> T_WLA<242> T_WLA<241> T_WLA<240> T_WLA<239> T_WLA<238> T_WLA<237> T_WLA<236> 
+ T_WLA<235> T_WLA<234> T_WLA<233> T_WLA<232> T_WLA<231> T_WLA<230> T_WLA<229> T_WLA<228> T_WLA<227> 
+ T_WLA<226> T_WLA<225> T_WLA<224> T_WLA<223> T_WLA<222> T_WLA<221> T_WLA<220> T_WLA<219> T_WLA<218> 
+ T_WLA<217> T_WLA<216> T_WLA<215> T_WLA<214> T_WLA<213> T_WLA<212> T_WLA<211> T_WLA<210> T_WLA<209> 
+ T_WLA<208> T_WLA<207> T_WLA<206> T_WLA<205> T_WLA<204> T_WLA<203> T_WLA<202> T_WLA<201> T_WLA<200> 
+ T_WLA<199> T_WLA<198> T_WLA<197> T_WLA<196> T_WLA<195> T_WLA<194> T_WLA<193> T_WLA<192> T_WLA<191> 
+ T_WLA<190> T_WLA<189> T_WLA<188> T_WLA<187> T_WLA<186> T_WLA<185> T_WLA<184> T_WLA<183> T_WLA<182> 
+ T_WLA<181> T_WLA<180> T_WLA<179> T_WLA<178> T_WLA<177> T_WLA<176> T_WLA<175> T_WLA<174> T_WLA<173> 
+ T_WLA<172> T_WLA<171> T_WLA<170> T_WLA<169> T_WLA<168> T_WLA<167> T_WLA<166> T_WLA<165> T_WLA<164> 
+ T_WLA<163> T_WLA<162> T_WLA<161> T_WLA<160> T_WLA<159> T_WLA<158> T_WLA<157> T_WLA<156> T_WLA<155> 
+ T_WLA<154> T_WLA<153> T_WLA<152> T_WLA<151> T_WLA<150> T_WLA<149> T_WLA<148> T_WLA<147> T_WLA<146> 
+ T_WLA<145> T_WLA<144> T_WLA<143> T_WLA<142> T_WLA<141> T_WLA<140> T_WLA<139> T_WLA<138> T_WLA<137> 
+ T_WLA<136> T_WLA<135> T_WLA<134> T_WLA<133> T_WLA<132> T_WLA<131> T_WLA<130> T_WLA<129> T_WLA<128> 
+ T_WLA<127> T_WLA<126> T_WLA<125> T_WLA<124> T_WLA<123> T_WLA<122> T_WLA<121> T_WLA<120> T_WLA<119> 
+ T_WLA<118> T_WLA<117> T_WLA<116> T_WLA<115> T_WLA<114> T_WLA<113> T_WLA<112> T_WLA<111> T_WLA<110> 
+ T_WLA<109> T_WLA<108> T_WLA<107> T_WLA<106> T_WLA<105> T_WLA<104> T_WLA<103> T_WLA<102> T_WLA<101> 
+ T_WLA<100> T_WLA<99> T_WLA<98> T_WLA<97> T_WLA<96> T_WLA<95> T_WLA<94> T_WLA<93> T_WLA<92> 
+ T_WLA<91> T_WLA<90> T_WLA<89> T_WLA<88> T_WLA<87> T_WLA<86> T_WLA<85> T_WLA<84> T_WLA<83> 
+ T_WLA<82> T_WLA<81> T_WLA<80> T_WLA<79> T_WLA<78> T_WLA<77> T_WLA<76> T_WLA<75> T_WLA<74> 
+ T_WLA<73> T_WLA<72> T_WLA<71> T_WLA<70> T_WLA<69> T_WLA<68> T_WLA<67> T_WLA<66> T_WLA<65> 
+ T_WLA<64> T_WLA<63> T_WLA<62> T_WLA<61> T_WLA<60> T_WLA<59> T_WLA<58> T_WLA<57> T_WLA<56> 
+ T_WLA<55> T_WLA<54> T_WLA<53> T_WLA<52> T_WLA<51> T_WLA<50> T_WLA<49> T_WLA<48> T_WLA<47> 
+ T_WLA<46> T_WLA<45> T_WLA<44> T_WLA<43> T_WLA<42> T_WLA<41> T_WLA<40> T_WLA<39> T_WLA<38> 
+ T_WLA<37> T_WLA<36> T_WLA<35> T_WLA<34> T_WLA<33> T_WLA<32> T_WLA<31> T_WLA<30> T_WLA<29> 
+ T_WLA<28> T_WLA<27> T_WLA<26> T_WLA<25> T_WLA<24> T_WLA<23> T_WLA<22> T_WLA<21> T_WLA<20> 
+ T_WLA<19> T_WLA<18> T_WLA<17> T_WLA<16> T_WLA<15> T_WLA<14> T_WLA<13> T_WLA<12> T_WLA<11> 
+ T_WLA<10> T_WLA<9> T_WLA<8> T_WLA<7> T_WLA<6> T_WLA<5> T_WLA<4> T_WLA<3> T_WLA<2> 
+ T_WLA<1> T_WLA<0> T_WLB<255> T_WLB<254> T_WLB<253> T_WLB<252> T_WLB<251> T_WLB<250> T_WLB<249> 
+ T_WLB<248> T_WLB<247> T_WLB<246> T_WLB<245> T_WLB<244> T_WLB<243> T_WLB<242> T_WLB<241> T_WLB<240> 
+ T_WLB<239> T_WLB<238> T_WLB<237> T_WLB<236> T_WLB<235> T_WLB<234> T_WLB<233> T_WLB<232> T_WLB<231> 
+ T_WLB<230> T_WLB<229> T_WLB<228> T_WLB<227> T_WLB<226> T_WLB<225> T_WLB<224> T_WLB<223> T_WLB<222> 
+ T_WLB<221> T_WLB<220> T_WLB<219> T_WLB<218> T_WLB<217> T_WLB<216> T_WLB<215> T_WLB<214> T_WLB<213> 
+ T_WLB<212> T_WLB<211> T_WLB<210> T_WLB<209> T_WLB<208> T_WLB<207> T_WLB<206> T_WLB<205> T_WLB<204> 
+ T_WLB<203> T_WLB<202> T_WLB<201> T_WLB<200> T_WLB<199> T_WLB<198> T_WLB<197> T_WLB<196> T_WLB<195> 
+ T_WLB<194> T_WLB<193> T_WLB<192> T_WLB<191> T_WLB<190> T_WLB<189> T_WLB<188> T_WLB<187> T_WLB<186> 
+ T_WLB<185> T_WLB<184> T_WLB<183> T_WLB<182> T_WLB<181> T_WLB<180> T_WLB<179> T_WLB<178> T_WLB<177> 
+ T_WLB<176> T_WLB<175> T_WLB<174> T_WLB<173> T_WLB<172> T_WLB<171> T_WLB<170> T_WLB<169> T_WLB<168> 
+ T_WLB<167> T_WLB<166> T_WLB<165> T_WLB<164> T_WLB<163> T_WLB<162> T_WLB<161> T_WLB<160> T_WLB<159> 
+ T_WLB<158> T_WLB<157> T_WLB<156> T_WLB<155> T_WLB<154> T_WLB<153> T_WLB<152> T_WLB<151> T_WLB<150> 
+ T_WLB<149> T_WLB<148> T_WLB<147> T_WLB<146> T_WLB<145> T_WLB<144> T_WLB<143> T_WLB<142> T_WLB<141> 
+ T_WLB<140> T_WLB<139> T_WLB<138> T_WLB<137> T_WLB<136> T_WLB<135> T_WLB<134> T_WLB<133> T_WLB<132> 
+ T_WLB<131> T_WLB<130> T_WLB<129> T_WLB<128> T_WLB<127> T_WLB<126> T_WLB<125> T_WLB<124> T_WLB<123> 
+ T_WLB<122> T_WLB<121> T_WLB<120> T_WLB<119> T_WLB<118> T_WLB<117> T_WLB<116> T_WLB<115> T_WLB<114> 
+ T_WLB<113> T_WLB<112> T_WLB<111> T_WLB<110> T_WLB<109> T_WLB<108> T_WLB<107> T_WLB<106> T_WLB<105> 
+ T_WLB<104> T_WLB<103> T_WLB<102> T_WLB<101> T_WLB<100> T_WLB<99> T_WLB<98> T_WLB<97> T_WLB<96> 
+ T_WLB<95> T_WLB<94> T_WLB<93> T_WLB<92> T_WLB<91> T_WLB<90> T_WLB<89> T_WLB<88> T_WLB<87> 
+ T_WLB<86> T_WLB<85> T_WLB<84> T_WLB<83> T_WLB<82> T_WLB<81> T_WLB<80> T_WLB<79> T_WLB<78> 
+ T_WLB<77> T_WLB<76> T_WLB<75> T_WLB<74> T_WLB<73> T_WLB<72> T_WLB<71> T_WLB<70> T_WLB<69> 
+ T_WLB<68> T_WLB<67> T_WLB<66> T_WLB<65> T_WLB<64> T_WLB<63> T_WLB<62> T_WLB<61> T_WLB<60> 
+ T_WLB<59> T_WLB<58> T_WLB<57> T_WLB<56> T_WLB<55> T_WLB<54> T_WLB<53> T_WLB<52> T_WLB<51> 
+ T_WLB<50> T_WLB<49> T_WLB<48> T_WLB<47> T_WLB<46> T_WLB<45> T_WLB<44> T_WLB<43> T_WLB<42> 
+ T_WLB<41> T_WLB<40> T_WLB<39> T_WLB<38> T_WLB<37> T_WLB<36> T_WLB<35> T_WLB<34> T_WLB<33> 
+ T_WLB<32> T_WLB<31> T_WLB<30> T_WLB<29> T_WLB<28> T_WLB<27> T_WLB<26> T_WLB<25> T_WLB<24> 
+ T_WLB<23> T_WLB<22> T_WLB<21> T_WLB<20> T_WLB<19> T_WLB<18> T_WLB<17> T_WLB<16> T_WLB<15> 
+ T_WLB<14> T_WLB<13> T_WLB<12> T_WLB<11> T_WLB<10> T_WLB<9> T_WLB<8> T_WLB<7> T_WLB<6> 
+ T_WLB<5> T_WLB<4> T_WLB<3> T_WLB<2> T_WLB<1> T_WLB<0> VDD VSS  / dpram16x4096_SingleCOL2X8_ROWX256
XCOL2<0>
+ RB_CA<3> RB_CA<2> RB_CA<1> RB_CA<0> RB_CB<3> RB_CB<2> RB_CB<1> RB_CB<0> RB_MA<3> 
+ RB_MA<2> RB_MA<1> RB_MA<0> RB_MB<3> RB_MB<2> RB_MB<1> RB_MB<0> RB_TM_PREB_N RB_TM_PREA_N 
+ B_WLA<255> B_WLA<254> B_WLA<253> B_WLA<252> B_WLA<251> B_WLA<250> B_WLA<249> B_WLA<248> B_WLA<247> 
+ B_WLA<246> B_WLA<245> B_WLA<244> B_WLA<243> B_WLA<242> B_WLA<241> B_WLA<240> B_WLA<239> B_WLA<238> 
+ B_WLA<237> B_WLA<236> B_WLA<235> B_WLA<234> B_WLA<233> B_WLA<232> B_WLA<231> B_WLA<230> B_WLA<229> 
+ B_WLA<228> B_WLA<227> B_WLA<226> B_WLA<225> B_WLA<224> B_WLA<223> B_WLA<222> B_WLA<221> B_WLA<220> 
+ B_WLA<219> B_WLA<218> B_WLA<217> B_WLA<216> B_WLA<215> B_WLA<214> B_WLA<213> B_WLA<212> B_WLA<211> 
+ B_WLA<210> B_WLA<209> B_WLA<208> B_WLA<207> B_WLA<206> B_WLA<205> B_WLA<204> B_WLA<203> B_WLA<202> 
+ B_WLA<201> B_WLA<200> B_WLA<199> B_WLA<198> B_WLA<197> B_WLA<196> B_WLA<195> B_WLA<194> B_WLA<193> 
+ B_WLA<192> B_WLA<191> B_WLA<190> B_WLA<189> B_WLA<188> B_WLA<187> B_WLA<186> B_WLA<185> B_WLA<184> 
+ B_WLA<183> B_WLA<182> B_WLA<181> B_WLA<180> B_WLA<179> B_WLA<178> B_WLA<177> B_WLA<176> B_WLA<175> 
+ B_WLA<174> B_WLA<173> B_WLA<172> B_WLA<171> B_WLA<170> B_WLA<169> B_WLA<168> B_WLA<167> B_WLA<166> 
+ B_WLA<165> B_WLA<164> B_WLA<163> B_WLA<162> B_WLA<161> B_WLA<160> B_WLA<159> B_WLA<158> B_WLA<157> 
+ B_WLA<156> B_WLA<155> B_WLA<154> B_WLA<153> B_WLA<152> B_WLA<151> B_WLA<150> B_WLA<149> B_WLA<148> 
+ B_WLA<147> B_WLA<146> B_WLA<145> B_WLA<144> B_WLA<143> B_WLA<142> B_WLA<141> B_WLA<140> B_WLA<139> 
+ B_WLA<138> B_WLA<137> B_WLA<136> B_WLA<135> B_WLA<134> B_WLA<133> B_WLA<132> B_WLA<131> B_WLA<130> 
+ B_WLA<129> B_WLA<128> B_WLA<127> B_WLA<126> B_WLA<125> B_WLA<124> B_WLA<123> B_WLA<122> B_WLA<121> 
+ B_WLA<120> B_WLA<119> B_WLA<118> B_WLA<117> B_WLA<116> B_WLA<115> B_WLA<114> B_WLA<113> B_WLA<112> 
+ B_WLA<111> B_WLA<110> B_WLA<109> B_WLA<108> B_WLA<107> B_WLA<106> B_WLA<105> B_WLA<104> B_WLA<103> 
+ B_WLA<102> B_WLA<101> B_WLA<100> B_WLA<99> B_WLA<98> B_WLA<97> B_WLA<96> B_WLA<95> B_WLA<94> 
+ B_WLA<93> B_WLA<92> B_WLA<91> B_WLA<90> B_WLA<89> B_WLA<88> B_WLA<87> B_WLA<86> B_WLA<85> 
+ B_WLA<84> B_WLA<83> B_WLA<82> B_WLA<81> B_WLA<80> B_WLA<79> B_WLA<78> B_WLA<77> B_WLA<76> 
+ B_WLA<75> B_WLA<74> B_WLA<73> B_WLA<72> B_WLA<71> B_WLA<70> B_WLA<69> B_WLA<68> B_WLA<67> 
+ B_WLA<66> B_WLA<65> B_WLA<64> B_WLA<63> B_WLA<62> B_WLA<61> B_WLA<60> B_WLA<59> B_WLA<58> 
+ B_WLA<57> B_WLA<56> B_WLA<55> B_WLA<54> B_WLA<53> B_WLA<52> B_WLA<51> B_WLA<50> B_WLA<49> 
+ B_WLA<48> B_WLA<47> B_WLA<46> B_WLA<45> B_WLA<44> B_WLA<43> B_WLA<42> B_WLA<41> B_WLA<40> 
+ B_WLA<39> B_WLA<38> B_WLA<37> B_WLA<36> B_WLA<35> B_WLA<34> B_WLA<33> B_WLA<32> B_WLA<31> 
+ B_WLA<30> B_WLA<29> B_WLA<28> B_WLA<27> B_WLA<26> B_WLA<25> B_WLA<24> B_WLA<23> B_WLA<22> 
+ B_WLA<21> B_WLA<20> B_WLA<19> B_WLA<18> B_WLA<17> B_WLA<16> B_WLA<15> B_WLA<14> B_WLA<13> 
+ B_WLA<12> B_WLA<11> B_WLA<10> B_WLA<9> B_WLA<8> B_WLA<7> B_WLA<6> B_WLA<5> B_WLA<4> 
+ B_WLA<3> B_WLA<2> B_WLA<1> B_WLA<0> B_WLB<255> B_WLB<254> B_WLB<253> B_WLB<252> B_WLB<251> 
+ B_WLB<250> B_WLB<249> B_WLB<248> B_WLB<247> B_WLB<246> B_WLB<245> B_WLB<244> B_WLB<243> B_WLB<242> 
+ B_WLB<241> B_WLB<240> B_WLB<239> B_WLB<238> B_WLB<237> B_WLB<236> B_WLB<235> B_WLB<234> B_WLB<233> 
+ B_WLB<232> B_WLB<231> B_WLB<230> B_WLB<229> B_WLB<228> B_WLB<227> B_WLB<226> B_WLB<225> B_WLB<224> 
+ B_WLB<223> B_WLB<222> B_WLB<221> B_WLB<220> B_WLB<219> B_WLB<218> B_WLB<217> B_WLB<216> B_WLB<215> 
+ B_WLB<214> B_WLB<213> B_WLB<212> B_WLB<211> B_WLB<210> B_WLB<209> B_WLB<208> B_WLB<207> B_WLB<206> 
+ B_WLB<205> B_WLB<204> B_WLB<203> B_WLB<202> B_WLB<201> B_WLB<200> B_WLB<199> B_WLB<198> B_WLB<197> 
+ B_WLB<196> B_WLB<195> B_WLB<194> B_WLB<193> B_WLB<192> B_WLB<191> B_WLB<190> B_WLB<189> B_WLB<188> 
+ B_WLB<187> B_WLB<186> B_WLB<185> B_WLB<184> B_WLB<183> B_WLB<182> B_WLB<181> B_WLB<180> B_WLB<179> 
+ B_WLB<178> B_WLB<177> B_WLB<176> B_WLB<175> B_WLB<174> B_WLB<173> B_WLB<172> B_WLB<171> B_WLB<170> 
+ B_WLB<169> B_WLB<168> B_WLB<167> B_WLB<166> B_WLB<165> B_WLB<164> B_WLB<163> B_WLB<162> B_WLB<161> 
+ B_WLB<160> B_WLB<159> B_WLB<158> B_WLB<157> B_WLB<156> B_WLB<155> B_WLB<154> B_WLB<153> B_WLB<152> 
+ B_WLB<151> B_WLB<150> B_WLB<149> B_WLB<148> B_WLB<147> B_WLB<146> B_WLB<145> B_WLB<144> B_WLB<143> 
+ B_WLB<142> B_WLB<141> B_WLB<140> B_WLB<139> B_WLB<138> B_WLB<137> B_WLB<136> B_WLB<135> B_WLB<134> 
+ B_WLB<133> B_WLB<132> B_WLB<131> B_WLB<130> B_WLB<129> B_WLB<128> B_WLB<127> B_WLB<126> B_WLB<125> 
+ B_WLB<124> B_WLB<123> B_WLB<122> B_WLB<121> B_WLB<120> B_WLB<119> B_WLB<118> B_WLB<117> B_WLB<116> 
+ B_WLB<115> B_WLB<114> B_WLB<113> B_WLB<112> B_WLB<111> B_WLB<110> B_WLB<109> B_WLB<108> B_WLB<107> 
+ B_WLB<106> B_WLB<105> B_WLB<104> B_WLB<103> B_WLB<102> B_WLB<101> B_WLB<100> B_WLB<99> B_WLB<98> 
+ B_WLB<97> B_WLB<96> B_WLB<95> B_WLB<94> B_WLB<93> B_WLB<92> B_WLB<91> B_WLB<90> B_WLB<89> 
+ B_WLB<88> B_WLB<87> B_WLB<86> B_WLB<85> B_WLB<84> B_WLB<83> B_WLB<82> B_WLB<81> B_WLB<80> 
+ B_WLB<79> B_WLB<78> B_WLB<77> B_WLB<76> B_WLB<75> B_WLB<74> B_WLB<73> B_WLB<72> B_WLB<71> 
+ B_WLB<70> B_WLB<69> B_WLB<68> B_WLB<67> B_WLB<66> B_WLB<65> B_WLB<64> B_WLB<63> B_WLB<62> 
+ B_WLB<61> B_WLB<60> B_WLB<59> B_WLB<58> B_WLB<57> B_WLB<56> B_WLB<55> B_WLB<54> B_WLB<53> 
+ B_WLB<52> B_WLB<51> B_WLB<50> B_WLB<49> B_WLB<48> B_WLB<47> B_WLB<46> B_WLB<45> B_WLB<44> 
+ B_WLB<43> B_WLB<42> B_WLB<41> B_WLB<40> B_WLB<39> B_WLB<38> B_WLB<37> B_WLB<36> B_WLB<35> 
+ B_WLB<34> B_WLB<33> B_WLB<32> B_WLB<31> B_WLB<30> B_WLB<29> B_WLB<28> B_WLB<27> B_WLB<26> 
+ B_WLB<25> B_WLB<24> B_WLB<23> B_WLB<22> B_WLB<21> B_WLB<20> B_WLB<19> B_WLB<18> B_WLB<17> 
+ B_WLB<16> B_WLB<15> B_WLB<14> B_WLB<13> B_WLB<12> B_WLB<11> B_WLB<10> B_WLB<9> B_WLB<8> 
+ B_WLB<7> B_WLB<6> B_WLB<5> B_WLB<4> B_WLB<3> B_WLB<2> B_WLB<1> B_WLB<0> BWENA<1> 
+ BWENA<0> BWENB<1> BWENB<0> R_CLK_DQA R_CLK_DQA_N R_CLK_DQB R_CLK_DQB_N DA<1> DA<0> 
+ DB<1> DB<0> DDQA<0> DDQA_N<0> DDQB<0> DDQB_N<0> R_LWEA R_LWEB QA<1> 
+ QA<0> QB<1> QB<0> R_SA_PREA_N R_SA_PREB_N R_SAEA_N R_SAEB_N RT_CA<3> RT_CA<2> 
+ RT_CA<1> RT_CA<0> RT_CB<3> RT_CB<2> RT_CB<1> RT_CB<0> RT_MA<3> RT_MA<2> RT_MA<1> 
+ RT_MA<0> RT_MB<3> RT_MB<2> RT_MB<1> RT_MB<0> R_TM_PREA_N R_TM_PREB_N T_WLA<255> T_WLA<254> 
+ T_WLA<253> T_WLA<252> T_WLA<251> T_WLA<250> T_WLA<249> T_WLA<248> T_WLA<247> T_WLA<246> T_WLA<245> 
+ T_WLA<244> T_WLA<243> T_WLA<242> T_WLA<241> T_WLA<240> T_WLA<239> T_WLA<238> T_WLA<237> T_WLA<236> 
+ T_WLA<235> T_WLA<234> T_WLA<233> T_WLA<232> T_WLA<231> T_WLA<230> T_WLA<229> T_WLA<228> T_WLA<227> 
+ T_WLA<226> T_WLA<225> T_WLA<224> T_WLA<223> T_WLA<222> T_WLA<221> T_WLA<220> T_WLA<219> T_WLA<218> 
+ T_WLA<217> T_WLA<216> T_WLA<215> T_WLA<214> T_WLA<213> T_WLA<212> T_WLA<211> T_WLA<210> T_WLA<209> 
+ T_WLA<208> T_WLA<207> T_WLA<206> T_WLA<205> T_WLA<204> T_WLA<203> T_WLA<202> T_WLA<201> T_WLA<200> 
+ T_WLA<199> T_WLA<198> T_WLA<197> T_WLA<196> T_WLA<195> T_WLA<194> T_WLA<193> T_WLA<192> T_WLA<191> 
+ T_WLA<190> T_WLA<189> T_WLA<188> T_WLA<187> T_WLA<186> T_WLA<185> T_WLA<184> T_WLA<183> T_WLA<182> 
+ T_WLA<181> T_WLA<180> T_WLA<179> T_WLA<178> T_WLA<177> T_WLA<176> T_WLA<175> T_WLA<174> T_WLA<173> 
+ T_WLA<172> T_WLA<171> T_WLA<170> T_WLA<169> T_WLA<168> T_WLA<167> T_WLA<166> T_WLA<165> T_WLA<164> 
+ T_WLA<163> T_WLA<162> T_WLA<161> T_WLA<160> T_WLA<159> T_WLA<158> T_WLA<157> T_WLA<156> T_WLA<155> 
+ T_WLA<154> T_WLA<153> T_WLA<152> T_WLA<151> T_WLA<150> T_WLA<149> T_WLA<148> T_WLA<147> T_WLA<146> 
+ T_WLA<145> T_WLA<144> T_WLA<143> T_WLA<142> T_WLA<141> T_WLA<140> T_WLA<139> T_WLA<138> T_WLA<137> 
+ T_WLA<136> T_WLA<135> T_WLA<134> T_WLA<133> T_WLA<132> T_WLA<131> T_WLA<130> T_WLA<129> T_WLA<128> 
+ T_WLA<127> T_WLA<126> T_WLA<125> T_WLA<124> T_WLA<123> T_WLA<122> T_WLA<121> T_WLA<120> T_WLA<119> 
+ T_WLA<118> T_WLA<117> T_WLA<116> T_WLA<115> T_WLA<114> T_WLA<113> T_WLA<112> T_WLA<111> T_WLA<110> 
+ T_WLA<109> T_WLA<108> T_WLA<107> T_WLA<106> T_WLA<105> T_WLA<104> T_WLA<103> T_WLA<102> T_WLA<101> 
+ T_WLA<100> T_WLA<99> T_WLA<98> T_WLA<97> T_WLA<96> T_WLA<95> T_WLA<94> T_WLA<93> T_WLA<92> 
+ T_WLA<91> T_WLA<90> T_WLA<89> T_WLA<88> T_WLA<87> T_WLA<86> T_WLA<85> T_WLA<84> T_WLA<83> 
+ T_WLA<82> T_WLA<81> T_WLA<80> T_WLA<79> T_WLA<78> T_WLA<77> T_WLA<76> T_WLA<75> T_WLA<74> 
+ T_WLA<73> T_WLA<72> T_WLA<71> T_WLA<70> T_WLA<69> T_WLA<68> T_WLA<67> T_WLA<66> T_WLA<65> 
+ T_WLA<64> T_WLA<63> T_WLA<62> T_WLA<61> T_WLA<60> T_WLA<59> T_WLA<58> T_WLA<57> T_WLA<56> 
+ T_WLA<55> T_WLA<54> T_WLA<53> T_WLA<52> T_WLA<51> T_WLA<50> T_WLA<49> T_WLA<48> T_WLA<47> 
+ T_WLA<46> T_WLA<45> T_WLA<44> T_WLA<43> T_WLA<42> T_WLA<41> T_WLA<40> T_WLA<39> T_WLA<38> 
+ T_WLA<37> T_WLA<36> T_WLA<35> T_WLA<34> T_WLA<33> T_WLA<32> T_WLA<31> T_WLA<30> T_WLA<29> 
+ T_WLA<28> T_WLA<27> T_WLA<26> T_WLA<25> T_WLA<24> T_WLA<23> T_WLA<22> T_WLA<21> T_WLA<20> 
+ T_WLA<19> T_WLA<18> T_WLA<17> T_WLA<16> T_WLA<15> T_WLA<14> T_WLA<13> T_WLA<12> T_WLA<11> 
+ T_WLA<10> T_WLA<9> T_WLA<8> T_WLA<7> T_WLA<6> T_WLA<5> T_WLA<4> T_WLA<3> T_WLA<2> 
+ T_WLA<1> T_WLA<0> T_WLB<255> T_WLB<254> T_WLB<253> T_WLB<252> T_WLB<251> T_WLB<250> T_WLB<249> 
+ T_WLB<248> T_WLB<247> T_WLB<246> T_WLB<245> T_WLB<244> T_WLB<243> T_WLB<242> T_WLB<241> T_WLB<240> 
+ T_WLB<239> T_WLB<238> T_WLB<237> T_WLB<236> T_WLB<235> T_WLB<234> T_WLB<233> T_WLB<232> T_WLB<231> 
+ T_WLB<230> T_WLB<229> T_WLB<228> T_WLB<227> T_WLB<226> T_WLB<225> T_WLB<224> T_WLB<223> T_WLB<222> 
+ T_WLB<221> T_WLB<220> T_WLB<219> T_WLB<218> T_WLB<217> T_WLB<216> T_WLB<215> T_WLB<214> T_WLB<213> 
+ T_WLB<212> T_WLB<211> T_WLB<210> T_WLB<209> T_WLB<208> T_WLB<207> T_WLB<206> T_WLB<205> T_WLB<204> 
+ T_WLB<203> T_WLB<202> T_WLB<201> T_WLB<200> T_WLB<199> T_WLB<198> T_WLB<197> T_WLB<196> T_WLB<195> 
+ T_WLB<194> T_WLB<193> T_WLB<192> T_WLB<191> T_WLB<190> T_WLB<189> T_WLB<188> T_WLB<187> T_WLB<186> 
+ T_WLB<185> T_WLB<184> T_WLB<183> T_WLB<182> T_WLB<181> T_WLB<180> T_WLB<179> T_WLB<178> T_WLB<177> 
+ T_WLB<176> T_WLB<175> T_WLB<174> T_WLB<173> T_WLB<172> T_WLB<171> T_WLB<170> T_WLB<169> T_WLB<168> 
+ T_WLB<167> T_WLB<166> T_WLB<165> T_WLB<164> T_WLB<163> T_WLB<162> T_WLB<161> T_WLB<160> T_WLB<159> 
+ T_WLB<158> T_WLB<157> T_WLB<156> T_WLB<155> T_WLB<154> T_WLB<153> T_WLB<152> T_WLB<151> T_WLB<150> 
+ T_WLB<149> T_WLB<148> T_WLB<147> T_WLB<146> T_WLB<145> T_WLB<144> T_WLB<143> T_WLB<142> T_WLB<141> 
+ T_WLB<140> T_WLB<139> T_WLB<138> T_WLB<137> T_WLB<136> T_WLB<135> T_WLB<134> T_WLB<133> T_WLB<132> 
+ T_WLB<131> T_WLB<130> T_WLB<129> T_WLB<128> T_WLB<127> T_WLB<126> T_WLB<125> T_WLB<124> T_WLB<123> 
+ T_WLB<122> T_WLB<121> T_WLB<120> T_WLB<119> T_WLB<118> T_WLB<117> T_WLB<116> T_WLB<115> T_WLB<114> 
+ T_WLB<113> T_WLB<112> T_WLB<111> T_WLB<110> T_WLB<109> T_WLB<108> T_WLB<107> T_WLB<106> T_WLB<105> 
+ T_WLB<104> T_WLB<103> T_WLB<102> T_WLB<101> T_WLB<100> T_WLB<99> T_WLB<98> T_WLB<97> T_WLB<96> 
+ T_WLB<95> T_WLB<94> T_WLB<93> T_WLB<92> T_WLB<91> T_WLB<90> T_WLB<89> T_WLB<88> T_WLB<87> 
+ T_WLB<86> T_WLB<85> T_WLB<84> T_WLB<83> T_WLB<82> T_WLB<81> T_WLB<80> T_WLB<79> T_WLB<78> 
+ T_WLB<77> T_WLB<76> T_WLB<75> T_WLB<74> T_WLB<73> T_WLB<72> T_WLB<71> T_WLB<70> T_WLB<69> 
+ T_WLB<68> T_WLB<67> T_WLB<66> T_WLB<65> T_WLB<64> T_WLB<63> T_WLB<62> T_WLB<61> T_WLB<60> 
+ T_WLB<59> T_WLB<58> T_WLB<57> T_WLB<56> T_WLB<55> T_WLB<54> T_WLB<53> T_WLB<52> T_WLB<51> 
+ T_WLB<50> T_WLB<49> T_WLB<48> T_WLB<47> T_WLB<46> T_WLB<45> T_WLB<44> T_WLB<43> T_WLB<42> 
+ T_WLB<41> T_WLB<40> T_WLB<39> T_WLB<38> T_WLB<37> T_WLB<36> T_WLB<35> T_WLB<34> T_WLB<33> 
+ T_WLB<32> T_WLB<31> T_WLB<30> T_WLB<29> T_WLB<28> T_WLB<27> T_WLB<26> T_WLB<25> T_WLB<24> 
+ T_WLB<23> T_WLB<22> T_WLB<21> T_WLB<20> T_WLB<19> T_WLB<18> T_WLB<17> T_WLB<16> T_WLB<15> 
+ T_WLB<14> T_WLB<13> T_WLB<12> T_WLB<11> T_WLB<10> T_WLB<9> T_WLB<8> T_WLB<7> T_WLB<6> 
+ T_WLB<5> T_WLB<4> T_WLB<3> T_WLB<2> T_WLB<1> T_WLB<0> VDD VSS  / dpram16x4096_SingleCOL2X8_ROWX256
XMID
+ AA<11> AA<10> AA<9> AA<8> AA<7> AA<6> AA<5> AA<4> AA<3> 
+ TIE_VSS AA<2> AA<1> AA<0> AB<11> AB<10> AB<9> AB<8> AB<7> 
+ AB<6> AB<5> AB<4> AB<3> TIE_VSS AB<2> AB<1> AB<0> B_WLA<255> 
+ B_WLA<254> B_WLA<253> B_WLA<252> B_WLA<251> B_WLA<250> B_WLA<249> B_WLA<248> B_WLA<247> B_WLA<246> 
+ B_WLA<245> B_WLA<244> B_WLA<243> B_WLA<242> B_WLA<241> B_WLA<240> B_WLA<239> B_WLA<238> B_WLA<237> 
+ B_WLA<236> B_WLA<235> B_WLA<234> B_WLA<233> B_WLA<232> B_WLA<231> B_WLA<230> B_WLA<229> B_WLA<228> 
+ B_WLA<227> B_WLA<226> B_WLA<225> B_WLA<224> B_WLA<223> B_WLA<222> B_WLA<221> B_WLA<220> B_WLA<219> 
+ B_WLA<218> B_WLA<217> B_WLA<216> B_WLA<215> B_WLA<214> B_WLA<213> B_WLA<212> B_WLA<211> B_WLA<210> 
+ B_WLA<209> B_WLA<208> B_WLA<207> B_WLA<206> B_WLA<205> B_WLA<204> B_WLA<203> B_WLA<202> B_WLA<201> 
+ B_WLA<200> B_WLA<199> B_WLA<198> B_WLA<197> B_WLA<196> B_WLA<195> B_WLA<194> B_WLA<193> B_WLA<192> 
+ B_WLA<191> B_WLA<190> B_WLA<189> B_WLA<188> B_WLA<187> B_WLA<186> B_WLA<185> B_WLA<184> B_WLA<183> 
+ B_WLA<182> B_WLA<181> B_WLA<180> B_WLA<179> B_WLA<178> B_WLA<177> B_WLA<176> B_WLA<175> B_WLA<174> 
+ B_WLA<173> B_WLA<172> B_WLA<171> B_WLA<170> B_WLA<169> B_WLA<168> B_WLA<167> B_WLA<166> B_WLA<165> 
+ B_WLA<164> B_WLA<163> B_WLA<162> B_WLA<161> B_WLA<160> B_WLA<159> B_WLA<158> B_WLA<157> B_WLA<156> 
+ B_WLA<155> B_WLA<154> B_WLA<153> B_WLA<152> B_WLA<151> B_WLA<150> B_WLA<149> B_WLA<148> B_WLA<147> 
+ B_WLA<146> B_WLA<145> B_WLA<144> B_WLA<143> B_WLA<142> B_WLA<141> B_WLA<140> B_WLA<139> B_WLA<138> 
+ B_WLA<137> B_WLA<136> B_WLA<135> B_WLA<134> B_WLA<133> B_WLA<132> B_WLA<131> B_WLA<130> B_WLA<129> 
+ B_WLA<128> B_WLA<127> B_WLA<126> B_WLA<125> B_WLA<124> B_WLA<123> B_WLA<122> B_WLA<121> B_WLA<120> 
+ B_WLA<119> B_WLA<118> B_WLA<117> B_WLA<116> B_WLA<115> B_WLA<114> B_WLA<113> B_WLA<112> B_WLA<111> 
+ B_WLA<110> B_WLA<109> B_WLA<108> B_WLA<107> B_WLA<106> B_WLA<105> B_WLA<104> B_WLA<103> B_WLA<102> 
+ B_WLA<101> B_WLA<100> B_WLA<99> B_WLA<98> B_WLA<97> B_WLA<96> B_WLA<95> B_WLA<94> B_WLA<93> 
+ B_WLA<92> B_WLA<91> B_WLA<90> B_WLA<89> B_WLA<88> B_WLA<87> B_WLA<86> B_WLA<85> B_WLA<84> 
+ B_WLA<83> B_WLA<82> B_WLA<81> B_WLA<80> B_WLA<79> B_WLA<78> B_WLA<77> B_WLA<76> B_WLA<75> 
+ B_WLA<74> B_WLA<73> B_WLA<72> B_WLA<71> B_WLA<70> B_WLA<69> B_WLA<68> B_WLA<67> B_WLA<66> 
+ B_WLA<65> B_WLA<64> B_WLA<63> B_WLA<62> B_WLA<61> B_WLA<60> B_WLA<59> B_WLA<58> B_WLA<57> 
+ B_WLA<56> B_WLA<55> B_WLA<54> B_WLA<53> B_WLA<52> B_WLA<51> B_WLA<50> B_WLA<49> B_WLA<48> 
+ B_WLA<47> B_WLA<46> B_WLA<45> B_WLA<44> B_WLA<43> B_WLA<42> B_WLA<41> B_WLA<40> B_WLA<39> 
+ B_WLA<38> B_WLA<37> B_WLA<36> B_WLA<35> B_WLA<34> B_WLA<33> B_WLA<32> B_WLA<31> B_WLA<30> 
+ B_WLA<29> B_WLA<28> B_WLA<27> B_WLA<26> B_WLA<25> B_WLA<24> B_WLA<23> B_WLA<22> B_WLA<21> 
+ B_WLA<20> B_WLA<19> B_WLA<18> B_WLA<17> B_WLA<16> B_WLA<15> B_WLA<14> B_WLA<13> B_WLA<12> 
+ B_WLA<11> B_WLA<10> B_WLA<9> B_WLA<8> B_WLA<7> B_WLA<6> B_WLA<5> B_WLA<4> B_WLA<3> 
+ B_WLA<2> B_WLA<1> B_WLA<0> B_WLB<255> B_WLB<254> B_WLB<253> B_WLB<252> B_WLB<251> B_WLB<250> 
+ B_WLB<249> B_WLB<248> B_WLB<247> B_WLB<246> B_WLB<245> B_WLB<244> B_WLB<243> B_WLB<242> B_WLB<241> 
+ B_WLB<240> B_WLB<239> B_WLB<238> B_WLB<237> B_WLB<236> B_WLB<235> B_WLB<234> B_WLB<233> B_WLB<232> 
+ B_WLB<231> B_WLB<230> B_WLB<229> B_WLB<228> B_WLB<227> B_WLB<226> B_WLB<225> B_WLB<224> B_WLB<223> 
+ B_WLB<222> B_WLB<221> B_WLB<220> B_WLB<219> B_WLB<218> B_WLB<217> B_WLB<216> B_WLB<215> B_WLB<214> 
+ B_WLB<213> B_WLB<212> B_WLB<211> B_WLB<210> B_WLB<209> B_WLB<208> B_WLB<207> B_WLB<206> B_WLB<205> 
+ B_WLB<204> B_WLB<203> B_WLB<202> B_WLB<201> B_WLB<200> B_WLB<199> B_WLB<198> B_WLB<197> B_WLB<196> 
+ B_WLB<195> B_WLB<194> B_WLB<193> B_WLB<192> B_WLB<191> B_WLB<190> B_WLB<189> B_WLB<188> B_WLB<187> 
+ B_WLB<186> B_WLB<185> B_WLB<184> B_WLB<183> B_WLB<182> B_WLB<181> B_WLB<180> B_WLB<179> B_WLB<178> 
+ B_WLB<177> B_WLB<176> B_WLB<175> B_WLB<174> B_WLB<173> B_WLB<172> B_WLB<171> B_WLB<170> B_WLB<169> 
+ B_WLB<168> B_WLB<167> B_WLB<166> B_WLB<165> B_WLB<164> B_WLB<163> B_WLB<162> B_WLB<161> B_WLB<160> 
+ B_WLB<159> B_WLB<158> B_WLB<157> B_WLB<156> B_WLB<155> B_WLB<154> B_WLB<153> B_WLB<152> B_WLB<151> 
+ B_WLB<150> B_WLB<149> B_WLB<148> B_WLB<147> B_WLB<146> B_WLB<145> B_WLB<144> B_WLB<143> B_WLB<142> 
+ B_WLB<141> B_WLB<140> B_WLB<139> B_WLB<138> B_WLB<137> B_WLB<136> B_WLB<135> B_WLB<134> B_WLB<133> 
+ B_WLB<132> B_WLB<131> B_WLB<130> B_WLB<129> B_WLB<128> B_WLB<127> B_WLB<126> B_WLB<125> B_WLB<124> 
+ B_WLB<123> B_WLB<122> B_WLB<121> B_WLB<120> B_WLB<119> B_WLB<118> B_WLB<117> B_WLB<116> B_WLB<115> 
+ B_WLB<114> B_WLB<113> B_WLB<112> B_WLB<111> B_WLB<110> B_WLB<109> B_WLB<108> B_WLB<107> B_WLB<106> 
+ B_WLB<105> B_WLB<104> B_WLB<103> B_WLB<102> B_WLB<101> B_WLB<100> B_WLB<99> B_WLB<98> B_WLB<97> 
+ B_WLB<96> B_WLB<95> B_WLB<94> B_WLB<93> B_WLB<92> B_WLB<91> B_WLB<90> B_WLB<89> B_WLB<88> 
+ B_WLB<87> B_WLB<86> B_WLB<85> B_WLB<84> B_WLB<83> B_WLB<82> B_WLB<81> B_WLB<80> B_WLB<79> 
+ B_WLB<78> B_WLB<77> B_WLB<76> B_WLB<75> B_WLB<74> B_WLB<73> B_WLB<72> B_WLB<71> B_WLB<70> 
+ B_WLB<69> B_WLB<68> B_WLB<67> B_WLB<66> B_WLB<65> B_WLB<64> B_WLB<63> B_WLB<62> B_WLB<61> 
+ B_WLB<60> B_WLB<59> B_WLB<58> B_WLB<57> B_WLB<56> B_WLB<55> B_WLB<54> B_WLB<53> B_WLB<52> 
+ B_WLB<51> B_WLB<50> B_WLB<49> B_WLB<48> B_WLB<47> B_WLB<46> B_WLB<45> B_WLB<44> B_WLB<43> 
+ B_WLB<42> B_WLB<41> B_WLB<40> B_WLB<39> B_WLB<38> B_WLB<37> B_WLB<36> B_WLB<35> B_WLB<34> 
+ B_WLB<33> B_WLB<32> B_WLB<31> B_WLB<30> B_WLB<29> B_WLB<28> B_WLB<27> B_WLB<26> B_WLB<25> 
+ B_WLB<24> B_WLB<23> B_WLB<22> B_WLB<21> B_WLB<20> B_WLB<19> B_WLB<18> B_WLB<17> B_WLB<16> 
+ B_WLB<15> B_WLB<14> B_WLB<13> B_WLB<12> B_WLB<11> B_WLB<10> B_WLB<9> B_WLB<8> B_WLB<7> 
+ B_WLB<6> B_WLB<5> B_WLB<4> B_WLB<3> B_WLB<2> B_WLB<1> B_WLB<0> CENA CENB 
+ CLKA CLKB DBL_PD_N<3> DBL_PD_N<2> DBL_PD_N<1> DBL_PD_N<0> DDQA<3> DDQA_N<3> DDQB<4> 
+ DDQB_N<4> DWLA<1> DWLA<0> DWLB<1> DWLB<0> L_CLK_DQA L_CLK_DQA_N L_CLK_DQB L_CLK_DQB_N 
+ L_LWEA L_LWEB L_SA_PREA_N L_SA_PREB_N L_SAEA_N L_SAEB_N LB_CA<3> LB_CA<2> LB_CA<1> 
+ LB_CA<0> LB_CB<3> LB_CB<2> LB_CB<1> LB_CB<0> LB_MA<3> LB_MA<2> LB_MA<1> LB_MA<0> 
+ LB_MB<3> LB_MB<2> LB_MB<1> LB_MB<0> LB_TM_PREA_N LB_TM_PREB_N LT_CA<3> LT_CA<2> LT_CA<1> 
+ LT_CA<0> LT_CB<3> LT_CB<2> LT_CB<1> LT_CB<0> LT_MA<3> LT_MA<2> LT_MA<1> LT_MA<0> 
+ LT_MB<3> LT_MB<2> LT_MB<1> LT_MB<0> LT_TM_PREA_N LT_TM_PREB_N R_CLK_DQA R_CLK_DQA_N R_CLK_DQB 
+ R_CLK_DQB_N R_LWEA R_LWEB R_SA_PREA_N R_SA_PREB_N R_SAEA_N R_SAEB_N RB_CA<3> RB_CA<2> 
+ RB_CA<1> RB_CA<0> RB_CB<3> RB_CB<2> RB_CB<1> RB_CB<0> RB_MA<3> RB_MA<2> RB_MA<1> 
+ RB_MA<0> RB_MB<3> RB_MB<2> RB_MB<1> RB_MB<0> RB_TM_PREB_N RB_TM_PREA_N RT_CA<3> RT_CA<2> 
+ RT_CA<1> RT_CA<0> RT_CB<3> RT_CB<2> RT_CB<1> RT_CB<0> RT_MA<3> RT_MA<2> RT_MA<1> 
+ RT_MA<0> RT_MB<3> RT_MB<2> RT_MB<1> RT_MB<0> R_TM_PREA_N R_TM_PREB_N STCLKA STCLKB 
+ T_WLA<255> T_WLA<254> T_WLA<253> T_WLA<252> T_WLA<251> T_WLA<250> T_WLA<249> T_WLA<248> T_WLA<247> 
+ T_WLA<246> T_WLA<245> T_WLA<244> T_WLA<243> T_WLA<242> T_WLA<241> T_WLA<240> T_WLA<239> T_WLA<238> 
+ T_WLA<237> T_WLA<236> T_WLA<235> T_WLA<234> T_WLA<233> T_WLA<232> T_WLA<231> T_WLA<230> T_WLA<229> 
+ T_WLA<228> T_WLA<227> T_WLA<226> T_WLA<225> T_WLA<224> T_WLA<223> T_WLA<222> T_WLA<221> T_WLA<220> 
+ T_WLA<219> T_WLA<218> T_WLA<217> T_WLA<216> T_WLA<215> T_WLA<214> T_WLA<213> T_WLA<212> T_WLA<211> 
+ T_WLA<210> T_WLA<209> T_WLA<208> T_WLA<207> T_WLA<206> T_WLA<205> T_WLA<204> T_WLA<203> T_WLA<202> 
+ T_WLA<201> T_WLA<200> T_WLA<199> T_WLA<198> T_WLA<197> T_WLA<196> T_WLA<195> T_WLA<194> T_WLA<193> 
+ T_WLA<192> T_WLA<191> T_WLA<190> T_WLA<189> T_WLA<188> T_WLA<187> T_WLA<186> T_WLA<185> T_WLA<184> 
+ T_WLA<183> T_WLA<182> T_WLA<181> T_WLA<180> T_WLA<179> T_WLA<178> T_WLA<177> T_WLA<176> T_WLA<175> 
+ T_WLA<174> T_WLA<173> T_WLA<172> T_WLA<171> T_WLA<170> T_WLA<169> T_WLA<168> T_WLA<167> T_WLA<166> 
+ T_WLA<165> T_WLA<164> T_WLA<163> T_WLA<162> T_WLA<161> T_WLA<160> T_WLA<159> T_WLA<158> T_WLA<157> 
+ T_WLA<156> T_WLA<155> T_WLA<154> T_WLA<153> T_WLA<152> T_WLA<151> T_WLA<150> T_WLA<149> T_WLA<148> 
+ T_WLA<147> T_WLA<146> T_WLA<145> T_WLA<144> T_WLA<143> T_WLA<142> T_WLA<141> T_WLA<140> T_WLA<139> 
+ T_WLA<138> T_WLA<137> T_WLA<136> T_WLA<135> T_WLA<134> T_WLA<133> T_WLA<132> T_WLA<131> T_WLA<130> 
+ T_WLA<129> T_WLA<128> T_WLA<127> T_WLA<126> T_WLA<125> T_WLA<124> T_WLA<123> T_WLA<122> T_WLA<121> 
+ T_WLA<120> T_WLA<119> T_WLA<118> T_WLA<117> T_WLA<116> T_WLA<115> T_WLA<114> T_WLA<113> T_WLA<112> 
+ T_WLA<111> T_WLA<110> T_WLA<109> T_WLA<108> T_WLA<107> T_WLA<106> T_WLA<105> T_WLA<104> T_WLA<103> 
+ T_WLA<102> T_WLA<101> T_WLA<100> T_WLA<99> T_WLA<98> T_WLA<97> T_WLA<96> T_WLA<95> T_WLA<94> 
+ T_WLA<93> T_WLA<92> T_WLA<91> T_WLA<90> T_WLA<89> T_WLA<88> T_WLA<87> T_WLA<86> T_WLA<85> 
+ T_WLA<84> T_WLA<83> T_WLA<82> T_WLA<81> T_WLA<80> T_WLA<79> T_WLA<78> T_WLA<77> T_WLA<76> 
+ T_WLA<75> T_WLA<74> T_WLA<73> T_WLA<72> T_WLA<71> T_WLA<70> T_WLA<69> T_WLA<68> T_WLA<67> 
+ T_WLA<66> T_WLA<65> T_WLA<64> T_WLA<63> T_WLA<62> T_WLA<61> T_WLA<60> T_WLA<59> T_WLA<58> 
+ T_WLA<57> T_WLA<56> T_WLA<55> T_WLA<54> T_WLA<53> T_WLA<52> T_WLA<51> T_WLA<50> T_WLA<49> 
+ T_WLA<48> T_WLA<47> T_WLA<46> T_WLA<45> T_WLA<44> T_WLA<43> T_WLA<42> T_WLA<41> T_WLA<40> 
+ T_WLA<39> T_WLA<38> T_WLA<37> T_WLA<36> T_WLA<35> T_WLA<34> T_WLA<33> T_WLA<32> T_WLA<31> 
+ T_WLA<30> T_WLA<29> T_WLA<28> T_WLA<27> T_WLA<26> T_WLA<25> T_WLA<24> T_WLA<23> T_WLA<22> 
+ T_WLA<21> T_WLA<20> T_WLA<19> T_WLA<18> T_WLA<17> T_WLA<16> T_WLA<15> T_WLA<14> T_WLA<13> 
+ T_WLA<12> T_WLA<11> T_WLA<10> T_WLA<9> T_WLA<8> T_WLA<7> T_WLA<6> T_WLA<5> T_WLA<4> 
+ T_WLA<3> T_WLA<2> T_WLA<1> T_WLA<0> T_WLB<255> T_WLB<254> T_WLB<253> T_WLB<252> T_WLB<251> 
+ T_WLB<250> T_WLB<249> T_WLB<248> T_WLB<247> T_WLB<246> T_WLB<245> T_WLB<244> T_WLB<243> T_WLB<242> 
+ T_WLB<241> T_WLB<240> T_WLB<239> T_WLB<238> T_WLB<237> T_WLB<236> T_WLB<235> T_WLB<234> T_WLB<233> 
+ T_WLB<232> T_WLB<231> T_WLB<230> T_WLB<229> T_WLB<228> T_WLB<227> T_WLB<226> T_WLB<225> T_WLB<224> 
+ T_WLB<223> T_WLB<222> T_WLB<221> T_WLB<220> T_WLB<219> T_WLB<218> T_WLB<217> T_WLB<216> T_WLB<215> 
+ T_WLB<214> T_WLB<213> T_WLB<212> T_WLB<211> T_WLB<210> T_WLB<209> T_WLB<208> T_WLB<207> T_WLB<206> 
+ T_WLB<205> T_WLB<204> T_WLB<203> T_WLB<202> T_WLB<201> T_WLB<200> T_WLB<199> T_WLB<198> T_WLB<197> 
+ T_WLB<196> T_WLB<195> T_WLB<194> T_WLB<193> T_WLB<192> T_WLB<191> T_WLB<190> T_WLB<189> T_WLB<188> 
+ T_WLB<187> T_WLB<186> T_WLB<185> T_WLB<184> T_WLB<183> T_WLB<182> T_WLB<181> T_WLB<180> T_WLB<179> 
+ T_WLB<178> T_WLB<177> T_WLB<176> T_WLB<175> T_WLB<174> T_WLB<173> T_WLB<172> T_WLB<171> T_WLB<170> 
+ T_WLB<169> T_WLB<168> T_WLB<167> T_WLB<166> T_WLB<165> T_WLB<164> T_WLB<163> T_WLB<162> T_WLB<161> 
+ T_WLB<160> T_WLB<159> T_WLB<158> T_WLB<157> T_WLB<156> T_WLB<155> T_WLB<154> T_WLB<153> T_WLB<152> 
+ T_WLB<151> T_WLB<150> T_WLB<149> T_WLB<148> T_WLB<147> T_WLB<146> T_WLB<145> T_WLB<144> T_WLB<143> 
+ T_WLB<142> T_WLB<141> T_WLB<140> T_WLB<139> T_WLB<138> T_WLB<137> T_WLB<136> T_WLB<135> T_WLB<134> 
+ T_WLB<133> T_WLB<132> T_WLB<131> T_WLB<130> T_WLB<129> T_WLB<128> T_WLB<127> T_WLB<126> T_WLB<125> 
+ T_WLB<124> T_WLB<123> T_WLB<122> T_WLB<121> T_WLB<120> T_WLB<119> T_WLB<118> T_WLB<117> T_WLB<116> 
+ T_WLB<115> T_WLB<114> T_WLB<113> T_WLB<112> T_WLB<111> T_WLB<110> T_WLB<109> T_WLB<108> T_WLB<107> 
+ T_WLB<106> T_WLB<105> T_WLB<104> T_WLB<103> T_WLB<102> T_WLB<101> T_WLB<100> T_WLB<99> T_WLB<98> 
+ T_WLB<97> T_WLB<96> T_WLB<95> T_WLB<94> T_WLB<93> T_WLB<92> T_WLB<91> T_WLB<90> T_WLB<89> 
+ T_WLB<88> T_WLB<87> T_WLB<86> T_WLB<85> T_WLB<84> T_WLB<83> T_WLB<82> T_WLB<81> T_WLB<80> 
+ T_WLB<79> T_WLB<78> T_WLB<77> T_WLB<76> T_WLB<75> T_WLB<74> T_WLB<73> T_WLB<72> T_WLB<71> 
+ T_WLB<70> T_WLB<69> T_WLB<68> T_WLB<67> T_WLB<66> T_WLB<65> T_WLB<64> T_WLB<63> T_WLB<62> 
+ T_WLB<61> T_WLB<60> T_WLB<59> T_WLB<58> T_WLB<57> T_WLB<56> T_WLB<55> T_WLB<54> T_WLB<53> 
+ T_WLB<52> T_WLB<51> T_WLB<50> T_WLB<49> T_WLB<48> T_WLB<47> T_WLB<46> T_WLB<45> T_WLB<44> 
+ T_WLB<43> T_WLB<42> T_WLB<41> T_WLB<40> T_WLB<39> T_WLB<38> T_WLB<37> T_WLB<36> T_WLB<35> 
+ T_WLB<34> T_WLB<33> T_WLB<32> T_WLB<31> T_WLB<30> T_WLB<29> T_WLB<28> T_WLB<27> T_WLB<26> 
+ T_WLB<25> T_WLB<24> T_WLB<23> T_WLB<22> T_WLB<21> T_WLB<20> T_WLB<19> T_WLB<18> T_WLB<17> 
+ T_WLB<16> T_WLB<15> T_WLB<14> T_WLB<13> T_WLB<12> T_WLB<11> T_WLB<10> T_WLB<9> T_WLB<8> 
+ T_WLB<7> T_WLB<6> T_WLB<5> T_WLB<4> T_WLB<3> T_WLB<2> T_WLB<1> T_WLB<0> TIE_VDD 
+ TIE_VSS TIE_VSS TIE_VSS TIE_VSS TIE_VSS TIE_VSS TIE_VSS TIE_VSS TIE_VSS 
+ TIE_VSS TIE_VSS VDD VSS WENA WENB  / dpram16x4096_MIDX8_ROWX256
.ENDS

