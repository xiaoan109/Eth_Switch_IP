// removed module with interface ports: DcpRdData16x16
