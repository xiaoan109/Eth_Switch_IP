// removed module with interface ports: DcpWrrArbiter
