VERSION 5.6 ;
NAMESCASESENSITIVE ON ; 
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

#Instance Name:  dpram16x4096
#Word Depth:     4096
#Word Width:     16
#ColMux:         8
#Bit Write:      on
#Test Mode:      off
#Created Data:   2024-3-29 10:29:186

MACRO dpram16x4096
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN dpram16x4096 0 0 ;
  SIZE 294.36 BY 326.068 ;
  SYMMETRY X Y R90 ;

  PIN AB[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 137.23 0.0 137.35 0.24 ;
      LAYER M2 ;
        RECT 137.23 0.0 137.35 0.24 ;
      LAYER M3 ;
        RECT 137.23 0.0 137.35 0.24 ;
    END
  END AB[11]
  PIN AA[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 157.01 0.0 157.13 0.24 ;
      LAYER M2 ;
        RECT 157.01 0.0 157.13 0.24 ;
      LAYER M3 ;
        RECT 157.01 0.0 157.13 0.24 ;
    END
  END AA[11]
  PIN AB[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 136.789 0.0 136.909 0.24 ;
      LAYER M2 ;
        RECT 136.789 0.0 136.909 0.24 ;
      LAYER M3 ;
        RECT 136.789 0.0 136.909 0.24 ;
    END
  END AB[10]
  PIN AA[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 157.451 0.0 157.571 0.24 ;
      LAYER M2 ;
        RECT 157.451 0.0 157.571 0.24 ;
      LAYER M3 ;
        RECT 157.451 0.0 157.571 0.24 ;
    END
  END AA[10]
  PIN AB[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 136.35 0.0 136.47 0.24 ;
      LAYER M2 ;
        RECT 136.35 0.0 136.47 0.24 ;
      LAYER M3 ;
        RECT 136.35 0.0 136.47 0.24 ;
    END
  END AB[9]
  PIN AA[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 157.89 0.0 158.01 0.24 ;
      LAYER M2 ;
        RECT 157.89 0.0 158.01 0.24 ;
      LAYER M3 ;
        RECT 157.89 0.0 158.01 0.24 ;
    END
  END AA[9]
  PIN AB[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 135.43 0.0 135.55 0.24 ;
      LAYER M2 ;
        RECT 135.43 0.0 135.55 0.24 ;
      LAYER M3 ;
        RECT 135.43 0.0 135.55 0.24 ;
    END
  END AB[8]
  PIN AA[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 158.81 0.0 158.93 0.24 ;
      LAYER M2 ;
        RECT 158.81 0.0 158.93 0.24 ;
      LAYER M3 ;
        RECT 158.81 0.0 158.93 0.24 ;
    END
  END AA[8]
  PIN AB[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 133.98 0.0 134.1 0.24 ;
      LAYER M2 ;
        RECT 133.98 0.0 134.1 0.24 ;
      LAYER M3 ;
        RECT 133.98 0.0 134.1 0.24 ;
    END
  END AB[7]
  PIN AA[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 160.26 0.0 160.38 0.24 ;
      LAYER M2 ;
        RECT 160.26 0.0 160.38 0.24 ;
      LAYER M3 ;
        RECT 160.26 0.0 160.38 0.24 ;
    END
  END AA[7]
  PIN AB[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 133.03 0.0 133.15 0.24 ;
      LAYER M2 ;
        RECT 133.03 0.0 133.15 0.24 ;
      LAYER M3 ;
        RECT 133.03 0.0 133.15 0.24 ;
    END
  END AB[6]
  PIN AA[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 161.21 0.0 161.33 0.24 ;
      LAYER M2 ;
        RECT 161.21 0.0 161.33 0.24 ;
      LAYER M3 ;
        RECT 161.21 0.0 161.33 0.24 ;
    END
  END AA[6]
  PIN AB[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 131.865 0.0 131.985 0.24 ;
      LAYER M2 ;
        RECT 131.865 0.0 131.985 0.24 ;
      LAYER M3 ;
        RECT 131.865 0.0 131.985 0.24 ;
    END
  END AB[5]
  PIN AA[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 162.375 0.0 162.495 0.24 ;
      LAYER M2 ;
        RECT 162.375 0.0 162.495 0.24 ;
      LAYER M3 ;
        RECT 162.375 0.0 162.495 0.24 ;
    END
  END AA[5]
  PIN AB[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 131.515 0.0 131.635 0.24 ;
      LAYER M2 ;
        RECT 131.515 0.0 131.635 0.24 ;
      LAYER M3 ;
        RECT 131.515 0.0 131.635 0.24 ;
    END
  END AB[4]
  PIN AA[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 162.725 0.0 162.845 0.24 ;
      LAYER M2 ;
        RECT 162.725 0.0 162.845 0.24 ;
      LAYER M3 ;
        RECT 162.725 0.0 162.845 0.24 ;
    END
  END AA[4]
  PIN AB[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 130.35 0.0 130.47 0.24 ;
      LAYER M2 ;
        RECT 130.35 0.0 130.47 0.24 ;
      LAYER M3 ;
        RECT 130.35 0.0 130.47 0.24 ;
    END
  END AB[3]
  PIN AA[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 163.89 0.0 164.01 0.24 ;
      LAYER M2 ;
        RECT 163.89 0.0 164.01 0.24 ;
      LAYER M3 ;
        RECT 163.89 0.0 164.01 0.24 ;
    END
  END AA[3]
  PIN AB[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 127.95 0.0 128.07 0.24 ;
      LAYER M2 ;
        RECT 127.95 0.0 128.07 0.24 ;
      LAYER M3 ;
        RECT 127.95 0.0 128.07 0.24 ;
    END
  END AB[2]
  PIN AA[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 166.29 0.0 166.41 0.24 ;
      LAYER M2 ;
        RECT 166.29 0.0 166.41 0.24 ;
      LAYER M3 ;
        RECT 166.29 0.0 166.41 0.24 ;
    END
  END AA[2]
  PIN AB[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 128.3 0.0 128.42 0.24 ;
      LAYER M2 ;
        RECT 128.3 0.0 128.42 0.24 ;
      LAYER M3 ;
        RECT 128.3 0.0 128.42 0.24 ;
    END
  END AB[1]
  PIN AA[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 165.94 0.0 166.06 0.24 ;
      LAYER M2 ;
        RECT 165.94 0.0 166.06 0.24 ;
      LAYER M3 ;
        RECT 165.94 0.0 166.06 0.24 ;
    END
  END AA[1]
  PIN AB[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 125.74 0.0 125.86 0.24 ;
      LAYER M2 ;
        RECT 125.74 0.0 125.86 0.24 ;
      LAYER M3 ;
        RECT 125.74 0.0 125.86 0.24 ;
    END
  END AB[0]
  PIN AA[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 168.5 0.0 168.62 0.24 ;
      LAYER M2 ;
        RECT 168.5 0.0 168.62 0.24 ;
      LAYER M3 ;
        RECT 168.5 0.0 168.62 0.24 ;
    END
  END AA[0]
  PIN QB[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 10.595 0.0 10.715 0.24 ;
      LAYER M2 ;
        RECT 10.595 0.0 10.715 0.24 ;
      LAYER M3 ;
        RECT 10.595 0.0 10.715 0.24 ;
    END
  END QB[15]
  PIN DB[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 9.64 0.0 9.76 0.24 ;
      LAYER M2 ;
        RECT 9.64 0.0 9.76 0.24 ;
      LAYER M3 ;
        RECT 9.64 0.0 9.76 0.24 ;
    END
  END DB[15]
  PIN QA[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.772 0.0 6.892 0.24 ;
      LAYER M2 ;
        RECT 6.772 0.0 6.892 0.24 ;
      LAYER M3 ;
        RECT 6.772 0.0 6.892 0.24 ;
    END
  END QA[15]
  PIN DA[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 7.722 0.0 7.842 0.24 ;
      LAYER M2 ;
        RECT 7.722 0.0 7.842 0.24 ;
      LAYER M3 ;
        RECT 7.722 0.0 7.842 0.24 ;
    END
  END DA[15]
  PIN QB[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 23.005 0.0 23.125 0.24 ;
      LAYER M2 ;
        RECT 23.005 0.0 23.125 0.24 ;
      LAYER M3 ;
        RECT 23.005 0.0 23.125 0.24 ;
    END
  END QB[14]
  PIN DB[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 23.96 0.0 24.08 0.24 ;
      LAYER M2 ;
        RECT 23.96 0.0 24.08 0.24 ;
      LAYER M3 ;
        RECT 23.96 0.0 24.08 0.24 ;
    END
  END DB[14]
  PIN QA[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 26.828 0.0 26.948 0.24 ;
      LAYER M2 ;
        RECT 26.828 0.0 26.948 0.24 ;
      LAYER M3 ;
        RECT 26.828 0.0 26.948 0.24 ;
    END
  END QA[14]
  PIN DA[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 25.878 0.0 25.998 0.24 ;
      LAYER M2 ;
        RECT 25.878 0.0 25.998 0.24 ;
      LAYER M3 ;
        RECT 25.878 0.0 25.998 0.24 ;
    END
  END DA[14]
  PIN QB[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 41.155 0.0 41.275 0.24 ;
      LAYER M2 ;
        RECT 41.155 0.0 41.275 0.24 ;
      LAYER M3 ;
        RECT 41.155 0.0 41.275 0.24 ;
    END
  END QB[13]
  PIN DB[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 40.2 0.0 40.32 0.24 ;
      LAYER M2 ;
        RECT 40.2 0.0 40.32 0.24 ;
      LAYER M3 ;
        RECT 40.2 0.0 40.32 0.24 ;
    END
  END DB[13]
  PIN QA[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 37.332 0.0 37.452 0.24 ;
      LAYER M2 ;
        RECT 37.332 0.0 37.452 0.24 ;
      LAYER M3 ;
        RECT 37.332 0.0 37.452 0.24 ;
    END
  END QA[13]
  PIN DA[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 38.282 0.0 38.402 0.24 ;
      LAYER M2 ;
        RECT 38.282 0.0 38.402 0.24 ;
      LAYER M3 ;
        RECT 38.282 0.0 38.402 0.24 ;
    END
  END DA[13]
  PIN QB[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 53.565 0.0 53.685 0.24 ;
      LAYER M2 ;
        RECT 53.565 0.0 53.685 0.24 ;
      LAYER M3 ;
        RECT 53.565 0.0 53.685 0.24 ;
    END
  END QB[12]
  PIN DB[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 54.52 0.0 54.64 0.24 ;
      LAYER M2 ;
        RECT 54.52 0.0 54.64 0.24 ;
      LAYER M3 ;
        RECT 54.52 0.0 54.64 0.24 ;
    END
  END DB[12]
  PIN QA[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 57.388 0.0 57.508 0.24 ;
      LAYER M2 ;
        RECT 57.388 0.0 57.508 0.24 ;
      LAYER M3 ;
        RECT 57.388 0.0 57.508 0.24 ;
    END
  END QA[12]
  PIN DA[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 56.438 0.0 56.558 0.24 ;
      LAYER M2 ;
        RECT 56.438 0.0 56.558 0.24 ;
      LAYER M3 ;
        RECT 56.438 0.0 56.558 0.24 ;
    END
  END DA[12]
  PIN QB[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 71.715 0.0 71.835 0.24 ;
      LAYER M2 ;
        RECT 71.715 0.0 71.835 0.24 ;
      LAYER M3 ;
        RECT 71.715 0.0 71.835 0.24 ;
    END
  END QB[11]
  PIN DB[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 70.76 0.0 70.88 0.24 ;
      LAYER M2 ;
        RECT 70.76 0.0 70.88 0.24 ;
      LAYER M3 ;
        RECT 70.76 0.0 70.88 0.24 ;
    END
  END DB[11]
  PIN QA[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 67.892 0.0 68.012 0.24 ;
      LAYER M2 ;
        RECT 67.892 0.0 68.012 0.24 ;
      LAYER M3 ;
        RECT 67.892 0.0 68.012 0.24 ;
    END
  END QA[11]
  PIN DA[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 68.842 0.0 68.962 0.24 ;
      LAYER M2 ;
        RECT 68.842 0.0 68.962 0.24 ;
      LAYER M3 ;
        RECT 68.842 0.0 68.962 0.24 ;
    END
  END DA[11]
  PIN QB[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 84.125 0.0 84.245 0.24 ;
      LAYER M2 ;
        RECT 84.125 0.0 84.245 0.24 ;
      LAYER M3 ;
        RECT 84.125 0.0 84.245 0.24 ;
    END
  END QB[10]
  PIN DB[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 85.08 0.0 85.2 0.24 ;
      LAYER M2 ;
        RECT 85.08 0.0 85.2 0.24 ;
      LAYER M3 ;
        RECT 85.08 0.0 85.2 0.24 ;
    END
  END DB[10]
  PIN QA[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 87.948 0.0 88.068 0.24 ;
      LAYER M2 ;
        RECT 87.948 0.0 88.068 0.24 ;
      LAYER M3 ;
        RECT 87.948 0.0 88.068 0.24 ;
    END
  END QA[10]
  PIN DA[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 86.998 0.0 87.118 0.24 ;
      LAYER M2 ;
        RECT 86.998 0.0 87.118 0.24 ;
      LAYER M3 ;
        RECT 86.998 0.0 87.118 0.24 ;
    END
  END DA[10]
  PIN QB[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 102.275 0.0 102.395 0.24 ;
      LAYER M2 ;
        RECT 102.275 0.0 102.395 0.24 ;
      LAYER M3 ;
        RECT 102.275 0.0 102.395 0.24 ;
    END
  END QB[9]
  PIN DB[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 101.32 0.0 101.44 0.24 ;
      LAYER M2 ;
        RECT 101.32 0.0 101.44 0.24 ;
      LAYER M3 ;
        RECT 101.32 0.0 101.44 0.24 ;
    END
  END DB[9]
  PIN QA[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 98.452 0.0 98.572 0.24 ;
      LAYER M2 ;
        RECT 98.452 0.0 98.572 0.24 ;
      LAYER M3 ;
        RECT 98.452 0.0 98.572 0.24 ;
    END
  END QA[9]
  PIN DA[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 99.402 0.0 99.522 0.24 ;
      LAYER M2 ;
        RECT 99.402 0.0 99.522 0.24 ;
      LAYER M3 ;
        RECT 99.402 0.0 99.522 0.24 ;
    END
  END DA[9]
  PIN QB[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 114.685 0.0 114.805 0.24 ;
      LAYER M2 ;
        RECT 114.685 0.0 114.805 0.24 ;
      LAYER M3 ;
        RECT 114.685 0.0 114.805 0.24 ;
    END
  END QB[8]
  PIN DB[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 115.64 0.0 115.76 0.24 ;
      LAYER M2 ;
        RECT 115.64 0.0 115.76 0.24 ;
      LAYER M3 ;
        RECT 115.64 0.0 115.76 0.24 ;
    END
  END DB[8]
  PIN QA[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 118.508 0.0 118.628 0.24 ;
      LAYER M2 ;
        RECT 118.508 0.0 118.628 0.24 ;
      LAYER M3 ;
        RECT 118.508 0.0 118.628 0.24 ;
    END
  END QA[8]
  PIN DA[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 117.558 0.0 117.678 0.24 ;
      LAYER M2 ;
        RECT 117.558 0.0 117.678 0.24 ;
      LAYER M3 ;
        RECT 117.558 0.0 117.678 0.24 ;
    END
  END DA[8]
  PIN QB[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 179.555 0.0 179.675 0.24 ;
      LAYER M2 ;
        RECT 179.555 0.0 179.675 0.24 ;
      LAYER M3 ;
        RECT 179.555 0.0 179.675 0.24 ;
    END
  END QB[7]
  PIN DB[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 178.6 0.0 178.72 0.24 ;
      LAYER M2 ;
        RECT 178.6 0.0 178.72 0.24 ;
      LAYER M3 ;
        RECT 178.6 0.0 178.72 0.24 ;
    END
  END DB[7]
  PIN QA[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 175.732 0.0 175.852 0.24 ;
      LAYER M2 ;
        RECT 175.732 0.0 175.852 0.24 ;
      LAYER M3 ;
        RECT 175.732 0.0 175.852 0.24 ;
    END
  END QA[7]
  PIN DA[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 176.682 0.0 176.802 0.24 ;
      LAYER M2 ;
        RECT 176.682 0.0 176.802 0.24 ;
      LAYER M3 ;
        RECT 176.682 0.0 176.802 0.24 ;
    END
  END DA[7]
  PIN QB[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 191.965 0.0 192.085 0.24 ;
      LAYER M2 ;
        RECT 191.965 0.0 192.085 0.24 ;
      LAYER M3 ;
        RECT 191.965 0.0 192.085 0.24 ;
    END
  END QB[6]
  PIN DB[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 192.92 0.0 193.04 0.24 ;
      LAYER M2 ;
        RECT 192.92 0.0 193.04 0.24 ;
      LAYER M3 ;
        RECT 192.92 0.0 193.04 0.24 ;
    END
  END DB[6]
  PIN QA[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 195.788 0.0 195.908 0.24 ;
      LAYER M2 ;
        RECT 195.788 0.0 195.908 0.24 ;
      LAYER M3 ;
        RECT 195.788 0.0 195.908 0.24 ;
    END
  END QA[6]
  PIN DA[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 194.838 0.0 194.958 0.24 ;
      LAYER M2 ;
        RECT 194.838 0.0 194.958 0.24 ;
      LAYER M3 ;
        RECT 194.838 0.0 194.958 0.24 ;
    END
  END DA[6]
  PIN QB[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 210.115 0.0 210.235 0.24 ;
      LAYER M2 ;
        RECT 210.115 0.0 210.235 0.24 ;
      LAYER M3 ;
        RECT 210.115 0.0 210.235 0.24 ;
    END
  END QB[5]
  PIN DB[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 209.16 0.0 209.28 0.24 ;
      LAYER M2 ;
        RECT 209.16 0.0 209.28 0.24 ;
      LAYER M3 ;
        RECT 209.16 0.0 209.28 0.24 ;
    END
  END DB[5]
  PIN QA[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 206.292 0.0 206.412 0.24 ;
      LAYER M2 ;
        RECT 206.292 0.0 206.412 0.24 ;
      LAYER M3 ;
        RECT 206.292 0.0 206.412 0.24 ;
    END
  END QA[5]
  PIN DA[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 207.242 0.0 207.362 0.24 ;
      LAYER M2 ;
        RECT 207.242 0.0 207.362 0.24 ;
      LAYER M3 ;
        RECT 207.242 0.0 207.362 0.24 ;
    END
  END DA[5]
  PIN QB[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 222.525 0.0 222.645 0.24 ;
      LAYER M2 ;
        RECT 222.525 0.0 222.645 0.24 ;
      LAYER M3 ;
        RECT 222.525 0.0 222.645 0.24 ;
    END
  END QB[4]
  PIN DB[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 223.48 0.0 223.6 0.24 ;
      LAYER M2 ;
        RECT 223.48 0.0 223.6 0.24 ;
      LAYER M3 ;
        RECT 223.48 0.0 223.6 0.24 ;
    END
  END DB[4]
  PIN QA[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 226.348 0.0 226.468 0.24 ;
      LAYER M2 ;
        RECT 226.348 0.0 226.468 0.24 ;
      LAYER M3 ;
        RECT 226.348 0.0 226.468 0.24 ;
    END
  END QA[4]
  PIN DA[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 225.398 0.0 225.518 0.24 ;
      LAYER M2 ;
        RECT 225.398 0.0 225.518 0.24 ;
      LAYER M3 ;
        RECT 225.398 0.0 225.518 0.24 ;
    END
  END DA[4]
  PIN QB[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 240.675 0.0 240.795 0.24 ;
      LAYER M2 ;
        RECT 240.675 0.0 240.795 0.24 ;
      LAYER M3 ;
        RECT 240.675 0.0 240.795 0.24 ;
    END
  END QB[3]
  PIN DB[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 239.72 0.0 239.84 0.24 ;
      LAYER M2 ;
        RECT 239.72 0.0 239.84 0.24 ;
      LAYER M3 ;
        RECT 239.72 0.0 239.84 0.24 ;
    END
  END DB[3]
  PIN QA[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 236.852 0.0 236.972 0.24 ;
      LAYER M2 ;
        RECT 236.852 0.0 236.972 0.24 ;
      LAYER M3 ;
        RECT 236.852 0.0 236.972 0.24 ;
    END
  END QA[3]
  PIN DA[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 237.802 0.0 237.922 0.24 ;
      LAYER M2 ;
        RECT 237.802 0.0 237.922 0.24 ;
      LAYER M3 ;
        RECT 237.802 0.0 237.922 0.24 ;
    END
  END DA[3]
  PIN QB[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 253.085 0.0 253.205 0.24 ;
      LAYER M2 ;
        RECT 253.085 0.0 253.205 0.24 ;
      LAYER M3 ;
        RECT 253.085 0.0 253.205 0.24 ;
    END
  END QB[2]
  PIN DB[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 254.04 0.0 254.16 0.24 ;
      LAYER M2 ;
        RECT 254.04 0.0 254.16 0.24 ;
      LAYER M3 ;
        RECT 254.04 0.0 254.16 0.24 ;
    END
  END DB[2]
  PIN QA[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 256.908 0.0 257.028 0.24 ;
      LAYER M2 ;
        RECT 256.908 0.0 257.028 0.24 ;
      LAYER M3 ;
        RECT 256.908 0.0 257.028 0.24 ;
    END
  END QA[2]
  PIN DA[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 255.958 0.0 256.078 0.24 ;
      LAYER M2 ;
        RECT 255.958 0.0 256.078 0.24 ;
      LAYER M3 ;
        RECT 255.958 0.0 256.078 0.24 ;
    END
  END DA[2]
  PIN QB[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 271.235 0.0 271.355 0.24 ;
      LAYER M2 ;
        RECT 271.235 0.0 271.355 0.24 ;
      LAYER M3 ;
        RECT 271.235 0.0 271.355 0.24 ;
    END
  END QB[1]
  PIN DB[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 270.28 0.0 270.4 0.24 ;
      LAYER M2 ;
        RECT 270.28 0.0 270.4 0.24 ;
      LAYER M3 ;
        RECT 270.28 0.0 270.4 0.24 ;
    END
  END DB[1]
  PIN QA[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 267.412 0.0 267.532 0.24 ;
      LAYER M2 ;
        RECT 267.412 0.0 267.532 0.24 ;
      LAYER M3 ;
        RECT 267.412 0.0 267.532 0.24 ;
    END
  END QA[1]
  PIN DA[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 268.362 0.0 268.482 0.24 ;
      LAYER M2 ;
        RECT 268.362 0.0 268.482 0.24 ;
      LAYER M3 ;
        RECT 268.362 0.0 268.482 0.24 ;
    END
  END DA[1]
  PIN QB[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 283.645 0.0 283.765 0.24 ;
      LAYER M2 ;
        RECT 283.645 0.0 283.765 0.24 ;
      LAYER M3 ;
        RECT 283.645 0.0 283.765 0.24 ;
    END
  END QB[0]
  PIN DB[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 284.6 0.0 284.72 0.24 ;
      LAYER M2 ;
        RECT 284.6 0.0 284.72 0.24 ;
      LAYER M3 ;
        RECT 284.6 0.0 284.72 0.24 ;
    END
  END DB[0]
  PIN QA[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 287.468 0.0 287.588 0.24 ;
      LAYER M2 ;
        RECT 287.468 0.0 287.588 0.24 ;
      LAYER M3 ;
        RECT 287.468 0.0 287.588 0.24 ;
    END
  END QA[0]
  PIN DA[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 286.518 0.0 286.638 0.24 ;
      LAYER M2 ;
        RECT 286.518 0.0 286.638 0.24 ;
      LAYER M3 ;
        RECT 286.518 0.0 286.638 0.24 ;
    END
  END DA[0]
  PIN BWENB[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 11.545 0.0 11.665 0.24 ;
      LAYER M2 ;
        RECT 11.545 0.0 11.665 0.24 ;
      LAYER M3 ;
        RECT 11.545 0.0 11.665 0.24 ;
    END
  END BWENB[15]
  PIN BWENA[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.817 0.0 5.937 0.24 ;
      LAYER M2 ;
        RECT 5.817 0.0 5.937 0.24 ;
      LAYER M3 ;
        RECT 5.817 0.0 5.937 0.24 ;
    END
  END BWENA[15]
  PIN BWENB[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 22.055 0.0 22.175 0.24 ;
      LAYER M2 ;
        RECT 22.055 0.0 22.175 0.24 ;
      LAYER M3 ;
        RECT 22.055 0.0 22.175 0.24 ;
    END
  END BWENB[14]
  PIN BWENA[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 27.783 0.0 27.903 0.24 ;
      LAYER M2 ;
        RECT 27.783 0.0 27.903 0.24 ;
      LAYER M3 ;
        RECT 27.783 0.0 27.903 0.24 ;
    END
  END BWENA[14]
  PIN BWENB[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 42.105 0.0 42.225 0.24 ;
      LAYER M2 ;
        RECT 42.105 0.0 42.225 0.24 ;
      LAYER M3 ;
        RECT 42.105 0.0 42.225 0.24 ;
    END
  END BWENB[13]
  PIN BWENA[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 36.377 0.0 36.497 0.24 ;
      LAYER M2 ;
        RECT 36.377 0.0 36.497 0.24 ;
      LAYER M3 ;
        RECT 36.377 0.0 36.497 0.24 ;
    END
  END BWENA[13]
  PIN BWENB[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 52.615 0.0 52.735 0.24 ;
      LAYER M2 ;
        RECT 52.615 0.0 52.735 0.24 ;
      LAYER M3 ;
        RECT 52.615 0.0 52.735 0.24 ;
    END
  END BWENB[12]
  PIN BWENA[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 58.343 0.0 58.463 0.24 ;
      LAYER M2 ;
        RECT 58.343 0.0 58.463 0.24 ;
      LAYER M3 ;
        RECT 58.343 0.0 58.463 0.24 ;
    END
  END BWENA[12]
  PIN BWENB[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 72.665 0.0 72.785 0.24 ;
      LAYER M2 ;
        RECT 72.665 0.0 72.785 0.24 ;
      LAYER M3 ;
        RECT 72.665 0.0 72.785 0.24 ;
    END
  END BWENB[11]
  PIN BWENA[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 66.937 0.0 67.057 0.24 ;
      LAYER M2 ;
        RECT 66.937 0.0 67.057 0.24 ;
      LAYER M3 ;
        RECT 66.937 0.0 67.057 0.24 ;
    END
  END BWENA[11]
  PIN BWENB[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 83.175 0.0 83.295 0.24 ;
      LAYER M2 ;
        RECT 83.175 0.0 83.295 0.24 ;
      LAYER M3 ;
        RECT 83.175 0.0 83.295 0.24 ;
    END
  END BWENB[10]
  PIN BWENA[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 88.903 0.0 89.023 0.24 ;
      LAYER M2 ;
        RECT 88.903 0.0 89.023 0.24 ;
      LAYER M3 ;
        RECT 88.903 0.0 89.023 0.24 ;
    END
  END BWENA[10]
  PIN BWENB[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 103.225 0.0 103.345 0.24 ;
      LAYER M2 ;
        RECT 103.225 0.0 103.345 0.24 ;
      LAYER M3 ;
        RECT 103.225 0.0 103.345 0.24 ;
    END
  END BWENB[9]
  PIN BWENA[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 97.497 0.0 97.617 0.24 ;
      LAYER M2 ;
        RECT 97.497 0.0 97.617 0.24 ;
      LAYER M3 ;
        RECT 97.497 0.0 97.617 0.24 ;
    END
  END BWENA[9]
  PIN BWENB[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 113.735 0.0 113.855 0.24 ;
      LAYER M2 ;
        RECT 113.735 0.0 113.855 0.24 ;
      LAYER M3 ;
        RECT 113.735 0.0 113.855 0.24 ;
    END
  END BWENB[8]
  PIN BWENA[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 119.463 0.0 119.583 0.24 ;
      LAYER M2 ;
        RECT 119.463 0.0 119.583 0.24 ;
      LAYER M3 ;
        RECT 119.463 0.0 119.583 0.24 ;
    END
  END BWENA[8]
  PIN BWENB[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 180.505 0.0 180.625 0.24 ;
      LAYER M2 ;
        RECT 180.505 0.0 180.625 0.24 ;
      LAYER M3 ;
        RECT 180.505 0.0 180.625 0.24 ;
    END
  END BWENB[7]
  PIN BWENA[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 174.777 0.0 174.897 0.24 ;
      LAYER M2 ;
        RECT 174.777 0.0 174.897 0.24 ;
      LAYER M3 ;
        RECT 174.777 0.0 174.897 0.24 ;
    END
  END BWENA[7]
  PIN BWENB[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 191.015 0.0 191.135 0.24 ;
      LAYER M2 ;
        RECT 191.015 0.0 191.135 0.24 ;
      LAYER M3 ;
        RECT 191.015 0.0 191.135 0.24 ;
    END
  END BWENB[6]
  PIN BWENA[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 196.743 0.0 196.863 0.24 ;
      LAYER M2 ;
        RECT 196.743 0.0 196.863 0.24 ;
      LAYER M3 ;
        RECT 196.743 0.0 196.863 0.24 ;
    END
  END BWENA[6]
  PIN BWENB[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 211.065 0.0 211.185 0.24 ;
      LAYER M2 ;
        RECT 211.065 0.0 211.185 0.24 ;
      LAYER M3 ;
        RECT 211.065 0.0 211.185 0.24 ;
    END
  END BWENB[5]
  PIN BWENA[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 205.337 0.0 205.457 0.24 ;
      LAYER M2 ;
        RECT 205.337 0.0 205.457 0.24 ;
      LAYER M3 ;
        RECT 205.337 0.0 205.457 0.24 ;
    END
  END BWENA[5]
  PIN BWENB[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 221.575 0.0 221.695 0.24 ;
      LAYER M2 ;
        RECT 221.575 0.0 221.695 0.24 ;
      LAYER M3 ;
        RECT 221.575 0.0 221.695 0.24 ;
    END
  END BWENB[4]
  PIN BWENA[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 227.303 0.0 227.423 0.24 ;
      LAYER M2 ;
        RECT 227.303 0.0 227.423 0.24 ;
      LAYER M3 ;
        RECT 227.303 0.0 227.423 0.24 ;
    END
  END BWENA[4]
  PIN BWENB[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 241.625 0.0 241.745 0.24 ;
      LAYER M2 ;
        RECT 241.625 0.0 241.745 0.24 ;
      LAYER M3 ;
        RECT 241.625 0.0 241.745 0.24 ;
    END
  END BWENB[3]
  PIN BWENA[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 235.897 0.0 236.017 0.24 ;
      LAYER M2 ;
        RECT 235.897 0.0 236.017 0.24 ;
      LAYER M3 ;
        RECT 235.897 0.0 236.017 0.24 ;
    END
  END BWENA[3]
  PIN BWENB[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 252.135 0.0 252.255 0.24 ;
      LAYER M2 ;
        RECT 252.135 0.0 252.255 0.24 ;
      LAYER M3 ;
        RECT 252.135 0.0 252.255 0.24 ;
    END
  END BWENB[2]
  PIN BWENA[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 257.863 0.0 257.983 0.24 ;
      LAYER M2 ;
        RECT 257.863 0.0 257.983 0.24 ;
      LAYER M3 ;
        RECT 257.863 0.0 257.983 0.24 ;
    END
  END BWENA[2]
  PIN BWENB[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 272.185 0.0 272.305 0.24 ;
      LAYER M2 ;
        RECT 272.185 0.0 272.305 0.24 ;
      LAYER M3 ;
        RECT 272.185 0.0 272.305 0.24 ;
    END
  END BWENB[1]
  PIN BWENA[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 266.457 0.0 266.577 0.24 ;
      LAYER M2 ;
        RECT 266.457 0.0 266.577 0.24 ;
      LAYER M3 ;
        RECT 266.457 0.0 266.577 0.24 ;
    END
  END BWENA[1]
  PIN BWENB[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 282.695 0.0 282.815 0.24 ;
      LAYER M2 ;
        RECT 282.695 0.0 282.815 0.24 ;
      LAYER M3 ;
        RECT 282.695 0.0 282.815 0.24 ;
    END
  END BWENB[0]
  PIN BWENA[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 288.423 0.0 288.543 0.24 ;
      LAYER M2 ;
        RECT 288.423 0.0 288.543 0.24 ;
      LAYER M3 ;
        RECT 288.423 0.0 288.543 0.24 ;
    END
  END BWENA[0]
  PIN WENB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 139.63 0.0 139.75 0.24 ;
      LAYER M2 ;
        RECT 139.63 0.0 139.75 0.24 ;
      LAYER M3 ;
        RECT 139.63 0.0 139.75 0.24 ;
    END
  END WENB
  PIN CENB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 140.55 0.0 140.67 0.24 ;
      LAYER M2 ;
        RECT 140.55 0.0 140.67 0.24 ;
      LAYER M3 ;
        RECT 140.55 0.0 140.67 0.24 ;
    END
  END CENB
  PIN CLKB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 142.15 0.0 142.27 0.24 ;
      LAYER M2 ;
        RECT 142.15 0.0 142.27 0.24 ;
      LAYER M3 ;
        RECT 142.15 0.0 142.27 0.24 ;
    END
  END CLKB
  PIN WENA
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 154.61 0.0 154.73 0.24 ;
      LAYER M2 ;
        RECT 154.61 0.0 154.73 0.24 ;
      LAYER M3 ;
        RECT 154.61 0.0 154.73 0.24 ;
    END
  END WENA
  PIN CENA
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 153.69 0.0 153.81 0.24 ;
      LAYER M2 ;
        RECT 153.69 0.0 153.81 0.24 ;
      LAYER M3 ;
        RECT 153.69 0.0 153.81 0.24 ;
    END
  END CENA
  PIN CLKA
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 152.09 0.0 152.21 0.24 ;
      LAYER M2 ;
        RECT 152.09 0.0 152.21 0.24 ;
      LAYER M3 ;
        RECT 152.09 0.0 152.21 0.24 ;
    END
  END CLKA
  PIN VDD 
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M4 ;
        RECT 0.45 0 0.8 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 2.36 0 2.71 139.69 ;
        RECT 2.4299999999999997 139.69 2.64 190.823 ;
        RECT 2.36 190.823 2.71 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 4.27 0 4.62 139.69 ;
        RECT 4.34 139.69 4.55 190.823 ;
        RECT 4.27 190.823 4.62 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 6.18 0 6.53 139.69 ;
        RECT 6.25 139.69 6.46 190.823 ;
        RECT 6.18 190.823 6.53 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 8.09 0 8.44 139.69 ;
        RECT 8.16 139.69 8.37 190.823 ;
        RECT 8.09 190.823 8.44 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 10.0 0 10.35 139.69 ;
        RECT 10.07 139.69 10.28 190.823 ;
        RECT 10.0 190.823 10.35 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 11.91 0 12.26 139.69 ;
        RECT 11.98 139.69 12.19 190.823 ;
        RECT 11.91 190.823 12.26 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 13.82 0 14.17 139.69 ;
        RECT 13.89 139.69 14.1 190.823 ;
        RECT 13.82 190.823 14.17 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 15.73 0 16.08 139.69 ;
        RECT 15.8 139.69 16.009999999999998 190.823 ;
        RECT 15.73 190.823 16.08 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 31.01 0 31.36 139.69 ;
        RECT 31.080000000000002 139.69 31.29 190.823 ;
        RECT 31.01 190.823 31.36 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 29.1 0 29.45 139.69 ;
        RECT 29.17 139.69 29.38 190.823 ;
        RECT 29.1 190.823 29.45 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 27.19 0 27.54 139.69 ;
        RECT 27.26 139.69 27.47 190.823 ;
        RECT 27.19 190.823 27.54 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 25.28 0 25.63 139.69 ;
        RECT 25.35 139.69 25.56 190.823 ;
        RECT 25.28 190.823 25.63 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 23.37 0 23.72 139.69 ;
        RECT 23.44 139.69 23.65 190.823 ;
        RECT 23.37 190.823 23.72 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 21.46 0 21.81 139.69 ;
        RECT 21.53 139.69 21.74 190.823 ;
        RECT 21.46 190.823 21.81 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 19.55 0 19.9 139.69 ;
        RECT 19.62 139.69 19.83 190.823 ;
        RECT 19.55 190.823 19.9 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 17.64 0 17.99 139.69 ;
        RECT 17.71 139.69 17.919999999999998 190.823 ;
        RECT 17.64 190.823 17.99 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 32.92 0 33.27 139.69 ;
        RECT 32.99 139.69 33.2 190.823 ;
        RECT 32.92 190.823 33.27 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 34.83 0 35.18 139.69 ;
        RECT 34.9 139.69 35.11 190.823 ;
        RECT 34.83 190.823 35.18 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 36.74 0 37.09 139.69 ;
        RECT 36.81 139.69 37.02 190.823 ;
        RECT 36.74 190.823 37.09 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 38.65 0 39.0 139.69 ;
        RECT 38.72 139.69 38.93 190.823 ;
        RECT 38.65 190.823 39.0 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 40.56 0 40.91 139.69 ;
        RECT 40.63 139.69 40.839999999999996 190.823 ;
        RECT 40.56 190.823 40.91 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 42.47 0 42.82 139.69 ;
        RECT 42.54 139.69 42.75 190.823 ;
        RECT 42.47 190.823 42.82 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 44.38 0 44.73 139.69 ;
        RECT 44.45 139.69 44.66 190.823 ;
        RECT 44.38 190.823 44.73 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 46.29 0 46.64 139.69 ;
        RECT 46.36 139.69 46.57 190.823 ;
        RECT 46.29 190.823 46.64 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 61.57 0 61.92 139.69 ;
        RECT 61.64 139.69 61.85 190.823 ;
        RECT 61.57 190.823 61.92 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 59.66 0 60.01 139.69 ;
        RECT 59.73 139.69 59.94 190.823 ;
        RECT 59.66 190.823 60.01 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 57.75 0 58.1 139.69 ;
        RECT 57.82 139.69 58.03 190.823 ;
        RECT 57.75 190.823 58.1 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 55.84 0 56.19 139.69 ;
        RECT 55.910000000000004 139.69 56.12 190.823 ;
        RECT 55.84 190.823 56.19 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 53.93 0 54.28 139.69 ;
        RECT 54.0 139.69 54.21 190.823 ;
        RECT 53.93 190.823 54.28 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 52.02 0 52.37 139.69 ;
        RECT 52.09 139.69 52.3 190.823 ;
        RECT 52.02 190.823 52.37 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 50.11 0 50.46 139.69 ;
        RECT 50.18 139.69 50.39 190.823 ;
        RECT 50.11 190.823 50.46 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 48.2 0 48.55 139.69 ;
        RECT 48.27 139.69 48.48 190.823 ;
        RECT 48.2 190.823 48.55 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 63.48 0 63.83 139.69 ;
        RECT 63.55 139.69 63.76 190.823 ;
        RECT 63.48 190.823 63.83 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 65.39 0 65.74 139.69 ;
        RECT 65.46 139.69 65.67 190.823 ;
        RECT 65.39 190.823 65.74 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 67.3 0 67.65 139.69 ;
        RECT 67.36999999999999 139.69 67.58000000000001 190.823 ;
        RECT 67.3 190.823 67.65 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 69.21 0 69.56 139.69 ;
        RECT 69.27999999999999 139.69 69.49000000000001 190.823 ;
        RECT 69.21 190.823 69.56 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 71.12 0 71.47 139.69 ;
        RECT 71.19 139.69 71.4 190.823 ;
        RECT 71.12 190.823 71.47 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 73.03 0 73.38 139.69 ;
        RECT 73.1 139.69 73.31 190.823 ;
        RECT 73.03 190.823 73.38 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 74.94 0 75.29 139.69 ;
        RECT 75.00999999999999 139.69 75.22000000000001 190.823 ;
        RECT 74.94 190.823 75.29 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 76.85 0 77.2 139.69 ;
        RECT 76.91999999999999 139.69 77.13000000000001 190.823 ;
        RECT 76.85 190.823 77.2 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 92.13 0 92.48 139.69 ;
        RECT 92.19999999999999 139.69 92.41000000000001 190.823 ;
        RECT 92.13 190.823 92.48 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 90.22 0 90.57 139.69 ;
        RECT 90.28999999999999 139.69 90.5 190.823 ;
        RECT 90.22 190.823 90.57 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 88.31 0 88.66 139.69 ;
        RECT 88.38 139.69 88.59 190.823 ;
        RECT 88.31 190.823 88.66 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 86.4 0 86.75 139.69 ;
        RECT 86.47 139.69 86.68 190.823 ;
        RECT 86.4 190.823 86.75 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 84.49 0 84.84 139.69 ;
        RECT 84.55999999999999 139.69 84.77000000000001 190.823 ;
        RECT 84.49 190.823 84.84 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 82.58 0 82.93 139.69 ;
        RECT 82.64999999999999 139.69 82.86000000000001 190.823 ;
        RECT 82.58 190.823 82.93 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 80.67 0 81.02 139.69 ;
        RECT 80.74 139.69 80.95 190.823 ;
        RECT 80.67 190.823 81.02 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 78.76 0 79.11 139.69 ;
        RECT 78.83 139.69 79.04 190.823 ;
        RECT 78.76 190.823 79.11 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 94.04 0 94.39 139.69 ;
        RECT 94.11 139.69 94.32000000000001 190.823 ;
        RECT 94.04 190.823 94.39 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 95.95 0 96.3 139.69 ;
        RECT 96.02 139.69 96.23 190.823 ;
        RECT 95.95 190.823 96.3 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 97.86 0 98.21 139.69 ;
        RECT 97.92999999999999 139.69 98.14 190.823 ;
        RECT 97.86 190.823 98.21 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 99.77 0 100.12 139.69 ;
        RECT 99.83999999999999 139.69 100.05000000000001 190.823 ;
        RECT 99.77 190.823 100.12 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 101.68 0 102.03 139.69 ;
        RECT 101.75 139.69 101.96000000000001 190.823 ;
        RECT 101.68 190.823 102.03 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 103.59 0 103.94 139.69 ;
        RECT 103.66 139.69 103.87 190.823 ;
        RECT 103.59 190.823 103.94 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 105.5 0 105.85 139.69 ;
        RECT 105.57 139.69 105.78 190.823 ;
        RECT 105.5 190.823 105.85 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 107.41 0 107.76 139.69 ;
        RECT 107.47999999999999 139.69 107.69000000000001 190.823 ;
        RECT 107.41 190.823 107.76 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 122.69 0 123.04 139.69 ;
        RECT 122.75999999999999 139.69 122.97000000000001 190.823 ;
        RECT 122.69 190.823 123.04 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 120.78 0 121.13 139.69 ;
        RECT 120.85 139.69 121.06 190.823 ;
        RECT 120.78 190.823 121.13 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 118.87 0 119.22 139.69 ;
        RECT 118.94 139.69 119.15 190.823 ;
        RECT 118.87 190.823 119.22 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 116.96 0 117.31 139.69 ;
        RECT 117.02999999999999 139.69 117.24000000000001 190.823 ;
        RECT 116.96 190.823 117.31 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 115.05 0 115.4 139.69 ;
        RECT 115.11999999999999 139.69 115.33000000000001 190.823 ;
        RECT 115.05 190.823 115.4 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 113.14 0 113.49 139.69 ;
        RECT 113.21 139.69 113.42 190.823 ;
        RECT 113.14 190.823 113.49 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 111.23 0 111.58 139.69 ;
        RECT 111.3 139.69 111.51 190.823 ;
        RECT 111.23 190.823 111.58 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 109.32 0 109.67 139.69 ;
        RECT 109.38999999999999 139.69 109.60000000000001 190.823 ;
        RECT 109.32 190.823 109.67 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 124.6 0 124.95 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 166.61 0 167.01 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 148.61 0 149.01 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 148.01 0 148.41 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 165.41 0 165.81 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 147.41 0 147.81 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 145.35 0 145.75 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 145.95 0 146.35 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 146.55 0 146.95 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 127.35 0 127.75 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 156.41 0 156.81 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 155.81 0 156.21 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 155.21 0 155.61 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 128.55 0 128.95 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 137.55 0 137.95 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 138.15 0 138.55 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 138.75 0 139.15 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 164.21 0 164.61 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 129.75 0 130.15 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 169.41 0 169.76 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 171.32 0 171.67 139.69 ;
        RECT 171.39 139.69 171.6 190.823 ;
        RECT 171.32 190.823 171.67 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 173.23 0 173.58 139.69 ;
        RECT 173.29999999999998 139.69 173.51000000000002 190.823 ;
        RECT 173.23 190.823 173.58 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 175.14 0 175.49 139.69 ;
        RECT 175.20999999999998 139.69 175.42000000000002 190.823 ;
        RECT 175.14 190.823 175.49 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 177.05 0 177.4 139.69 ;
        RECT 177.12 139.69 177.33 190.823 ;
        RECT 177.05 190.823 177.4 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 178.96 0 179.31 139.69 ;
        RECT 179.03 139.69 179.24 190.823 ;
        RECT 178.96 190.823 179.31 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 180.87 0 181.22 139.69 ;
        RECT 180.94 139.69 181.15 190.823 ;
        RECT 180.87 190.823 181.22 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 182.78 0 183.13 139.69 ;
        RECT 182.85 139.69 183.06 190.823 ;
        RECT 182.78 190.823 183.13 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 184.69 0 185.04 139.69 ;
        RECT 184.76 139.69 184.97 190.823 ;
        RECT 184.69 190.823 185.04 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 199.97 0 200.32 139.69 ;
        RECT 200.04 139.69 200.25 190.823 ;
        RECT 199.97 190.823 200.32 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 198.06 0 198.41 139.69 ;
        RECT 198.13 139.69 198.34 190.823 ;
        RECT 198.06 190.823 198.41 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 196.15 0 196.5 139.69 ;
        RECT 196.22 139.69 196.43 190.823 ;
        RECT 196.15 190.823 196.5 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 194.24 0 194.59 139.69 ;
        RECT 194.31 139.69 194.52 190.823 ;
        RECT 194.24 190.823 194.59 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 192.33 0 192.68 139.69 ;
        RECT 192.4 139.69 192.61 190.823 ;
        RECT 192.33 190.823 192.68 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 190.42 0 190.77 139.69 ;
        RECT 190.48999999999998 139.69 190.70000000000002 190.823 ;
        RECT 190.42 190.823 190.77 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 188.51 0 188.86 139.69 ;
        RECT 188.57999999999998 139.69 188.79000000000002 190.823 ;
        RECT 188.51 190.823 188.86 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 186.6 0 186.95 139.69 ;
        RECT 186.67 139.69 186.88 190.823 ;
        RECT 186.6 190.823 186.95 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 201.88 0 202.23 139.69 ;
        RECT 201.95 139.69 202.16 190.823 ;
        RECT 201.88 190.823 202.23 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 203.79 0 204.14 139.69 ;
        RECT 203.85999999999999 139.69 204.07 190.823 ;
        RECT 203.79 190.823 204.14 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 205.7 0 206.05 139.69 ;
        RECT 205.76999999999998 139.69 205.98000000000002 190.823 ;
        RECT 205.7 190.823 206.05 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 207.61 0 207.96 139.69 ;
        RECT 207.68 139.69 207.89000000000001 190.823 ;
        RECT 207.61 190.823 207.96 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 209.52 0 209.87 139.69 ;
        RECT 209.59 139.69 209.8 190.823 ;
        RECT 209.52 190.823 209.87 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 211.43 0 211.78 139.69 ;
        RECT 211.5 139.69 211.71 190.823 ;
        RECT 211.43 190.823 211.78 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 213.34 0 213.69 139.69 ;
        RECT 213.41 139.69 213.62 190.823 ;
        RECT 213.34 190.823 213.69 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 215.25 0 215.6 139.69 ;
        RECT 215.32 139.69 215.53 190.823 ;
        RECT 215.25 190.823 215.6 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 230.53 0 230.88 139.69 ;
        RECT 230.6 139.69 230.81 190.823 ;
        RECT 230.53 190.823 230.88 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 228.62 0 228.97 139.69 ;
        RECT 228.69 139.69 228.9 190.823 ;
        RECT 228.62 190.823 228.97 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 226.71 0 227.06 139.69 ;
        RECT 226.78 139.69 226.99 190.823 ;
        RECT 226.71 190.823 227.06 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 224.8 0 225.15 139.69 ;
        RECT 224.87 139.69 225.08 190.823 ;
        RECT 224.8 190.823 225.15 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 222.89 0 223.24 139.69 ;
        RECT 222.95999999999998 139.69 223.17000000000002 190.823 ;
        RECT 222.89 190.823 223.24 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 220.98 0 221.33 139.69 ;
        RECT 221.04999999999998 139.69 221.26000000000002 190.823 ;
        RECT 220.98 190.823 221.33 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 219.07 0 219.42 139.69 ;
        RECT 219.14 139.69 219.35 190.823 ;
        RECT 219.07 190.823 219.42 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 217.16 0 217.51 139.69 ;
        RECT 217.23 139.69 217.44 190.823 ;
        RECT 217.16 190.823 217.51 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 232.44 0 232.79 139.69 ;
        RECT 232.51 139.69 232.72 190.823 ;
        RECT 232.44 190.823 232.79 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 234.35 0 234.7 139.69 ;
        RECT 234.42 139.69 234.63 190.823 ;
        RECT 234.35 190.823 234.7 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 236.26 0 236.61 139.69 ;
        RECT 236.32999999999998 139.69 236.54000000000002 190.823 ;
        RECT 236.26 190.823 236.61 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 238.17 0 238.52 139.69 ;
        RECT 238.23999999999998 139.69 238.45000000000002 190.823 ;
        RECT 238.17 190.823 238.52 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 240.08 0 240.43 139.69 ;
        RECT 240.15 139.69 240.36 190.823 ;
        RECT 240.08 190.823 240.43 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 241.99 0 242.34 139.69 ;
        RECT 242.06 139.69 242.27 190.823 ;
        RECT 241.99 190.823 242.34 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 243.9 0 244.25 139.69 ;
        RECT 243.97 139.69 244.18 190.823 ;
        RECT 243.9 190.823 244.25 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 245.81 0 246.16 139.69 ;
        RECT 245.88 139.69 246.09 190.823 ;
        RECT 245.81 190.823 246.16 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 261.09 0 261.44 139.69 ;
        RECT 261.15999999999997 139.69 261.37 190.823 ;
        RECT 261.09 190.823 261.44 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 259.18 0 259.53 139.69 ;
        RECT 259.25 139.69 259.46 190.823 ;
        RECT 259.18 190.823 259.53 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 257.27 0 257.62 139.69 ;
        RECT 257.34 139.69 257.55 190.823 ;
        RECT 257.27 190.823 257.62 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 255.36 0 255.71 139.69 ;
        RECT 255.43 139.69 255.64000000000001 190.823 ;
        RECT 255.36 190.823 255.71 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 253.45 0 253.8 139.69 ;
        RECT 253.51999999999998 139.69 253.73000000000002 190.823 ;
        RECT 253.45 190.823 253.8 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 251.54 0 251.89 139.69 ;
        RECT 251.60999999999999 139.69 251.82 190.823 ;
        RECT 251.54 190.823 251.89 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 249.63 0 249.98 139.69 ;
        RECT 249.7 139.69 249.91 190.823 ;
        RECT 249.63 190.823 249.98 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 247.72 0 248.07 139.69 ;
        RECT 247.79 139.69 248.0 190.823 ;
        RECT 247.72 190.823 248.07 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 263.0 0 263.35 139.69 ;
        RECT 263.07 139.69 263.28000000000003 190.823 ;
        RECT 263.0 190.823 263.35 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 264.91 0 265.26 139.69 ;
        RECT 264.98 139.69 265.19 190.823 ;
        RECT 264.91 190.823 265.26 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 266.82 0 267.17 139.69 ;
        RECT 266.89 139.69 267.1 190.823 ;
        RECT 266.82 190.823 267.17 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 268.73 0 269.08 139.69 ;
        RECT 268.8 139.69 269.01 190.823 ;
        RECT 268.73 190.823 269.08 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 270.64 0 270.99 139.69 ;
        RECT 270.71 139.69 270.92 190.823 ;
        RECT 270.64 190.823 270.99 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 272.55 0 272.9 139.69 ;
        RECT 272.62 139.69 272.83 190.823 ;
        RECT 272.55 190.823 272.9 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 274.46 0 274.81 139.69 ;
        RECT 274.53 139.69 274.74 190.823 ;
        RECT 274.46 190.823 274.81 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 276.37 0 276.72 139.69 ;
        RECT 276.44 139.69 276.65000000000003 190.823 ;
        RECT 276.37 190.823 276.72 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 291.65 0 292.0 139.69 ;
        RECT 291.71999999999997 139.69 291.93 190.823 ;
        RECT 291.65 190.823 292.0 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 289.74 0 290.09 139.69 ;
        RECT 289.81 139.69 290.02 190.823 ;
        RECT 289.74 190.823 290.09 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 287.83 0 288.18 139.69 ;
        RECT 287.9 139.69 288.11 190.823 ;
        RECT 287.83 190.823 288.18 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 285.92 0 286.27 139.69 ;
        RECT 285.99 139.69 286.2 190.823 ;
        RECT 285.92 190.823 286.27 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 284.01 0 284.36 139.69 ;
        RECT 284.08 139.69 284.29 190.823 ;
        RECT 284.01 190.823 284.36 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 282.1 0 282.45 139.69 ;
        RECT 282.17 139.69 282.38 190.823 ;
        RECT 282.1 190.823 282.45 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 280.19 0 280.54 139.69 ;
        RECT 280.26 139.69 280.47 190.823 ;
        RECT 280.19 190.823 280.54 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 278.28 0 278.63 139.69 ;
        RECT 278.34999999999997 139.69 278.56 190.823 ;
        RECT 278.28 190.823 278.63 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 293.56 0 293.91 326.068 ;
    END 
  END VDD 
  PIN VSS 
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M4 ;
        RECT 1.405 0 1.755 139.69 ;
        RECT 1.475 139.69 1.6849999999999998 190.823 ;
        RECT 1.405 190.823 1.755 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 3.315 0 3.665 139.69 ;
        RECT 3.385 139.69 3.595 190.823 ;
        RECT 3.315 190.823 3.665 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 5.225 0 5.575 139.69 ;
        RECT 5.295 139.69 5.505 190.823 ;
        RECT 5.225 190.823 5.575 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 5.225 0 5.575 139.69 ;
        RECT 5.295 139.69 5.505 190.823 ;
        RECT 5.225 190.823 5.575 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 7.135 0 7.485 139.69 ;
        RECT 7.205 139.69 7.415 190.823 ;
        RECT 7.135 190.823 7.485 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 9.045 0 9.395 139.69 ;
        RECT 9.115 139.69 9.325 190.823 ;
        RECT 9.045 190.823 9.395 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 9.045 0 9.395 139.69 ;
        RECT 9.115 139.69 9.325 190.823 ;
        RECT 9.045 190.823 9.395 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 10.955 0 11.305 139.69 ;
        RECT 11.025 139.69 11.235 190.823 ;
        RECT 10.955 190.823 11.305 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 12.865 0 13.215 139.69 ;
        RECT 12.935 139.69 13.145 190.823 ;
        RECT 12.865 190.823 13.215 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 12.865 0 13.215 139.69 ;
        RECT 12.935 139.69 13.145 190.823 ;
        RECT 12.865 190.823 13.215 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 14.775 0 15.125 139.69 ;
        RECT 14.845 139.69 15.055 190.823 ;
        RECT 14.775 190.823 15.125 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 16.685 0 17.035 139.69 ;
        RECT 16.755 139.69 16.965 190.823 ;
        RECT 16.685 190.823 17.035 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 31.965 0 32.315 139.69 ;
        RECT 32.035 139.69 32.245 190.823 ;
        RECT 31.965 190.823 32.315 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 30.055 0 30.405 139.69 ;
        RECT 30.125 139.69 30.335 190.823 ;
        RECT 30.055 190.823 30.405 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 28.145 0 28.495 139.69 ;
        RECT 28.215 139.69 28.425 190.823 ;
        RECT 28.145 190.823 28.495 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 28.145 0 28.495 139.69 ;
        RECT 28.215 139.69 28.425 190.823 ;
        RECT 28.145 190.823 28.495 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 26.235 0 26.585 139.69 ;
        RECT 26.305 139.69 26.515 190.823 ;
        RECT 26.235 190.823 26.585 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 24.325 0 24.675 139.69 ;
        RECT 24.395 139.69 24.605 190.823 ;
        RECT 24.325 190.823 24.675 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 24.325 0 24.675 139.69 ;
        RECT 24.395 139.69 24.605 190.823 ;
        RECT 24.325 190.823 24.675 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 22.415 0 22.765 139.69 ;
        RECT 22.485 139.69 22.695 190.823 ;
        RECT 22.415 190.823 22.765 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 20.505 0 20.855 139.69 ;
        RECT 20.575 139.69 20.785 190.823 ;
        RECT 20.505 190.823 20.855 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 20.505 0 20.855 139.69 ;
        RECT 20.575 139.69 20.785 190.823 ;
        RECT 20.505 190.823 20.855 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 18.595 0 18.945 139.69 ;
        RECT 18.665 139.69 18.875 190.823 ;
        RECT 18.595 190.823 18.945 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 16.685 0 17.035 139.69 ;
        RECT 16.755 139.69 16.965 190.823 ;
        RECT 16.685 190.823 17.035 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 31.965 0 32.315 139.69 ;
        RECT 32.035 139.69 32.245 190.823 ;
        RECT 31.965 190.823 32.315 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 33.875 0 34.225 139.69 ;
        RECT 33.945 139.69 34.155 190.823 ;
        RECT 33.875 190.823 34.225 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 35.785 0 36.135 139.69 ;
        RECT 35.855 139.69 36.065 190.823 ;
        RECT 35.785 190.823 36.135 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 35.785 0 36.135 139.69 ;
        RECT 35.855 139.69 36.065 190.823 ;
        RECT 35.785 190.823 36.135 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 37.695 0 38.045 139.69 ;
        RECT 37.765 139.69 37.975 190.823 ;
        RECT 37.695 190.823 38.045 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 39.605 0 39.955 139.69 ;
        RECT 39.675 139.69 39.885 190.823 ;
        RECT 39.605 190.823 39.955 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 39.605 0 39.955 139.69 ;
        RECT 39.675 139.69 39.885 190.823 ;
        RECT 39.605 190.823 39.955 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 41.515 0 41.865 139.69 ;
        RECT 41.585 139.69 41.795 190.823 ;
        RECT 41.515 190.823 41.865 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 43.425 0 43.775 139.69 ;
        RECT 43.495 139.69 43.705 190.823 ;
        RECT 43.425 190.823 43.775 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 43.425 0 43.775 139.69 ;
        RECT 43.495 139.69 43.705 190.823 ;
        RECT 43.425 190.823 43.775 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 45.335 0 45.685 139.69 ;
        RECT 45.405 139.69 45.615 190.823 ;
        RECT 45.335 190.823 45.685 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 47.245 0 47.595 139.69 ;
        RECT 47.315 139.69 47.525 190.823 ;
        RECT 47.245 190.823 47.595 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 62.525 0 62.875 139.69 ;
        RECT 62.595 139.69 62.805 190.823 ;
        RECT 62.525 190.823 62.875 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 60.615 0 60.965 139.69 ;
        RECT 60.685 139.69 60.895 190.823 ;
        RECT 60.615 190.823 60.965 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 58.705 0 59.055 139.69 ;
        RECT 58.775 139.69 58.985 190.823 ;
        RECT 58.705 190.823 59.055 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 58.705 0 59.055 139.69 ;
        RECT 58.775 139.69 58.985 190.823 ;
        RECT 58.705 190.823 59.055 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 56.795 0 57.145 139.69 ;
        RECT 56.865 139.69 57.075 190.823 ;
        RECT 56.795 190.823 57.145 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 54.885 0 55.235 139.69 ;
        RECT 54.955 139.69 55.165 190.823 ;
        RECT 54.885 190.823 55.235 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 54.885 0 55.235 139.69 ;
        RECT 54.955 139.69 55.165 190.823 ;
        RECT 54.885 190.823 55.235 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 52.975 0 53.325 139.69 ;
        RECT 53.045 139.69 53.255 190.823 ;
        RECT 52.975 190.823 53.325 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 51.065 0 51.415 139.69 ;
        RECT 51.135 139.69 51.345 190.823 ;
        RECT 51.065 190.823 51.415 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 51.065 0 51.415 139.69 ;
        RECT 51.135 139.69 51.345 190.823 ;
        RECT 51.065 190.823 51.415 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 49.155 0 49.505 139.69 ;
        RECT 49.225 139.69 49.435 190.823 ;
        RECT 49.155 190.823 49.505 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 47.245 0 47.595 139.69 ;
        RECT 47.315 139.69 47.525 190.823 ;
        RECT 47.245 190.823 47.595 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 62.525 0 62.875 139.69 ;
        RECT 62.595 139.69 62.805 190.823 ;
        RECT 62.525 190.823 62.875 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 64.435 0 64.785 139.69 ;
        RECT 64.505 139.69 64.715 190.823 ;
        RECT 64.435 190.823 64.785 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 66.345 0 66.695 139.69 ;
        RECT 66.41499999999999 139.69 66.625 190.823 ;
        RECT 66.345 190.823 66.695 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 66.345 0 66.695 139.69 ;
        RECT 66.41499999999999 139.69 66.625 190.823 ;
        RECT 66.345 190.823 66.695 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 68.255 0 68.605 139.69 ;
        RECT 68.32499999999999 139.69 68.53500000000001 190.823 ;
        RECT 68.255 190.823 68.605 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 70.165 0 70.515 139.69 ;
        RECT 70.235 139.69 70.44500000000001 190.823 ;
        RECT 70.165 190.823 70.515 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 70.165 0 70.515 139.69 ;
        RECT 70.235 139.69 70.44500000000001 190.823 ;
        RECT 70.165 190.823 70.515 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 72.075 0 72.425 139.69 ;
        RECT 72.145 139.69 72.355 190.823 ;
        RECT 72.075 190.823 72.425 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 73.985 0 74.335 139.69 ;
        RECT 74.05499999999999 139.69 74.265 190.823 ;
        RECT 73.985 190.823 74.335 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 73.985 0 74.335 139.69 ;
        RECT 74.05499999999999 139.69 74.265 190.823 ;
        RECT 73.985 190.823 74.335 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 75.895 0 76.245 139.69 ;
        RECT 75.96499999999999 139.69 76.17500000000001 190.823 ;
        RECT 75.895 190.823 76.245 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 77.805 0 78.155 139.69 ;
        RECT 77.875 139.69 78.08500000000001 190.823 ;
        RECT 77.805 190.823 78.155 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 93.085 0 93.435 139.69 ;
        RECT 93.15499999999999 139.69 93.36500000000001 190.823 ;
        RECT 93.085 190.823 93.435 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 91.175 0 91.525 139.69 ;
        RECT 91.24499999999999 139.69 91.45500000000001 190.823 ;
        RECT 91.175 190.823 91.525 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 89.265 0 89.615 139.69 ;
        RECT 89.335 139.69 89.545 190.823 ;
        RECT 89.265 190.823 89.615 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 89.265 0 89.615 139.69 ;
        RECT 89.335 139.69 89.545 190.823 ;
        RECT 89.265 190.823 89.615 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 87.355 0 87.705 139.69 ;
        RECT 87.425 139.69 87.635 190.823 ;
        RECT 87.355 190.823 87.705 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 85.445 0 85.795 139.69 ;
        RECT 85.51499999999999 139.69 85.72500000000001 190.823 ;
        RECT 85.445 190.823 85.795 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 85.445 0 85.795 139.69 ;
        RECT 85.51499999999999 139.69 85.72500000000001 190.823 ;
        RECT 85.445 190.823 85.795 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 83.535 0 83.885 139.69 ;
        RECT 83.60499999999999 139.69 83.81500000000001 190.823 ;
        RECT 83.535 190.823 83.885 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 81.625 0 81.975 139.69 ;
        RECT 81.695 139.69 81.905 190.823 ;
        RECT 81.625 190.823 81.975 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 81.625 0 81.975 139.69 ;
        RECT 81.695 139.69 81.905 190.823 ;
        RECT 81.625 190.823 81.975 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 79.715 0 80.065 139.69 ;
        RECT 79.785 139.69 79.995 190.823 ;
        RECT 79.715 190.823 80.065 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 77.805 0 78.155 139.69 ;
        RECT 77.875 139.69 78.08500000000001 190.823 ;
        RECT 77.805 190.823 78.155 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 93.085 0 93.435 139.69 ;
        RECT 93.15499999999999 139.69 93.36500000000001 190.823 ;
        RECT 93.085 190.823 93.435 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 94.995 0 95.345 139.69 ;
        RECT 95.065 139.69 95.275 190.823 ;
        RECT 94.995 190.823 95.345 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 96.905 0 97.255 139.69 ;
        RECT 96.975 139.69 97.185 190.823 ;
        RECT 96.905 190.823 97.255 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 96.905 0 97.255 139.69 ;
        RECT 96.975 139.69 97.185 190.823 ;
        RECT 96.905 190.823 97.255 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 98.815 0 99.165 139.69 ;
        RECT 98.88499999999999 139.69 99.09500000000001 190.823 ;
        RECT 98.815 190.823 99.165 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 100.725 0 101.075 139.69 ;
        RECT 100.79499999999999 139.69 101.00500000000001 190.823 ;
        RECT 100.725 190.823 101.075 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 100.725 0 101.075 139.69 ;
        RECT 100.79499999999999 139.69 101.00500000000001 190.823 ;
        RECT 100.725 190.823 101.075 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 102.635 0 102.985 139.69 ;
        RECT 102.705 139.69 102.915 190.823 ;
        RECT 102.635 190.823 102.985 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 104.545 0 104.895 139.69 ;
        RECT 104.615 139.69 104.825 190.823 ;
        RECT 104.545 190.823 104.895 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 104.545 0 104.895 139.69 ;
        RECT 104.615 139.69 104.825 190.823 ;
        RECT 104.545 190.823 104.895 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 106.455 0 106.805 139.69 ;
        RECT 106.52499999999999 139.69 106.73500000000001 190.823 ;
        RECT 106.455 190.823 106.805 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 108.365 0 108.715 139.69 ;
        RECT 108.43499999999999 139.69 108.64500000000001 190.823 ;
        RECT 108.365 190.823 108.715 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 123.645 0 123.995 139.69 ;
        RECT 123.71499999999999 139.69 123.92500000000001 190.823 ;
        RECT 123.645 190.823 123.995 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 121.735 0 122.085 139.69 ;
        RECT 121.80499999999999 139.69 122.015 190.823 ;
        RECT 121.735 190.823 122.085 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 119.825 0 120.175 139.69 ;
        RECT 119.895 139.69 120.105 190.823 ;
        RECT 119.825 190.823 120.175 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 119.825 0 120.175 139.69 ;
        RECT 119.895 139.69 120.105 190.823 ;
        RECT 119.825 190.823 120.175 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 117.915 0 118.265 139.69 ;
        RECT 117.985 139.69 118.19500000000001 190.823 ;
        RECT 117.915 190.823 118.265 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 116.005 0 116.355 139.69 ;
        RECT 116.07499999999999 139.69 116.28500000000001 190.823 ;
        RECT 116.005 190.823 116.355 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 116.005 0 116.355 139.69 ;
        RECT 116.07499999999999 139.69 116.28500000000001 190.823 ;
        RECT 116.005 190.823 116.355 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 114.095 0 114.445 139.69 ;
        RECT 114.16499999999999 139.69 114.375 190.823 ;
        RECT 114.095 190.823 114.445 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 112.185 0 112.535 139.69 ;
        RECT 112.255 139.69 112.465 190.823 ;
        RECT 112.185 190.823 112.535 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 112.185 0 112.535 139.69 ;
        RECT 112.255 139.69 112.465 190.823 ;
        RECT 112.185 190.823 112.535 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 110.275 0 110.625 139.69 ;
        RECT 110.345 139.69 110.555 190.823 ;
        RECT 110.275 190.823 110.625 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 108.365 0 108.715 139.69 ;
        RECT 108.43499999999999 139.69 108.64500000000001 190.823 ;
        RECT 108.365 190.823 108.715 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 167.21 0 167.61 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 126.75 0 127.15 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 126.15 0 126.55 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 167.81 0 168.21 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 152.81 0 153.21 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 149.81 0 150.21 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 154.01 0 154.41 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 139.95 0 140.35 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 141.15 0 141.55 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 158.21 0 158.61 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 159.41 0 159.81 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 160.61 0 161.01 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 161.81 0 162.21 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 163.01 0 163.41 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 144.15 0 144.55 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 142.95 0 143.35 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 135.75 0 136.15 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 134.55 0 134.95 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 133.35 0 133.75 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 132.15 0 132.55 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 130.95 0 131.35 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 151.01 0 151.41 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 170.365 0 170.715 139.69 ;
        RECT 170.435 139.69 170.645 190.823 ;
        RECT 170.365 190.823 170.715 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 172.275 0 172.625 139.69 ;
        RECT 172.345 139.69 172.555 190.823 ;
        RECT 172.275 190.823 172.625 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 174.185 0 174.535 139.69 ;
        RECT 174.255 139.69 174.465 190.823 ;
        RECT 174.185 190.823 174.535 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 174.185 0 174.535 139.69 ;
        RECT 174.255 139.69 174.465 190.823 ;
        RECT 174.185 190.823 174.535 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 176.095 0 176.445 139.69 ;
        RECT 176.165 139.69 176.375 190.823 ;
        RECT 176.095 190.823 176.445 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 178.005 0 178.355 139.69 ;
        RECT 178.075 139.69 178.285 190.823 ;
        RECT 178.005 190.823 178.355 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 178.005 0 178.355 139.69 ;
        RECT 178.075 139.69 178.285 190.823 ;
        RECT 178.005 190.823 178.355 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 179.915 0 180.265 139.69 ;
        RECT 179.98499999999999 139.69 180.195 190.823 ;
        RECT 179.915 190.823 180.265 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 181.825 0 182.175 139.69 ;
        RECT 181.89499999999998 139.69 182.10500000000002 190.823 ;
        RECT 181.825 190.823 182.175 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 181.825 0 182.175 139.69 ;
        RECT 181.89499999999998 139.69 182.10500000000002 190.823 ;
        RECT 181.825 190.823 182.175 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 183.735 0 184.085 139.69 ;
        RECT 183.805 139.69 184.01500000000001 190.823 ;
        RECT 183.735 190.823 184.085 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 185.645 0 185.995 139.69 ;
        RECT 185.715 139.69 185.925 190.823 ;
        RECT 185.645 190.823 185.995 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 200.925 0 201.275 139.69 ;
        RECT 200.995 139.69 201.205 190.823 ;
        RECT 200.925 190.823 201.275 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 199.015 0 199.365 139.69 ;
        RECT 199.08499999999998 139.69 199.29500000000002 190.823 ;
        RECT 199.015 190.823 199.365 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 197.105 0 197.455 139.69 ;
        RECT 197.17499999999998 139.69 197.38500000000002 190.823 ;
        RECT 197.105 190.823 197.455 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 197.105 0 197.455 139.69 ;
        RECT 197.17499999999998 139.69 197.38500000000002 190.823 ;
        RECT 197.105 190.823 197.455 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 195.195 0 195.545 139.69 ;
        RECT 195.265 139.69 195.475 190.823 ;
        RECT 195.195 190.823 195.545 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 193.285 0 193.635 139.69 ;
        RECT 193.355 139.69 193.565 190.823 ;
        RECT 193.285 190.823 193.635 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 193.285 0 193.635 139.69 ;
        RECT 193.355 139.69 193.565 190.823 ;
        RECT 193.285 190.823 193.635 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 191.375 0 191.725 139.69 ;
        RECT 191.445 139.69 191.655 190.823 ;
        RECT 191.375 190.823 191.725 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 189.465 0 189.815 139.69 ;
        RECT 189.535 139.69 189.745 190.823 ;
        RECT 189.465 190.823 189.815 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 189.465 0 189.815 139.69 ;
        RECT 189.535 139.69 189.745 190.823 ;
        RECT 189.465 190.823 189.815 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 187.555 0 187.905 139.69 ;
        RECT 187.625 139.69 187.835 190.823 ;
        RECT 187.555 190.823 187.905 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 185.645 0 185.995 139.69 ;
        RECT 185.715 139.69 185.925 190.823 ;
        RECT 185.645 190.823 185.995 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 200.925 0 201.275 139.69 ;
        RECT 200.995 139.69 201.205 190.823 ;
        RECT 200.925 190.823 201.275 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 202.835 0 203.185 139.69 ;
        RECT 202.905 139.69 203.115 190.823 ;
        RECT 202.835 190.823 203.185 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 204.745 0 205.095 139.69 ;
        RECT 204.815 139.69 205.025 190.823 ;
        RECT 204.745 190.823 205.095 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 204.745 0 205.095 139.69 ;
        RECT 204.815 139.69 205.025 190.823 ;
        RECT 204.745 190.823 205.095 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 206.655 0 207.005 139.69 ;
        RECT 206.725 139.69 206.935 190.823 ;
        RECT 206.655 190.823 207.005 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 208.565 0 208.915 139.69 ;
        RECT 208.635 139.69 208.845 190.823 ;
        RECT 208.565 190.823 208.915 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 208.565 0 208.915 139.69 ;
        RECT 208.635 139.69 208.845 190.823 ;
        RECT 208.565 190.823 208.915 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 210.475 0 210.825 139.69 ;
        RECT 210.545 139.69 210.755 190.823 ;
        RECT 210.475 190.823 210.825 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 212.385 0 212.735 139.69 ;
        RECT 212.45499999999998 139.69 212.66500000000002 190.823 ;
        RECT 212.385 190.823 212.735 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 212.385 0 212.735 139.69 ;
        RECT 212.45499999999998 139.69 212.66500000000002 190.823 ;
        RECT 212.385 190.823 212.735 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 214.295 0 214.645 139.69 ;
        RECT 214.36499999999998 139.69 214.57500000000002 190.823 ;
        RECT 214.295 190.823 214.645 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 216.205 0 216.555 139.69 ;
        RECT 216.275 139.69 216.485 190.823 ;
        RECT 216.205 190.823 216.555 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 231.485 0 231.835 139.69 ;
        RECT 231.555 139.69 231.76500000000001 190.823 ;
        RECT 231.485 190.823 231.835 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 229.575 0 229.925 139.69 ;
        RECT 229.64499999999998 139.69 229.85500000000002 190.823 ;
        RECT 229.575 190.823 229.925 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 227.665 0 228.015 139.69 ;
        RECT 227.73499999999999 139.69 227.945 190.823 ;
        RECT 227.665 190.823 228.015 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 227.665 0 228.015 139.69 ;
        RECT 227.73499999999999 139.69 227.945 190.823 ;
        RECT 227.665 190.823 228.015 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 225.755 0 226.105 139.69 ;
        RECT 225.825 139.69 226.035 190.823 ;
        RECT 225.755 190.823 226.105 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 223.845 0 224.195 139.69 ;
        RECT 223.915 139.69 224.125 190.823 ;
        RECT 223.845 190.823 224.195 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 223.845 0 224.195 139.69 ;
        RECT 223.915 139.69 224.125 190.823 ;
        RECT 223.845 190.823 224.195 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 221.935 0 222.285 139.69 ;
        RECT 222.005 139.69 222.215 190.823 ;
        RECT 221.935 190.823 222.285 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 220.025 0 220.375 139.69 ;
        RECT 220.095 139.69 220.305 190.823 ;
        RECT 220.025 190.823 220.375 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 220.025 0 220.375 139.69 ;
        RECT 220.095 139.69 220.305 190.823 ;
        RECT 220.025 190.823 220.375 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 218.115 0 218.465 139.69 ;
        RECT 218.185 139.69 218.395 190.823 ;
        RECT 218.115 190.823 218.465 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 216.205 0 216.555 139.69 ;
        RECT 216.275 139.69 216.485 190.823 ;
        RECT 216.205 190.823 216.555 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 231.485 0 231.835 139.69 ;
        RECT 231.555 139.69 231.76500000000001 190.823 ;
        RECT 231.485 190.823 231.835 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 233.395 0 233.745 139.69 ;
        RECT 233.465 139.69 233.675 190.823 ;
        RECT 233.395 190.823 233.745 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 235.305 0 235.655 139.69 ;
        RECT 235.375 139.69 235.585 190.823 ;
        RECT 235.305 190.823 235.655 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 235.305 0 235.655 139.69 ;
        RECT 235.375 139.69 235.585 190.823 ;
        RECT 235.305 190.823 235.655 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 237.215 0 237.565 139.69 ;
        RECT 237.285 139.69 237.495 190.823 ;
        RECT 237.215 190.823 237.565 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 239.125 0 239.475 139.69 ;
        RECT 239.195 139.69 239.405 190.823 ;
        RECT 239.125 190.823 239.475 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 239.125 0 239.475 139.69 ;
        RECT 239.195 139.69 239.405 190.823 ;
        RECT 239.125 190.823 239.475 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 241.035 0 241.385 139.69 ;
        RECT 241.105 139.69 241.315 190.823 ;
        RECT 241.035 190.823 241.385 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 242.945 0 243.295 139.69 ;
        RECT 243.015 139.69 243.225 190.823 ;
        RECT 242.945 190.823 243.295 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 242.945 0 243.295 139.69 ;
        RECT 243.015 139.69 243.225 190.823 ;
        RECT 242.945 190.823 243.295 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 244.855 0 245.205 139.69 ;
        RECT 244.92499999999998 139.69 245.13500000000002 190.823 ;
        RECT 244.855 190.823 245.205 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 246.765 0 247.115 139.69 ;
        RECT 246.83499999999998 139.69 247.04500000000002 190.823 ;
        RECT 246.765 190.823 247.115 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 262.045 0 262.395 139.69 ;
        RECT 262.115 139.69 262.325 190.823 ;
        RECT 262.045 190.823 262.395 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 260.135 0 260.485 139.69 ;
        RECT 260.205 139.69 260.415 190.823 ;
        RECT 260.135 190.823 260.485 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 258.225 0 258.575 139.69 ;
        RECT 258.295 139.69 258.505 190.823 ;
        RECT 258.225 190.823 258.575 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 258.225 0 258.575 139.69 ;
        RECT 258.295 139.69 258.505 190.823 ;
        RECT 258.225 190.823 258.575 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 256.315 0 256.665 139.69 ;
        RECT 256.385 139.69 256.595 190.823 ;
        RECT 256.315 190.823 256.665 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 254.405 0 254.755 139.69 ;
        RECT 254.475 139.69 254.685 190.823 ;
        RECT 254.405 190.823 254.755 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 254.405 0 254.755 139.69 ;
        RECT 254.475 139.69 254.685 190.823 ;
        RECT 254.405 190.823 254.755 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 252.495 0 252.845 139.69 ;
        RECT 252.565 139.69 252.775 190.823 ;
        RECT 252.495 190.823 252.845 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 250.585 0 250.935 139.69 ;
        RECT 250.655 139.69 250.865 190.823 ;
        RECT 250.585 190.823 250.935 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 250.585 0 250.935 139.69 ;
        RECT 250.655 139.69 250.865 190.823 ;
        RECT 250.585 190.823 250.935 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 248.675 0 249.025 139.69 ;
        RECT 248.745 139.69 248.955 190.823 ;
        RECT 248.675 190.823 249.025 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 246.765 0 247.115 139.69 ;
        RECT 246.83499999999998 139.69 247.04500000000002 190.823 ;
        RECT 246.765 190.823 247.115 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 262.045 0 262.395 139.69 ;
        RECT 262.115 139.69 262.325 190.823 ;
        RECT 262.045 190.823 262.395 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 263.955 0 264.305 139.69 ;
        RECT 264.025 139.69 264.235 190.823 ;
        RECT 263.955 190.823 264.305 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 265.865 0 266.215 139.69 ;
        RECT 265.935 139.69 266.145 190.823 ;
        RECT 265.865 190.823 266.215 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 265.865 0 266.215 139.69 ;
        RECT 265.935 139.69 266.145 190.823 ;
        RECT 265.865 190.823 266.215 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 267.775 0 268.125 139.69 ;
        RECT 267.84499999999997 139.69 268.055 190.823 ;
        RECT 267.775 190.823 268.125 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 269.685 0 270.035 139.69 ;
        RECT 269.755 139.69 269.96500000000003 190.823 ;
        RECT 269.685 190.823 270.035 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 269.685 0 270.035 139.69 ;
        RECT 269.755 139.69 269.96500000000003 190.823 ;
        RECT 269.685 190.823 270.035 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 271.595 0 271.945 139.69 ;
        RECT 271.665 139.69 271.875 190.823 ;
        RECT 271.595 190.823 271.945 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 273.505 0 273.855 139.69 ;
        RECT 273.575 139.69 273.785 190.823 ;
        RECT 273.505 190.823 273.855 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 273.505 0 273.855 139.69 ;
        RECT 273.575 139.69 273.785 190.823 ;
        RECT 273.505 190.823 273.855 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 275.415 0 275.765 139.69 ;
        RECT 275.485 139.69 275.695 190.823 ;
        RECT 275.415 190.823 275.765 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 277.325 0 277.675 139.69 ;
        RECT 277.395 139.69 277.605 190.823 ;
        RECT 277.325 190.823 277.675 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 292.605 0 292.955 139.69 ;
        RECT 292.675 139.69 292.885 190.823 ;
        RECT 292.605 190.823 292.955 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 290.695 0 291.045 139.69 ;
        RECT 290.765 139.69 290.975 190.823 ;
        RECT 290.695 190.823 291.045 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 288.785 0 289.135 139.69 ;
        RECT 288.855 139.69 289.065 190.823 ;
        RECT 288.785 190.823 289.135 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 288.785 0 289.135 139.69 ;
        RECT 288.855 139.69 289.065 190.823 ;
        RECT 288.785 190.823 289.135 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 286.875 0 287.225 139.69 ;
        RECT 286.945 139.69 287.15500000000003 190.823 ;
        RECT 286.875 190.823 287.225 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 284.965 0 285.315 139.69 ;
        RECT 285.03499999999997 139.69 285.245 190.823 ;
        RECT 284.965 190.823 285.315 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 284.965 0 285.315 139.69 ;
        RECT 285.03499999999997 139.69 285.245 190.823 ;
        RECT 284.965 190.823 285.315 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 283.055 0 283.405 139.69 ;
        RECT 283.125 139.69 283.335 190.823 ;
        RECT 283.055 190.823 283.405 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 281.145 0 281.495 139.69 ;
        RECT 281.215 139.69 281.425 190.823 ;
        RECT 281.145 190.823 281.495 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 281.145 0 281.495 139.69 ;
        RECT 281.215 139.69 281.425 190.823 ;
        RECT 281.145 190.823 281.495 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 279.235 0 279.585 139.69 ;
        RECT 279.305 139.69 279.515 190.823 ;
        RECT 279.235 190.823 279.585 326.068 ;
    END 
    PORT
      LAYER M4 ;
        RECT 277.325 0 277.675 139.69 ;
        RECT 277.395 139.69 277.605 190.823 ;
        RECT 277.325 190.823 277.675 326.068 ;
    END 
  END VSS 
  OBS
    LAYER M1 SPACING 0.1 ;
      RECT  0.00 0.33999999999999997 294.36 326.068 ;
      RECT 0.0 0.0 5.7170000000000005 0.33999999999999997 ;
      RECT 6.037 0.0 6.672000000000001 0.33999999999999997 ;
      RECT 6.992 0.0 7.622000000000001 0.33999999999999997 ;
      RECT 7.941999999999999 0.0 9.540000000000001 0.33999999999999997 ;
      RECT 9.86 0.0 10.495000000000001 0.33999999999999997 ;
      RECT 10.815 0.0 11.445 0.33999999999999997 ;
      RECT 11.764999999999999 0.0 21.955 0.33999999999999997 ;
      RECT 22.275000000000002 0.0 22.904999999999998 0.33999999999999997 ;
      RECT 23.225 0.0 23.86 0.33999999999999997 ;
      RECT 24.18 0.0 25.778 0.33999999999999997 ;
      RECT 26.098000000000003 0.0 26.727999999999998 0.33999999999999997 ;
      RECT 27.048000000000002 0.0 27.683 0.33999999999999997 ;
      RECT 28.003 0.0 36.277 0.33999999999999997 ;
      RECT 36.597 0.0 37.232 0.33999999999999997 ;
      RECT 37.552 0.0 38.181999999999995 0.33999999999999997 ;
      RECT 38.502 0.0 40.1 0.33999999999999997 ;
      RECT 40.42 0.0 41.055 0.33999999999999997 ;
      RECT 41.375 0.0 42.004999999999995 0.33999999999999997 ;
      RECT 42.325 0.0 52.515 0.33999999999999997 ;
      RECT 52.835 0.0 53.464999999999996 0.33999999999999997 ;
      RECT 53.785000000000004 0.0 54.42 0.33999999999999997 ;
      RECT 54.74 0.0 56.338 0.33999999999999997 ;
      RECT 56.658 0.0 57.288 0.33999999999999997 ;
      RECT 57.608000000000004 0.0 58.243 0.33999999999999997 ;
      RECT 58.563 0.0 66.837 0.33999999999999997 ;
      RECT 67.157 0.0 67.792 0.33999999999999997 ;
      RECT 68.112 0.0 68.742 0.33999999999999997 ;
      RECT 69.062 0.0 70.66000000000001 0.33999999999999997 ;
      RECT 70.97999999999999 0.0 71.61500000000001 0.33999999999999997 ;
      RECT 71.93499999999999 0.0 72.56500000000001 0.33999999999999997 ;
      RECT 72.88499999999999 0.0 83.075 0.33999999999999997 ;
      RECT 83.395 0.0 84.025 0.33999999999999997 ;
      RECT 84.345 0.0 84.98 0.33999999999999997 ;
      RECT 85.3 0.0 86.89800000000001 0.33999999999999997 ;
      RECT 87.21799999999999 0.0 87.848 0.33999999999999997 ;
      RECT 88.16799999999999 0.0 88.80300000000001 0.33999999999999997 ;
      RECT 89.12299999999999 0.0 97.397 0.33999999999999997 ;
      RECT 97.717 0.0 98.352 0.33999999999999997 ;
      RECT 98.672 0.0 99.302 0.33999999999999997 ;
      RECT 99.622 0.0 101.22 0.33999999999999997 ;
      RECT 101.53999999999999 0.0 102.17500000000001 0.33999999999999997 ;
      RECT 102.49499999999999 0.0 103.125 0.33999999999999997 ;
      RECT 103.445 0.0 113.635 0.33999999999999997 ;
      RECT 113.955 0.0 114.58500000000001 0.33999999999999997 ;
      RECT 114.905 0.0 115.54 0.33999999999999997 ;
      RECT 115.86 0.0 117.45800000000001 0.33999999999999997 ;
      RECT 117.77799999999999 0.0 118.408 0.33999999999999997 ;
      RECT 118.728 0.0 119.363 0.33999999999999997 ;
      RECT 119.68299999999999 0.0 125.64 0.33999999999999997 ;
      RECT 125.96 0.0 127.85000000000001 0.33999999999999997 ;
      RECT 128.17 0.0 128.20000000000002 0.33999999999999997 ;
      RECT 128.51999999999998 0.0 130.25 0.33999999999999997 ;
      RECT 130.57 0.0 131.415 0.33999999999999997 ;
      RECT 131.73499999999999 0.0 131.76500000000001 0.33999999999999997 ;
      RECT 132.085 0.0 132.93 0.33999999999999997 ;
      RECT 133.25 0.0 133.88 0.33999999999999997 ;
      RECT 134.2 0.0 135.33 0.33999999999999997 ;
      RECT 135.65 0.0 136.25 0.33999999999999997 ;
      RECT 136.57 0.0 136.689 0.33999999999999997 ;
      RECT 137.009 0.0 137.13 0.33999999999999997 ;
      RECT 137.45 0.0 139.53 0.33999999999999997 ;
      RECT 139.85 0.0 140.45000000000002 0.33999999999999997 ;
      RECT 140.76999999999998 0.0 142.05 0.33999999999999997 ;
      RECT 142.37 0.0 151.99 0.33999999999999997 ;
      RECT 152.31 0.0 153.59 0.33999999999999997 ;
      RECT 153.91 0.0 154.51000000000002 0.33999999999999997 ;
      RECT 154.82999999999998 0.0 156.91 0.33999999999999997 ;
      RECT 157.23 0.0 157.351 0.33999999999999997 ;
      RECT 157.671 0.0 157.79 0.33999999999999997 ;
      RECT 158.10999999999999 0.0 158.71 0.33999999999999997 ;
      RECT 159.03 0.0 160.16 0.33999999999999997 ;
      RECT 160.48 0.0 161.11 0.33999999999999997 ;
      RECT 161.43 0.0 162.275 0.33999999999999997 ;
      RECT 162.595 0.0 162.625 0.33999999999999997 ;
      RECT 162.945 0.0 163.79 0.33999999999999997 ;
      RECT 164.10999999999999 0.0 165.84 0.33999999999999997 ;
      RECT 166.16 0.0 166.19 0.33999999999999997 ;
      RECT 166.51 0.0 168.4 0.33999999999999997 ;
      RECT 168.72 0.0 174.677 0.33999999999999997 ;
      RECT 174.99699999999999 0.0 175.632 0.33999999999999997 ;
      RECT 175.952 0.0 176.582 0.33999999999999997 ;
      RECT 176.902 0.0 178.5 0.33999999999999997 ;
      RECT 178.82 0.0 179.455 0.33999999999999997 ;
      RECT 179.775 0.0 180.405 0.33999999999999997 ;
      RECT 180.725 0.0 190.915 0.33999999999999997 ;
      RECT 191.23499999999999 0.0 191.865 0.33999999999999997 ;
      RECT 192.185 0.0 192.82 0.33999999999999997 ;
      RECT 193.14 0.0 194.738 0.33999999999999997 ;
      RECT 195.058 0.0 195.68800000000002 0.33999999999999997 ;
      RECT 196.00799999999998 0.0 196.643 0.33999999999999997 ;
      RECT 196.963 0.0 205.237 0.33999999999999997 ;
      RECT 205.557 0.0 206.192 0.33999999999999997 ;
      RECT 206.512 0.0 207.142 0.33999999999999997 ;
      RECT 207.462 0.0 209.06 0.33999999999999997 ;
      RECT 209.38 0.0 210.01500000000001 0.33999999999999997 ;
      RECT 210.335 0.0 210.965 0.33999999999999997 ;
      RECT 211.285 0.0 221.475 0.33999999999999997 ;
      RECT 221.795 0.0 222.425 0.33999999999999997 ;
      RECT 222.745 0.0 223.38 0.33999999999999997 ;
      RECT 223.7 0.0 225.298 0.33999999999999997 ;
      RECT 225.618 0.0 226.24800000000002 0.33999999999999997 ;
      RECT 226.56799999999998 0.0 227.203 0.33999999999999997 ;
      RECT 227.523 0.0 235.797 0.33999999999999997 ;
      RECT 236.117 0.0 236.752 0.33999999999999997 ;
      RECT 237.072 0.0 237.702 0.33999999999999997 ;
      RECT 238.022 0.0 239.62 0.33999999999999997 ;
      RECT 239.94 0.0 240.57500000000002 0.33999999999999997 ;
      RECT 240.89499999999998 0.0 241.525 0.33999999999999997 ;
      RECT 241.845 0.0 252.035 0.33999999999999997 ;
      RECT 252.355 0.0 252.985 0.33999999999999997 ;
      RECT 253.305 0.0 253.94 0.33999999999999997 ;
      RECT 254.26 0.0 255.858 0.33999999999999997 ;
      RECT 256.178 0.0 256.808 0.33999999999999997 ;
      RECT 257.12800000000004 0.0 257.763 0.33999999999999997 ;
      RECT 258.083 0.0 266.35699999999997 0.33999999999999997 ;
      RECT 266.677 0.0 267.31199999999995 0.33999999999999997 ;
      RECT 267.632 0.0 268.262 0.33999999999999997 ;
      RECT 268.58200000000005 0.0 270.17999999999995 0.33999999999999997 ;
      RECT 270.5 0.0 271.135 0.33999999999999997 ;
      RECT 271.45500000000004 0.0 272.085 0.33999999999999997 ;
      RECT 272.40500000000003 0.0 282.59499999999997 0.33999999999999997 ;
      RECT 282.915 0.0 283.54499999999996 0.33999999999999997 ;
      RECT 283.865 0.0 284.5 0.33999999999999997 ;
      RECT 284.82000000000005 0.0 286.41799999999995 0.33999999999999997 ;
      RECT 286.738 0.0 287.368 0.33999999999999997 ;
      RECT 287.68800000000005 0.0 288.323 0.33999999999999997 ;
      RECT 288.64300000000003 0.0 294.36 0.33999999999999997 ;
    LAYER M2 SPACING 0.1 ;
      RECT  0.00 0.33999999999999997 294.36 326.068 ;
      RECT 0.0 0.0 5.7170000000000005 0.33999999999999997 ;
      RECT 6.037 0.0 6.672000000000001 0.33999999999999997 ;
      RECT 6.992 0.0 7.622000000000001 0.33999999999999997 ;
      RECT 7.941999999999999 0.0 9.540000000000001 0.33999999999999997 ;
      RECT 9.86 0.0 10.495000000000001 0.33999999999999997 ;
      RECT 10.815 0.0 11.445 0.33999999999999997 ;
      RECT 11.764999999999999 0.0 21.955 0.33999999999999997 ;
      RECT 22.275000000000002 0.0 22.904999999999998 0.33999999999999997 ;
      RECT 23.225 0.0 23.86 0.33999999999999997 ;
      RECT 24.18 0.0 25.778 0.33999999999999997 ;
      RECT 26.098000000000003 0.0 26.727999999999998 0.33999999999999997 ;
      RECT 27.048000000000002 0.0 27.683 0.33999999999999997 ;
      RECT 28.003 0.0 36.277 0.33999999999999997 ;
      RECT 36.597 0.0 37.232 0.33999999999999997 ;
      RECT 37.552 0.0 38.181999999999995 0.33999999999999997 ;
      RECT 38.502 0.0 40.1 0.33999999999999997 ;
      RECT 40.42 0.0 41.055 0.33999999999999997 ;
      RECT 41.375 0.0 42.004999999999995 0.33999999999999997 ;
      RECT 42.325 0.0 52.515 0.33999999999999997 ;
      RECT 52.835 0.0 53.464999999999996 0.33999999999999997 ;
      RECT 53.785000000000004 0.0 54.42 0.33999999999999997 ;
      RECT 54.74 0.0 56.338 0.33999999999999997 ;
      RECT 56.658 0.0 57.288 0.33999999999999997 ;
      RECT 57.608000000000004 0.0 58.243 0.33999999999999997 ;
      RECT 58.563 0.0 66.837 0.33999999999999997 ;
      RECT 67.157 0.0 67.792 0.33999999999999997 ;
      RECT 68.112 0.0 68.742 0.33999999999999997 ;
      RECT 69.062 0.0 70.66000000000001 0.33999999999999997 ;
      RECT 70.97999999999999 0.0 71.61500000000001 0.33999999999999997 ;
      RECT 71.93499999999999 0.0 72.56500000000001 0.33999999999999997 ;
      RECT 72.88499999999999 0.0 83.075 0.33999999999999997 ;
      RECT 83.395 0.0 84.025 0.33999999999999997 ;
      RECT 84.345 0.0 84.98 0.33999999999999997 ;
      RECT 85.3 0.0 86.89800000000001 0.33999999999999997 ;
      RECT 87.21799999999999 0.0 87.848 0.33999999999999997 ;
      RECT 88.16799999999999 0.0 88.80300000000001 0.33999999999999997 ;
      RECT 89.12299999999999 0.0 97.397 0.33999999999999997 ;
      RECT 97.717 0.0 98.352 0.33999999999999997 ;
      RECT 98.672 0.0 99.302 0.33999999999999997 ;
      RECT 99.622 0.0 101.22 0.33999999999999997 ;
      RECT 101.53999999999999 0.0 102.17500000000001 0.33999999999999997 ;
      RECT 102.49499999999999 0.0 103.125 0.33999999999999997 ;
      RECT 103.445 0.0 113.635 0.33999999999999997 ;
      RECT 113.955 0.0 114.58500000000001 0.33999999999999997 ;
      RECT 114.905 0.0 115.54 0.33999999999999997 ;
      RECT 115.86 0.0 117.45800000000001 0.33999999999999997 ;
      RECT 117.77799999999999 0.0 118.408 0.33999999999999997 ;
      RECT 118.728 0.0 119.363 0.33999999999999997 ;
      RECT 119.68299999999999 0.0 125.64 0.33999999999999997 ;
      RECT 125.96 0.0 127.85000000000001 0.33999999999999997 ;
      RECT 128.17 0.0 128.20000000000002 0.33999999999999997 ;
      RECT 128.51999999999998 0.0 130.25 0.33999999999999997 ;
      RECT 130.57 0.0 131.415 0.33999999999999997 ;
      RECT 131.73499999999999 0.0 131.76500000000001 0.33999999999999997 ;
      RECT 132.085 0.0 132.93 0.33999999999999997 ;
      RECT 133.25 0.0 133.88 0.33999999999999997 ;
      RECT 134.2 0.0 135.33 0.33999999999999997 ;
      RECT 135.65 0.0 136.25 0.33999999999999997 ;
      RECT 136.57 0.0 136.689 0.33999999999999997 ;
      RECT 137.009 0.0 137.13 0.33999999999999997 ;
      RECT 137.45 0.0 139.53 0.33999999999999997 ;
      RECT 139.85 0.0 140.45000000000002 0.33999999999999997 ;
      RECT 140.76999999999998 0.0 142.05 0.33999999999999997 ;
      RECT 142.37 0.0 151.99 0.33999999999999997 ;
      RECT 152.31 0.0 153.59 0.33999999999999997 ;
      RECT 153.91 0.0 154.51000000000002 0.33999999999999997 ;
      RECT 154.82999999999998 0.0 156.91 0.33999999999999997 ;
      RECT 157.23 0.0 157.351 0.33999999999999997 ;
      RECT 157.671 0.0 157.79 0.33999999999999997 ;
      RECT 158.10999999999999 0.0 158.71 0.33999999999999997 ;
      RECT 159.03 0.0 160.16 0.33999999999999997 ;
      RECT 160.48 0.0 161.11 0.33999999999999997 ;
      RECT 161.43 0.0 162.275 0.33999999999999997 ;
      RECT 162.595 0.0 162.625 0.33999999999999997 ;
      RECT 162.945 0.0 163.79 0.33999999999999997 ;
      RECT 164.10999999999999 0.0 165.84 0.33999999999999997 ;
      RECT 166.16 0.0 166.19 0.33999999999999997 ;
      RECT 166.51 0.0 168.4 0.33999999999999997 ;
      RECT 168.72 0.0 174.677 0.33999999999999997 ;
      RECT 174.99699999999999 0.0 175.632 0.33999999999999997 ;
      RECT 175.952 0.0 176.582 0.33999999999999997 ;
      RECT 176.902 0.0 178.5 0.33999999999999997 ;
      RECT 178.82 0.0 179.455 0.33999999999999997 ;
      RECT 179.775 0.0 180.405 0.33999999999999997 ;
      RECT 180.725 0.0 190.915 0.33999999999999997 ;
      RECT 191.23499999999999 0.0 191.865 0.33999999999999997 ;
      RECT 192.185 0.0 192.82 0.33999999999999997 ;
      RECT 193.14 0.0 194.738 0.33999999999999997 ;
      RECT 195.058 0.0 195.68800000000002 0.33999999999999997 ;
      RECT 196.00799999999998 0.0 196.643 0.33999999999999997 ;
      RECT 196.963 0.0 205.237 0.33999999999999997 ;
      RECT 205.557 0.0 206.192 0.33999999999999997 ;
      RECT 206.512 0.0 207.142 0.33999999999999997 ;
      RECT 207.462 0.0 209.06 0.33999999999999997 ;
      RECT 209.38 0.0 210.01500000000001 0.33999999999999997 ;
      RECT 210.335 0.0 210.965 0.33999999999999997 ;
      RECT 211.285 0.0 221.475 0.33999999999999997 ;
      RECT 221.795 0.0 222.425 0.33999999999999997 ;
      RECT 222.745 0.0 223.38 0.33999999999999997 ;
      RECT 223.7 0.0 225.298 0.33999999999999997 ;
      RECT 225.618 0.0 226.24800000000002 0.33999999999999997 ;
      RECT 226.56799999999998 0.0 227.203 0.33999999999999997 ;
      RECT 227.523 0.0 235.797 0.33999999999999997 ;
      RECT 236.117 0.0 236.752 0.33999999999999997 ;
      RECT 237.072 0.0 237.702 0.33999999999999997 ;
      RECT 238.022 0.0 239.62 0.33999999999999997 ;
      RECT 239.94 0.0 240.57500000000002 0.33999999999999997 ;
      RECT 240.89499999999998 0.0 241.525 0.33999999999999997 ;
      RECT 241.845 0.0 252.035 0.33999999999999997 ;
      RECT 252.355 0.0 252.985 0.33999999999999997 ;
      RECT 253.305 0.0 253.94 0.33999999999999997 ;
      RECT 254.26 0.0 255.858 0.33999999999999997 ;
      RECT 256.178 0.0 256.808 0.33999999999999997 ;
      RECT 257.12800000000004 0.0 257.763 0.33999999999999997 ;
      RECT 258.083 0.0 266.35699999999997 0.33999999999999997 ;
      RECT 266.677 0.0 267.31199999999995 0.33999999999999997 ;
      RECT 267.632 0.0 268.262 0.33999999999999997 ;
      RECT 268.58200000000005 0.0 270.17999999999995 0.33999999999999997 ;
      RECT 270.5 0.0 271.135 0.33999999999999997 ;
      RECT 271.45500000000004 0.0 272.085 0.33999999999999997 ;
      RECT 272.40500000000003 0.0 282.59499999999997 0.33999999999999997 ;
      RECT 282.915 0.0 283.54499999999996 0.33999999999999997 ;
      RECT 283.865 0.0 284.5 0.33999999999999997 ;
      RECT 284.82000000000005 0.0 286.41799999999995 0.33999999999999997 ;
      RECT 286.738 0.0 287.368 0.33999999999999997 ;
      RECT 287.68800000000005 0.0 288.323 0.33999999999999997 ;
      RECT 288.64300000000003 0.0 294.36 0.33999999999999997 ;
    LAYER M3 SPACING 0.1 ;
      RECT  0.00 0.33999999999999997 294.36 326.068 ;
      RECT 0.0 0.0 5.7170000000000005 0.33999999999999997 ;
      RECT 6.037 0.0 6.672000000000001 0.33999999999999997 ;
      RECT 6.992 0.0 7.622000000000001 0.33999999999999997 ;
      RECT 7.941999999999999 0.0 9.540000000000001 0.33999999999999997 ;
      RECT 9.86 0.0 10.495000000000001 0.33999999999999997 ;
      RECT 10.815 0.0 11.445 0.33999999999999997 ;
      RECT 11.764999999999999 0.0 21.955 0.33999999999999997 ;
      RECT 22.275000000000002 0.0 22.904999999999998 0.33999999999999997 ;
      RECT 23.225 0.0 23.86 0.33999999999999997 ;
      RECT 24.18 0.0 25.778 0.33999999999999997 ;
      RECT 26.098000000000003 0.0 26.727999999999998 0.33999999999999997 ;
      RECT 27.048000000000002 0.0 27.683 0.33999999999999997 ;
      RECT 28.003 0.0 36.277 0.33999999999999997 ;
      RECT 36.597 0.0 37.232 0.33999999999999997 ;
      RECT 37.552 0.0 38.181999999999995 0.33999999999999997 ;
      RECT 38.502 0.0 40.1 0.33999999999999997 ;
      RECT 40.42 0.0 41.055 0.33999999999999997 ;
      RECT 41.375 0.0 42.004999999999995 0.33999999999999997 ;
      RECT 42.325 0.0 52.515 0.33999999999999997 ;
      RECT 52.835 0.0 53.464999999999996 0.33999999999999997 ;
      RECT 53.785000000000004 0.0 54.42 0.33999999999999997 ;
      RECT 54.74 0.0 56.338 0.33999999999999997 ;
      RECT 56.658 0.0 57.288 0.33999999999999997 ;
      RECT 57.608000000000004 0.0 58.243 0.33999999999999997 ;
      RECT 58.563 0.0 66.837 0.33999999999999997 ;
      RECT 67.157 0.0 67.792 0.33999999999999997 ;
      RECT 68.112 0.0 68.742 0.33999999999999997 ;
      RECT 69.062 0.0 70.66000000000001 0.33999999999999997 ;
      RECT 70.97999999999999 0.0 71.61500000000001 0.33999999999999997 ;
      RECT 71.93499999999999 0.0 72.56500000000001 0.33999999999999997 ;
      RECT 72.88499999999999 0.0 83.075 0.33999999999999997 ;
      RECT 83.395 0.0 84.025 0.33999999999999997 ;
      RECT 84.345 0.0 84.98 0.33999999999999997 ;
      RECT 85.3 0.0 86.89800000000001 0.33999999999999997 ;
      RECT 87.21799999999999 0.0 87.848 0.33999999999999997 ;
      RECT 88.16799999999999 0.0 88.80300000000001 0.33999999999999997 ;
      RECT 89.12299999999999 0.0 97.397 0.33999999999999997 ;
      RECT 97.717 0.0 98.352 0.33999999999999997 ;
      RECT 98.672 0.0 99.302 0.33999999999999997 ;
      RECT 99.622 0.0 101.22 0.33999999999999997 ;
      RECT 101.53999999999999 0.0 102.17500000000001 0.33999999999999997 ;
      RECT 102.49499999999999 0.0 103.125 0.33999999999999997 ;
      RECT 103.445 0.0 113.635 0.33999999999999997 ;
      RECT 113.955 0.0 114.58500000000001 0.33999999999999997 ;
      RECT 114.905 0.0 115.54 0.33999999999999997 ;
      RECT 115.86 0.0 117.45800000000001 0.33999999999999997 ;
      RECT 117.77799999999999 0.0 118.408 0.33999999999999997 ;
      RECT 118.728 0.0 119.363 0.33999999999999997 ;
      RECT 119.68299999999999 0.0 125.64 0.33999999999999997 ;
      RECT 125.96 0.0 127.85000000000001 0.33999999999999997 ;
      RECT 128.17 0.0 128.20000000000002 0.33999999999999997 ;
      RECT 128.51999999999998 0.0 130.25 0.33999999999999997 ;
      RECT 130.57 0.0 131.415 0.33999999999999997 ;
      RECT 131.73499999999999 0.0 131.76500000000001 0.33999999999999997 ;
      RECT 132.085 0.0 132.93 0.33999999999999997 ;
      RECT 133.25 0.0 133.88 0.33999999999999997 ;
      RECT 134.2 0.0 135.33 0.33999999999999997 ;
      RECT 135.65 0.0 136.25 0.33999999999999997 ;
      RECT 136.57 0.0 136.689 0.33999999999999997 ;
      RECT 137.009 0.0 137.13 0.33999999999999997 ;
      RECT 137.45 0.0 139.53 0.33999999999999997 ;
      RECT 139.85 0.0 140.45000000000002 0.33999999999999997 ;
      RECT 140.76999999999998 0.0 142.05 0.33999999999999997 ;
      RECT 142.37 0.0 151.99 0.33999999999999997 ;
      RECT 152.31 0.0 153.59 0.33999999999999997 ;
      RECT 153.91 0.0 154.51000000000002 0.33999999999999997 ;
      RECT 154.82999999999998 0.0 156.91 0.33999999999999997 ;
      RECT 157.23 0.0 157.351 0.33999999999999997 ;
      RECT 157.671 0.0 157.79 0.33999999999999997 ;
      RECT 158.10999999999999 0.0 158.71 0.33999999999999997 ;
      RECT 159.03 0.0 160.16 0.33999999999999997 ;
      RECT 160.48 0.0 161.11 0.33999999999999997 ;
      RECT 161.43 0.0 162.275 0.33999999999999997 ;
      RECT 162.595 0.0 162.625 0.33999999999999997 ;
      RECT 162.945 0.0 163.79 0.33999999999999997 ;
      RECT 164.10999999999999 0.0 165.84 0.33999999999999997 ;
      RECT 166.16 0.0 166.19 0.33999999999999997 ;
      RECT 166.51 0.0 168.4 0.33999999999999997 ;
      RECT 168.72 0.0 174.677 0.33999999999999997 ;
      RECT 174.99699999999999 0.0 175.632 0.33999999999999997 ;
      RECT 175.952 0.0 176.582 0.33999999999999997 ;
      RECT 176.902 0.0 178.5 0.33999999999999997 ;
      RECT 178.82 0.0 179.455 0.33999999999999997 ;
      RECT 179.775 0.0 180.405 0.33999999999999997 ;
      RECT 180.725 0.0 190.915 0.33999999999999997 ;
      RECT 191.23499999999999 0.0 191.865 0.33999999999999997 ;
      RECT 192.185 0.0 192.82 0.33999999999999997 ;
      RECT 193.14 0.0 194.738 0.33999999999999997 ;
      RECT 195.058 0.0 195.68800000000002 0.33999999999999997 ;
      RECT 196.00799999999998 0.0 196.643 0.33999999999999997 ;
      RECT 196.963 0.0 205.237 0.33999999999999997 ;
      RECT 205.557 0.0 206.192 0.33999999999999997 ;
      RECT 206.512 0.0 207.142 0.33999999999999997 ;
      RECT 207.462 0.0 209.06 0.33999999999999997 ;
      RECT 209.38 0.0 210.01500000000001 0.33999999999999997 ;
      RECT 210.335 0.0 210.965 0.33999999999999997 ;
      RECT 211.285 0.0 221.475 0.33999999999999997 ;
      RECT 221.795 0.0 222.425 0.33999999999999997 ;
      RECT 222.745 0.0 223.38 0.33999999999999997 ;
      RECT 223.7 0.0 225.298 0.33999999999999997 ;
      RECT 225.618 0.0 226.24800000000002 0.33999999999999997 ;
      RECT 226.56799999999998 0.0 227.203 0.33999999999999997 ;
      RECT 227.523 0.0 235.797 0.33999999999999997 ;
      RECT 236.117 0.0 236.752 0.33999999999999997 ;
      RECT 237.072 0.0 237.702 0.33999999999999997 ;
      RECT 238.022 0.0 239.62 0.33999999999999997 ;
      RECT 239.94 0.0 240.57500000000002 0.33999999999999997 ;
      RECT 240.89499999999998 0.0 241.525 0.33999999999999997 ;
      RECT 241.845 0.0 252.035 0.33999999999999997 ;
      RECT 252.355 0.0 252.985 0.33999999999999997 ;
      RECT 253.305 0.0 253.94 0.33999999999999997 ;
      RECT 254.26 0.0 255.858 0.33999999999999997 ;
      RECT 256.178 0.0 256.808 0.33999999999999997 ;
      RECT 257.12800000000004 0.0 257.763 0.33999999999999997 ;
      RECT 258.083 0.0 266.35699999999997 0.33999999999999997 ;
      RECT 266.677 0.0 267.31199999999995 0.33999999999999997 ;
      RECT 267.632 0.0 268.262 0.33999999999999997 ;
      RECT 268.58200000000005 0.0 270.17999999999995 0.33999999999999997 ;
      RECT 270.5 0.0 271.135 0.33999999999999997 ;
      RECT 271.45500000000004 0.0 272.085 0.33999999999999997 ;
      RECT 272.40500000000003 0.0 282.59499999999997 0.33999999999999997 ;
      RECT 282.915 0.0 283.54499999999996 0.33999999999999997 ;
      RECT 283.865 0.0 284.5 0.33999999999999997 ;
      RECT 284.82000000000005 0.0 286.41799999999995 0.33999999999999997 ;
      RECT 286.738 0.0 287.368 0.33999999999999997 ;
      RECT 287.68800000000005 0.0 288.323 0.33999999999999997 ;
      RECT 288.64300000000003 0.0 294.36 0.33999999999999997 ;
    LAYER M4 SPACING 0.1 ;
      RECT 2.26 139.79 2.3299999999999996 190.723 ;
      RECT 2.74 139.79 2.81 190.723 ;
      RECT 4.17 139.79 4.24 190.723 ;
      RECT 4.6499999999999995 139.79 4.72 190.723 ;
      RECT 6.08 139.79 6.15 190.723 ;
      RECT 6.56 139.79 6.63 190.723 ;
      RECT 7.99 139.79 8.06 190.723 ;
      RECT 8.469999999999999 139.79 8.54 190.723 ;
      RECT 9.9 139.79 9.97 190.723 ;
      RECT 10.379999999999999 139.79 10.45 190.723 ;
      RECT 11.81 139.79 11.88 190.723 ;
      RECT 12.29 139.79 12.36 190.723 ;
      RECT 13.72 139.79 13.790000000000001 190.723 ;
      RECT 14.2 139.79 14.27 190.723 ;
      RECT 15.63 139.79 15.700000000000001 190.723 ;
      RECT 16.11 139.79 16.18 190.723 ;
      RECT 30.91 139.79 30.98 190.723 ;
      RECT 31.39 139.79 31.46 190.723 ;
      RECT 29.0 139.79 29.07 190.723 ;
      RECT 29.48 139.79 29.55 190.723 ;
      RECT 27.09 139.79 27.16 190.723 ;
      RECT 27.57 139.79 27.64 190.723 ;
      RECT 25.18 139.79 25.25 190.723 ;
      RECT 25.66 139.79 25.73 190.723 ;
      RECT 23.27 139.79 23.34 190.723 ;
      RECT 23.75 139.79 23.82 190.723 ;
      RECT 21.36 139.79 21.43 190.723 ;
      RECT 21.84 139.79 21.91 190.723 ;
      RECT 19.45 139.79 19.52 190.723 ;
      RECT 19.93 139.79 20.0 190.723 ;
      RECT 17.54 139.79 17.61 190.723 ;
      RECT 18.02 139.79 18.09 190.723 ;
      RECT 32.82 139.79 32.89 190.723 ;
      RECT 33.300000000000004 139.79 33.370000000000005 190.723 ;
      RECT 34.73 139.79 34.8 190.723 ;
      RECT 35.21 139.79 35.28 190.723 ;
      RECT 36.64 139.79 36.71 190.723 ;
      RECT 37.120000000000005 139.79 37.190000000000005 190.723 ;
      RECT 38.55 139.79 38.62 190.723 ;
      RECT 39.03 139.79 39.1 190.723 ;
      RECT 40.46 139.79 40.53 190.723 ;
      RECT 40.94 139.79 41.01 190.723 ;
      RECT 42.37 139.79 42.44 190.723 ;
      RECT 42.85 139.79 42.92 190.723 ;
      RECT 44.28 139.79 44.35 190.723 ;
      RECT 44.76 139.79 44.83 190.723 ;
      RECT 46.19 139.79 46.26 190.723 ;
      RECT 46.67 139.79 46.74 190.723 ;
      RECT 61.47 139.79 61.54 190.723 ;
      RECT 61.95 139.79 62.02 190.723 ;
      RECT 59.559999999999995 139.79 59.629999999999995 190.723 ;
      RECT 60.04 139.79 60.11 190.723 ;
      RECT 57.65 139.79 57.72 190.723 ;
      RECT 58.13 139.79 58.2 190.723 ;
      RECT 55.74 139.79 55.81 190.723 ;
      RECT 56.22 139.79 56.29 190.723 ;
      RECT 53.83 139.79 53.9 190.723 ;
      RECT 54.31 139.79 54.38 190.723 ;
      RECT 51.92 139.79 51.99 190.723 ;
      RECT 52.4 139.79 52.47 190.723 ;
      RECT 50.01 139.79 50.08 190.723 ;
      RECT 50.49 139.79 50.56 190.723 ;
      RECT 48.1 139.79 48.17 190.723 ;
      RECT 48.58 139.79 48.65 190.723 ;
      RECT 63.379999999999995 139.79 63.449999999999996 190.723 ;
      RECT 63.86 139.79 63.93 190.723 ;
      RECT 65.29 139.79 65.36 190.723 ;
      RECT 65.77 139.79 65.83999999999999 190.723 ;
      RECT 67.2 139.79 67.27 190.723 ;
      RECT 67.68 139.79 67.75 190.723 ;
      RECT 69.11 139.79 69.17999999999999 190.723 ;
      RECT 69.59 139.79 69.66 190.723 ;
      RECT 71.02000000000001 139.79 71.09 190.723 ;
      RECT 71.5 139.79 71.57 190.723 ;
      RECT 72.93 139.79 73.0 190.723 ;
      RECT 73.41 139.79 73.47999999999999 190.723 ;
      RECT 74.84 139.79 74.91 190.723 ;
      RECT 75.32000000000001 139.79 75.39 190.723 ;
      RECT 76.75 139.79 76.82 190.723 ;
      RECT 77.23 139.79 77.3 190.723 ;
      RECT 92.03 139.79 92.1 190.723 ;
      RECT 92.51 139.79 92.58 190.723 ;
      RECT 90.12 139.79 90.19 190.723 ;
      RECT 90.6 139.79 90.66999999999999 190.723 ;
      RECT 88.21000000000001 139.79 88.28 190.723 ;
      RECT 88.69 139.79 88.75999999999999 190.723 ;
      RECT 86.30000000000001 139.79 86.37 190.723 ;
      RECT 86.78 139.79 86.85 190.723 ;
      RECT 84.39 139.79 84.46 190.723 ;
      RECT 84.87 139.79 84.94 190.723 ;
      RECT 82.48 139.79 82.55 190.723 ;
      RECT 82.96000000000001 139.79 83.03 190.723 ;
      RECT 80.57000000000001 139.79 80.64 190.723 ;
      RECT 81.05 139.79 81.11999999999999 190.723 ;
      RECT 78.66000000000001 139.79 78.73 190.723 ;
      RECT 79.14 139.79 79.21 190.723 ;
      RECT 93.94000000000001 139.79 94.01 190.723 ;
      RECT 94.42 139.79 94.49 190.723 ;
      RECT 95.85000000000001 139.79 95.92 190.723 ;
      RECT 96.33 139.79 96.39999999999999 190.723 ;
      RECT 97.76 139.79 97.83 190.723 ;
      RECT 98.24 139.79 98.30999999999999 190.723 ;
      RECT 99.67 139.79 99.74 190.723 ;
      RECT 100.15 139.79 100.22 190.723 ;
      RECT 101.58000000000001 139.79 101.65 190.723 ;
      RECT 102.06 139.79 102.13 190.723 ;
      RECT 103.49000000000001 139.79 103.56 190.723 ;
      RECT 103.97 139.79 104.03999999999999 190.723 ;
      RECT 105.4 139.79 105.47 190.723 ;
      RECT 105.88 139.79 105.94999999999999 190.723 ;
      RECT 107.31 139.79 107.38 190.723 ;
      RECT 107.79 139.79 107.86 190.723 ;
      RECT 122.59 139.79 122.66 190.723 ;
      RECT 123.07000000000001 139.79 123.14 190.723 ;
      RECT 120.68 139.79 120.75 190.723 ;
      RECT 121.16 139.79 121.22999999999999 190.723 ;
      RECT 118.77000000000001 139.79 118.84 190.723 ;
      RECT 119.25 139.79 119.32 190.723 ;
      RECT 116.86 139.79 116.92999999999999 190.723 ;
      RECT 117.34 139.79 117.41 190.723 ;
      RECT 114.95 139.79 115.02 190.723 ;
      RECT 115.43 139.79 115.5 190.723 ;
      RECT 113.04 139.79 113.11 190.723 ;
      RECT 113.52 139.79 113.58999999999999 190.723 ;
      RECT 111.13000000000001 139.79 111.2 190.723 ;
      RECT 111.61 139.79 111.67999999999999 190.723 ;
      RECT 109.22 139.79 109.28999999999999 190.723 ;
      RECT 109.7 139.79 109.77 190.723 ;
      RECT 171.22 139.79 171.29 190.723 ;
      RECT 171.7 139.79 171.76999999999998 190.723 ;
      RECT 173.13 139.79 173.2 190.723 ;
      RECT 173.61 139.79 173.68 190.723 ;
      RECT 175.04 139.79 175.10999999999999 190.723 ;
      RECT 175.52 139.79 175.59 190.723 ;
      RECT 176.95000000000002 139.79 177.02 190.723 ;
      RECT 177.43 139.79 177.5 190.723 ;
      RECT 178.86 139.79 178.93 190.723 ;
      RECT 179.34 139.79 179.41 190.723 ;
      RECT 180.77 139.79 180.84 190.723 ;
      RECT 181.25 139.79 181.32 190.723 ;
      RECT 182.68 139.79 182.75 190.723 ;
      RECT 183.16 139.79 183.23 190.723 ;
      RECT 184.59 139.79 184.66 190.723 ;
      RECT 185.07 139.79 185.14 190.723 ;
      RECT 199.87 139.79 199.94 190.723 ;
      RECT 200.35 139.79 200.42 190.723 ;
      RECT 197.96 139.79 198.03 190.723 ;
      RECT 198.44 139.79 198.51 190.723 ;
      RECT 196.05 139.79 196.12 190.723 ;
      RECT 196.53 139.79 196.6 190.723 ;
      RECT 194.14000000000001 139.79 194.21 190.723 ;
      RECT 194.62 139.79 194.69 190.723 ;
      RECT 192.23000000000002 139.79 192.3 190.723 ;
      RECT 192.71 139.79 192.78 190.723 ;
      RECT 190.32 139.79 190.39 190.723 ;
      RECT 190.8 139.79 190.87 190.723 ;
      RECT 188.41 139.79 188.48 190.723 ;
      RECT 188.89000000000001 139.79 188.96 190.723 ;
      RECT 186.5 139.79 186.57 190.723 ;
      RECT 186.98 139.79 187.04999999999998 190.723 ;
      RECT 201.78 139.79 201.85 190.723 ;
      RECT 202.26 139.79 202.32999999999998 190.723 ;
      RECT 203.69 139.79 203.76 190.723 ;
      RECT 204.17 139.79 204.23999999999998 190.723 ;
      RECT 205.6 139.79 205.67 190.723 ;
      RECT 206.08 139.79 206.15 190.723 ;
      RECT 207.51000000000002 139.79 207.58 190.723 ;
      RECT 207.99 139.79 208.06 190.723 ;
      RECT 209.42000000000002 139.79 209.49 190.723 ;
      RECT 209.9 139.79 209.97 190.723 ;
      RECT 211.33 139.79 211.4 190.723 ;
      RECT 211.81 139.79 211.88 190.723 ;
      RECT 213.24 139.79 213.31 190.723 ;
      RECT 213.72 139.79 213.79 190.723 ;
      RECT 215.15 139.79 215.22 190.723 ;
      RECT 215.63 139.79 215.7 190.723 ;
      RECT 230.43 139.79 230.5 190.723 ;
      RECT 230.91 139.79 230.98 190.723 ;
      RECT 228.52 139.79 228.59 190.723 ;
      RECT 229.0 139.79 229.07 190.723 ;
      RECT 226.61 139.79 226.68 190.723 ;
      RECT 227.09 139.79 227.16 190.723 ;
      RECT 224.70000000000002 139.79 224.77 190.723 ;
      RECT 225.18 139.79 225.25 190.723 ;
      RECT 222.79 139.79 222.85999999999999 190.723 ;
      RECT 223.27 139.79 223.34 190.723 ;
      RECT 220.88 139.79 220.95 190.723 ;
      RECT 221.36 139.79 221.43 190.723 ;
      RECT 218.97 139.79 219.04 190.723 ;
      RECT 219.45 139.79 219.51999999999998 190.723 ;
      RECT 217.06 139.79 217.13 190.723 ;
      RECT 217.54 139.79 217.60999999999999 190.723 ;
      RECT 232.34 139.79 232.41 190.723 ;
      RECT 232.82 139.79 232.89 190.723 ;
      RECT 234.25 139.79 234.32 190.723 ;
      RECT 234.73 139.79 234.79999999999998 190.723 ;
      RECT 236.16 139.79 236.23 190.723 ;
      RECT 236.64000000000001 139.79 236.71 190.723 ;
      RECT 238.07 139.79 238.14 190.723 ;
      RECT 238.55 139.79 238.62 190.723 ;
      RECT 239.98000000000002 139.79 240.05 190.723 ;
      RECT 240.46 139.79 240.53 190.723 ;
      RECT 241.89000000000001 139.79 241.96 190.723 ;
      RECT 242.37 139.79 242.44 190.723 ;
      RECT 243.8 139.79 243.87 190.723 ;
      RECT 244.28 139.79 244.35 190.723 ;
      RECT 245.71 139.79 245.78 190.723 ;
      RECT 246.19 139.79 246.26 190.723 ;
      RECT 260.98999999999995 139.79 261.05999999999995 190.723 ;
      RECT 261.47 139.79 261.54 190.723 ;
      RECT 259.08 139.79 259.15 190.723 ;
      RECT 259.56 139.79 259.63 190.723 ;
      RECT 257.16999999999996 139.79 257.23999999999995 190.723 ;
      RECT 257.65000000000003 139.79 257.72 190.723 ;
      RECT 255.26000000000002 139.79 255.33 190.723 ;
      RECT 255.74 139.79 255.81 190.723 ;
      RECT 253.35 139.79 253.42 190.723 ;
      RECT 253.83 139.79 253.9 190.723 ;
      RECT 251.44 139.79 251.51 190.723 ;
      RECT 251.92 139.79 251.98999999999998 190.723 ;
      RECT 249.53 139.79 249.6 190.723 ;
      RECT 250.01 139.79 250.07999999999998 190.723 ;
      RECT 247.62 139.79 247.69 190.723 ;
      RECT 248.1 139.79 248.17 190.723 ;
      RECT 262.9 139.79 262.96999999999997 190.723 ;
      RECT 263.38000000000005 139.79 263.45000000000005 190.723 ;
      RECT 264.81 139.79 264.88 190.723 ;
      RECT 265.29 139.79 265.36 190.723 ;
      RECT 266.71999999999997 139.79 266.78999999999996 190.723 ;
      RECT 267.20000000000005 139.79 267.27000000000004 190.723 ;
      RECT 268.63 139.79 268.7 190.723 ;
      RECT 269.11 139.79 269.18 190.723 ;
      RECT 270.53999999999996 139.79 270.60999999999996 190.723 ;
      RECT 271.02000000000004 139.79 271.09000000000003 190.723 ;
      RECT 272.45 139.79 272.52 190.723 ;
      RECT 272.93 139.79 273.0 190.723 ;
      RECT 274.35999999999996 139.79 274.42999999999995 190.723 ;
      RECT 274.84000000000003 139.79 274.91 190.723 ;
      RECT 276.27 139.79 276.34 190.723 ;
      RECT 276.75000000000006 139.79 276.82000000000005 190.723 ;
      RECT 291.54999999999995 139.79 291.61999999999995 190.723 ;
      RECT 292.03000000000003 139.79 292.1 190.723 ;
      RECT 289.64 139.79 289.71 190.723 ;
      RECT 290.12 139.79 290.19 190.723 ;
      RECT 287.72999999999996 139.79 287.79999999999995 190.723 ;
      RECT 288.21000000000004 139.79 288.28000000000003 190.723 ;
      RECT 285.82 139.79 285.89 190.723 ;
      RECT 286.3 139.79 286.37 190.723 ;
      RECT 283.90999999999997 139.79 283.97999999999996 190.723 ;
      RECT 284.39000000000004 139.79 284.46000000000004 190.723 ;
      RECT 282.0 139.79 282.07 190.723 ;
      RECT 282.48 139.79 282.55 190.723 ;
      RECT 280.09 139.79 280.15999999999997 190.723 ;
      RECT 280.57000000000005 139.79 280.64000000000004 190.723 ;
      RECT 278.17999999999995 139.79 278.24999999999994 190.723 ;
      RECT 278.66 139.79 278.73 190.723 ;
      RECT 1.305 139.79 1.375 190.723 ;
      RECT 1.785 139.79 1.855 190.723 ;
      RECT 3.215 139.79 3.2849999999999997 190.723 ;
      RECT 3.6950000000000003 139.79 3.765 190.723 ;
      RECT 5.125 139.79 5.195 190.723 ;
      RECT 5.6049999999999995 139.79 5.675 190.723 ;
      RECT 5.125 139.79 5.195 190.723 ;
      RECT 5.6049999999999995 139.79 5.675 190.723 ;
      RECT 7.035 139.79 7.105 190.723 ;
      RECT 7.515 139.79 7.585 190.723 ;
      RECT 8.945 139.79 9.015 190.723 ;
      RECT 9.424999999999999 139.79 9.495 190.723 ;
      RECT 8.945 139.79 9.015 190.723 ;
      RECT 9.424999999999999 139.79 9.495 190.723 ;
      RECT 10.855 139.79 10.925 190.723 ;
      RECT 11.334999999999999 139.79 11.405 190.723 ;
      RECT 12.765 139.79 12.835 190.723 ;
      RECT 13.245 139.79 13.315 190.723 ;
      RECT 12.765 139.79 12.835 190.723 ;
      RECT 13.245 139.79 13.315 190.723 ;
      RECT 14.675 139.79 14.745000000000001 190.723 ;
      RECT 15.155 139.79 15.225 190.723 ;
      RECT 16.584999999999997 139.79 16.654999999999998 190.723 ;
      RECT 17.065 139.79 17.135 190.723 ;
      RECT 31.865 139.79 31.935 190.723 ;
      RECT 32.345 139.79 32.415 190.723 ;
      RECT 29.955 139.79 30.025 190.723 ;
      RECT 30.435000000000002 139.79 30.505000000000003 190.723 ;
      RECT 28.044999999999998 139.79 28.115 190.723 ;
      RECT 28.525000000000002 139.79 28.595000000000002 190.723 ;
      RECT 28.044999999999998 139.79 28.115 190.723 ;
      RECT 28.525000000000002 139.79 28.595000000000002 190.723 ;
      RECT 26.134999999999998 139.79 26.205 190.723 ;
      RECT 26.615000000000002 139.79 26.685000000000002 190.723 ;
      RECT 24.224999999999998 139.79 24.294999999999998 190.723 ;
      RECT 24.705000000000002 139.79 24.775000000000002 190.723 ;
      RECT 24.224999999999998 139.79 24.294999999999998 190.723 ;
      RECT 24.705000000000002 139.79 24.775000000000002 190.723 ;
      RECT 22.314999999999998 139.79 22.384999999999998 190.723 ;
      RECT 22.795 139.79 22.865000000000002 190.723 ;
      RECT 20.404999999999998 139.79 20.474999999999998 190.723 ;
      RECT 20.885 139.79 20.955000000000002 190.723 ;
      RECT 20.404999999999998 139.79 20.474999999999998 190.723 ;
      RECT 20.885 139.79 20.955000000000002 190.723 ;
      RECT 18.494999999999997 139.79 18.564999999999998 190.723 ;
      RECT 18.975 139.79 19.045 190.723 ;
      RECT 16.584999999999997 139.79 16.654999999999998 190.723 ;
      RECT 17.065 139.79 17.135 190.723 ;
      RECT 31.865 139.79 31.935 190.723 ;
      RECT 32.345 139.79 32.415 190.723 ;
      RECT 33.775 139.79 33.845 190.723 ;
      RECT 34.255 139.79 34.325 190.723 ;
      RECT 35.684999999999995 139.79 35.754999999999995 190.723 ;
      RECT 36.165 139.79 36.235 190.723 ;
      RECT 35.684999999999995 139.79 35.754999999999995 190.723 ;
      RECT 36.165 139.79 36.235 190.723 ;
      RECT 37.595 139.79 37.665 190.723 ;
      RECT 38.075 139.79 38.145 190.723 ;
      RECT 39.504999999999995 139.79 39.574999999999996 190.723 ;
      RECT 39.985 139.79 40.055 190.723 ;
      RECT 39.504999999999995 139.79 39.574999999999996 190.723 ;
      RECT 39.985 139.79 40.055 190.723 ;
      RECT 41.415 139.79 41.485 190.723 ;
      RECT 41.895 139.79 41.965 190.723 ;
      RECT 43.324999999999996 139.79 43.394999999999996 190.723 ;
      RECT 43.805 139.79 43.875 190.723 ;
      RECT 43.324999999999996 139.79 43.394999999999996 190.723 ;
      RECT 43.805 139.79 43.875 190.723 ;
      RECT 45.235 139.79 45.305 190.723 ;
      RECT 45.715 139.79 45.785000000000004 190.723 ;
      RECT 47.144999999999996 139.79 47.214999999999996 190.723 ;
      RECT 47.625 139.79 47.695 190.723 ;
      RECT 62.425 139.79 62.495 190.723 ;
      RECT 62.905 139.79 62.975 190.723 ;
      RECT 60.515 139.79 60.585 190.723 ;
      RECT 60.995000000000005 139.79 61.065000000000005 190.723 ;
      RECT 58.605 139.79 58.675 190.723 ;
      RECT 59.085 139.79 59.155 190.723 ;
      RECT 58.605 139.79 58.675 190.723 ;
      RECT 59.085 139.79 59.155 190.723 ;
      RECT 56.695 139.79 56.765 190.723 ;
      RECT 57.175000000000004 139.79 57.245000000000005 190.723 ;
      RECT 54.785 139.79 54.855 190.723 ;
      RECT 55.265 139.79 55.335 190.723 ;
      RECT 54.785 139.79 54.855 190.723 ;
      RECT 55.265 139.79 55.335 190.723 ;
      RECT 52.875 139.79 52.945 190.723 ;
      RECT 53.355000000000004 139.79 53.425000000000004 190.723 ;
      RECT 50.964999999999996 139.79 51.035 190.723 ;
      RECT 51.445 139.79 51.515 190.723 ;
      RECT 50.964999999999996 139.79 51.035 190.723 ;
      RECT 51.445 139.79 51.515 190.723 ;
      RECT 49.055 139.79 49.125 190.723 ;
      RECT 49.535000000000004 139.79 49.605000000000004 190.723 ;
      RECT 47.144999999999996 139.79 47.214999999999996 190.723 ;
      RECT 47.625 139.79 47.695 190.723 ;
      RECT 62.425 139.79 62.495 190.723 ;
      RECT 62.905 139.79 62.975 190.723 ;
      RECT 64.33500000000001 139.79 64.405 190.723 ;
      RECT 64.815 139.79 64.88499999999999 190.723 ;
      RECT 66.245 139.79 66.315 190.723 ;
      RECT 66.725 139.79 66.79499999999999 190.723 ;
      RECT 66.245 139.79 66.315 190.723 ;
      RECT 66.725 139.79 66.79499999999999 190.723 ;
      RECT 68.155 139.79 68.225 190.723 ;
      RECT 68.635 139.79 68.705 190.723 ;
      RECT 70.06500000000001 139.79 70.135 190.723 ;
      RECT 70.545 139.79 70.615 190.723 ;
      RECT 70.06500000000001 139.79 70.135 190.723 ;
      RECT 70.545 139.79 70.615 190.723 ;
      RECT 71.97500000000001 139.79 72.045 190.723 ;
      RECT 72.455 139.79 72.52499999999999 190.723 ;
      RECT 73.885 139.79 73.955 190.723 ;
      RECT 74.365 139.79 74.43499999999999 190.723 ;
      RECT 73.885 139.79 73.955 190.723 ;
      RECT 74.365 139.79 74.43499999999999 190.723 ;
      RECT 75.795 139.79 75.865 190.723 ;
      RECT 76.275 139.79 76.345 190.723 ;
      RECT 77.70500000000001 139.79 77.775 190.723 ;
      RECT 78.185 139.79 78.255 190.723 ;
      RECT 92.985 139.79 93.05499999999999 190.723 ;
      RECT 93.465 139.79 93.535 190.723 ;
      RECT 91.075 139.79 91.145 190.723 ;
      RECT 91.555 139.79 91.625 190.723 ;
      RECT 89.165 139.79 89.235 190.723 ;
      RECT 89.645 139.79 89.71499999999999 190.723 ;
      RECT 89.165 139.79 89.235 190.723 ;
      RECT 89.645 139.79 89.71499999999999 190.723 ;
      RECT 87.25500000000001 139.79 87.325 190.723 ;
      RECT 87.735 139.79 87.80499999999999 190.723 ;
      RECT 85.345 139.79 85.41499999999999 190.723 ;
      RECT 85.825 139.79 85.895 190.723 ;
      RECT 85.345 139.79 85.41499999999999 190.723 ;
      RECT 85.825 139.79 85.895 190.723 ;
      RECT 83.435 139.79 83.505 190.723 ;
      RECT 83.915 139.79 83.985 190.723 ;
      RECT 81.525 139.79 81.595 190.723 ;
      RECT 82.005 139.79 82.07499999999999 190.723 ;
      RECT 81.525 139.79 81.595 190.723 ;
      RECT 82.005 139.79 82.07499999999999 190.723 ;
      RECT 79.61500000000001 139.79 79.685 190.723 ;
      RECT 80.095 139.79 80.16499999999999 190.723 ;
      RECT 77.70500000000001 139.79 77.775 190.723 ;
      RECT 78.185 139.79 78.255 190.723 ;
      RECT 92.985 139.79 93.05499999999999 190.723 ;
      RECT 93.465 139.79 93.535 190.723 ;
      RECT 94.89500000000001 139.79 94.965 190.723 ;
      RECT 95.375 139.79 95.445 190.723 ;
      RECT 96.805 139.79 96.875 190.723 ;
      RECT 97.285 139.79 97.35499999999999 190.723 ;
      RECT 96.805 139.79 96.875 190.723 ;
      RECT 97.285 139.79 97.35499999999999 190.723 ;
      RECT 98.715 139.79 98.785 190.723 ;
      RECT 99.19500000000001 139.79 99.265 190.723 ;
      RECT 100.625 139.79 100.695 190.723 ;
      RECT 101.105 139.79 101.175 190.723 ;
      RECT 100.625 139.79 100.695 190.723 ;
      RECT 101.105 139.79 101.175 190.723 ;
      RECT 102.53500000000001 139.79 102.605 190.723 ;
      RECT 103.015 139.79 103.085 190.723 ;
      RECT 104.44500000000001 139.79 104.515 190.723 ;
      RECT 104.925 139.79 104.99499999999999 190.723 ;
      RECT 104.44500000000001 139.79 104.515 190.723 ;
      RECT 104.925 139.79 104.99499999999999 190.723 ;
      RECT 106.355 139.79 106.425 190.723 ;
      RECT 106.83500000000001 139.79 106.905 190.723 ;
      RECT 108.265 139.79 108.335 190.723 ;
      RECT 108.745 139.79 108.815 190.723 ;
      RECT 123.545 139.79 123.615 190.723 ;
      RECT 124.025 139.79 124.095 190.723 ;
      RECT 121.635 139.79 121.705 190.723 ;
      RECT 122.115 139.79 122.18499999999999 190.723 ;
      RECT 119.72500000000001 139.79 119.795 190.723 ;
      RECT 120.205 139.79 120.27499999999999 190.723 ;
      RECT 119.72500000000001 139.79 119.795 190.723 ;
      RECT 120.205 139.79 120.27499999999999 190.723 ;
      RECT 117.81500000000001 139.79 117.885 190.723 ;
      RECT 118.295 139.79 118.365 190.723 ;
      RECT 115.905 139.79 115.975 190.723 ;
      RECT 116.385 139.79 116.455 190.723 ;
      RECT 115.905 139.79 115.975 190.723 ;
      RECT 116.385 139.79 116.455 190.723 ;
      RECT 113.995 139.79 114.065 190.723 ;
      RECT 114.475 139.79 114.54499999999999 190.723 ;
      RECT 112.08500000000001 139.79 112.155 190.723 ;
      RECT 112.565 139.79 112.63499999999999 190.723 ;
      RECT 112.08500000000001 139.79 112.155 190.723 ;
      RECT 112.565 139.79 112.63499999999999 190.723 ;
      RECT 110.17500000000001 139.79 110.245 190.723 ;
      RECT 110.655 139.79 110.725 190.723 ;
      RECT 108.265 139.79 108.335 190.723 ;
      RECT 108.745 139.79 108.815 190.723 ;
      RECT 170.26500000000001 139.79 170.335 190.723 ;
      RECT 170.745 139.79 170.815 190.723 ;
      RECT 172.175 139.79 172.245 190.723 ;
      RECT 172.655 139.79 172.725 190.723 ;
      RECT 174.085 139.79 174.155 190.723 ;
      RECT 174.565 139.79 174.635 190.723 ;
      RECT 174.085 139.79 174.155 190.723 ;
      RECT 174.565 139.79 174.635 190.723 ;
      RECT 175.995 139.79 176.065 190.723 ;
      RECT 176.475 139.79 176.545 190.723 ;
      RECT 177.905 139.79 177.975 190.723 ;
      RECT 178.385 139.79 178.45499999999998 190.723 ;
      RECT 177.905 139.79 177.975 190.723 ;
      RECT 178.385 139.79 178.45499999999998 190.723 ;
      RECT 179.815 139.79 179.885 190.723 ;
      RECT 180.295 139.79 180.36499999999998 190.723 ;
      RECT 181.725 139.79 181.795 190.723 ;
      RECT 182.205 139.79 182.275 190.723 ;
      RECT 181.725 139.79 181.795 190.723 ;
      RECT 182.205 139.79 182.275 190.723 ;
      RECT 183.63500000000002 139.79 183.705 190.723 ;
      RECT 184.115 139.79 184.185 190.723 ;
      RECT 185.54500000000002 139.79 185.615 190.723 ;
      RECT 186.025 139.79 186.095 190.723 ;
      RECT 200.82500000000002 139.79 200.895 190.723 ;
      RECT 201.305 139.79 201.375 190.723 ;
      RECT 198.915 139.79 198.98499999999999 190.723 ;
      RECT 199.395 139.79 199.465 190.723 ;
      RECT 197.005 139.79 197.075 190.723 ;
      RECT 197.485 139.79 197.555 190.723 ;
      RECT 197.005 139.79 197.075 190.723 ;
      RECT 197.485 139.79 197.555 190.723 ;
      RECT 195.095 139.79 195.165 190.723 ;
      RECT 195.575 139.79 195.64499999999998 190.723 ;
      RECT 193.185 139.79 193.255 190.723 ;
      RECT 193.665 139.79 193.73499999999999 190.723 ;
      RECT 193.185 139.79 193.255 190.723 ;
      RECT 193.665 139.79 193.73499999999999 190.723 ;
      RECT 191.275 139.79 191.345 190.723 ;
      RECT 191.755 139.79 191.825 190.723 ;
      RECT 189.365 139.79 189.435 190.723 ;
      RECT 189.845 139.79 189.915 190.723 ;
      RECT 189.365 139.79 189.435 190.723 ;
      RECT 189.845 139.79 189.915 190.723 ;
      RECT 187.455 139.79 187.525 190.723 ;
      RECT 187.935 139.79 188.005 190.723 ;
      RECT 185.54500000000002 139.79 185.615 190.723 ;
      RECT 186.025 139.79 186.095 190.723 ;
      RECT 200.82500000000002 139.79 200.895 190.723 ;
      RECT 201.305 139.79 201.375 190.723 ;
      RECT 202.735 139.79 202.805 190.723 ;
      RECT 203.215 139.79 203.285 190.723 ;
      RECT 204.645 139.79 204.715 190.723 ;
      RECT 205.125 139.79 205.195 190.723 ;
      RECT 204.645 139.79 204.715 190.723 ;
      RECT 205.125 139.79 205.195 190.723 ;
      RECT 206.555 139.79 206.625 190.723 ;
      RECT 207.035 139.79 207.105 190.723 ;
      RECT 208.465 139.79 208.535 190.723 ;
      RECT 208.945 139.79 209.015 190.723 ;
      RECT 208.465 139.79 208.535 190.723 ;
      RECT 208.945 139.79 209.015 190.723 ;
      RECT 210.375 139.79 210.445 190.723 ;
      RECT 210.855 139.79 210.92499999999998 190.723 ;
      RECT 212.285 139.79 212.355 190.723 ;
      RECT 212.76500000000001 139.79 212.835 190.723 ;
      RECT 212.285 139.79 212.355 190.723 ;
      RECT 212.76500000000001 139.79 212.835 190.723 ;
      RECT 214.195 139.79 214.265 190.723 ;
      RECT 214.675 139.79 214.745 190.723 ;
      RECT 216.10500000000002 139.79 216.175 190.723 ;
      RECT 216.585 139.79 216.655 190.723 ;
      RECT 231.38500000000002 139.79 231.455 190.723 ;
      RECT 231.865 139.79 231.935 190.723 ;
      RECT 229.475 139.79 229.545 190.723 ;
      RECT 229.955 139.79 230.025 190.723 ;
      RECT 227.565 139.79 227.635 190.723 ;
      RECT 228.045 139.79 228.11499999999998 190.723 ;
      RECT 227.565 139.79 227.635 190.723 ;
      RECT 228.045 139.79 228.11499999999998 190.723 ;
      RECT 225.655 139.79 225.725 190.723 ;
      RECT 226.135 139.79 226.20499999999998 190.723 ;
      RECT 223.745 139.79 223.815 190.723 ;
      RECT 224.225 139.79 224.295 190.723 ;
      RECT 223.745 139.79 223.815 190.723 ;
      RECT 224.225 139.79 224.295 190.723 ;
      RECT 221.835 139.79 221.905 190.723 ;
      RECT 222.315 139.79 222.385 190.723 ;
      RECT 219.925 139.79 219.995 190.723 ;
      RECT 220.405 139.79 220.475 190.723 ;
      RECT 219.925 139.79 219.995 190.723 ;
      RECT 220.405 139.79 220.475 190.723 ;
      RECT 218.01500000000001 139.79 218.085 190.723 ;
      RECT 218.495 139.79 218.565 190.723 ;
      RECT 216.10500000000002 139.79 216.175 190.723 ;
      RECT 216.585 139.79 216.655 190.723 ;
      RECT 231.38500000000002 139.79 231.455 190.723 ;
      RECT 231.865 139.79 231.935 190.723 ;
      RECT 233.29500000000002 139.79 233.365 190.723 ;
      RECT 233.775 139.79 233.845 190.723 ;
      RECT 235.205 139.79 235.275 190.723 ;
      RECT 235.685 139.79 235.755 190.723 ;
      RECT 235.205 139.79 235.275 190.723 ;
      RECT 235.685 139.79 235.755 190.723 ;
      RECT 237.115 139.79 237.185 190.723 ;
      RECT 237.595 139.79 237.665 190.723 ;
      RECT 239.025 139.79 239.095 190.723 ;
      RECT 239.505 139.79 239.575 190.723 ;
      RECT 239.025 139.79 239.095 190.723 ;
      RECT 239.505 139.79 239.575 190.723 ;
      RECT 240.935 139.79 241.005 190.723 ;
      RECT 241.415 139.79 241.48499999999999 190.723 ;
      RECT 242.845 139.79 242.915 190.723 ;
      RECT 243.325 139.79 243.39499999999998 190.723 ;
      RECT 242.845 139.79 242.915 190.723 ;
      RECT 243.325 139.79 243.39499999999998 190.723 ;
      RECT 244.755 139.79 244.825 190.723 ;
      RECT 245.235 139.79 245.305 190.723 ;
      RECT 246.665 139.79 246.73499999999999 190.723 ;
      RECT 247.145 139.79 247.215 190.723 ;
      RECT 261.945 139.79 262.015 190.723 ;
      RECT 262.425 139.79 262.495 190.723 ;
      RECT 260.03499999999997 139.79 260.10499999999996 190.723 ;
      RECT 260.51500000000004 139.79 260.58500000000004 190.723 ;
      RECT 258.125 139.79 258.195 190.723 ;
      RECT 258.605 139.79 258.675 190.723 ;
      RECT 258.125 139.79 258.195 190.723 ;
      RECT 258.605 139.79 258.675 190.723 ;
      RECT 256.215 139.79 256.28499999999997 190.723 ;
      RECT 256.69500000000005 139.79 256.76500000000004 190.723 ;
      RECT 254.305 139.79 254.375 190.723 ;
      RECT 254.785 139.79 254.855 190.723 ;
      RECT 254.305 139.79 254.375 190.723 ;
      RECT 254.785 139.79 254.855 190.723 ;
      RECT 252.395 139.79 252.465 190.723 ;
      RECT 252.875 139.79 252.945 190.723 ;
      RECT 250.485 139.79 250.555 190.723 ;
      RECT 250.965 139.79 251.035 190.723 ;
      RECT 250.485 139.79 250.555 190.723 ;
      RECT 250.965 139.79 251.035 190.723 ;
      RECT 248.57500000000002 139.79 248.645 190.723 ;
      RECT 249.055 139.79 249.125 190.723 ;
      RECT 246.665 139.79 246.73499999999999 190.723 ;
      RECT 247.145 139.79 247.215 190.723 ;
      RECT 261.945 139.79 262.015 190.723 ;
      RECT 262.425 139.79 262.495 190.723 ;
      RECT 263.85499999999996 139.79 263.92499999999995 190.723 ;
      RECT 264.33500000000004 139.79 264.40500000000003 190.723 ;
      RECT 265.765 139.79 265.835 190.723 ;
      RECT 266.245 139.79 266.315 190.723 ;
      RECT 265.765 139.79 265.835 190.723 ;
      RECT 266.245 139.79 266.315 190.723 ;
      RECT 267.67499999999995 139.79 267.74499999999995 190.723 ;
      RECT 268.15500000000003 139.79 268.225 190.723 ;
      RECT 269.585 139.79 269.655 190.723 ;
      RECT 270.06500000000005 139.79 270.13500000000005 190.723 ;
      RECT 269.585 139.79 269.655 190.723 ;
      RECT 270.06500000000005 139.79 270.13500000000005 190.723 ;
      RECT 271.495 139.79 271.565 190.723 ;
      RECT 271.975 139.79 272.045 190.723 ;
      RECT 273.405 139.79 273.47499999999997 190.723 ;
      RECT 273.88500000000005 139.79 273.95500000000004 190.723 ;
      RECT 273.405 139.79 273.47499999999997 190.723 ;
      RECT 273.88500000000005 139.79 273.95500000000004 190.723 ;
      RECT 275.315 139.79 275.385 190.723 ;
      RECT 275.795 139.79 275.865 190.723 ;
      RECT 277.22499999999997 139.79 277.29499999999996 190.723 ;
      RECT 277.70500000000004 139.79 277.77500000000003 190.723 ;
      RECT 292.505 139.79 292.575 190.723 ;
      RECT 292.985 139.79 293.055 190.723 ;
      RECT 290.59499999999997 139.79 290.66499999999996 190.723 ;
      RECT 291.07500000000005 139.79 291.14500000000004 190.723 ;
      RECT 288.685 139.79 288.755 190.723 ;
      RECT 289.165 139.79 289.235 190.723 ;
      RECT 288.685 139.79 288.755 190.723 ;
      RECT 289.165 139.79 289.235 190.723 ;
      RECT 286.775 139.79 286.84499999999997 190.723 ;
      RECT 287.25500000000005 139.79 287.32500000000005 190.723 ;
      RECT 284.86499999999995 139.79 284.93499999999995 190.723 ;
      RECT 285.345 139.79 285.415 190.723 ;
      RECT 284.86499999999995 139.79 284.93499999999995 190.723 ;
      RECT 285.345 139.79 285.415 190.723 ;
      RECT 282.955 139.79 283.025 190.723 ;
      RECT 283.435 139.79 283.505 190.723 ;
      RECT 281.04499999999996 139.79 281.11499999999995 190.723 ;
      RECT 281.52500000000003 139.79 281.595 190.723 ;
      RECT 281.04499999999996 139.79 281.11499999999995 190.723 ;
      RECT 281.52500000000003 139.79 281.595 190.723 ;
      RECT 279.135 139.79 279.205 190.723 ;
      RECT 279.615 139.79 279.685 190.723 ;
      RECT 277.22499999999997 139.79 277.29499999999996 190.723 ;
      RECT 277.70500000000004 139.79 277.77500000000003 190.723 ;
      RECT 0.0 0.0 0.35 326.068 ;
      RECT 0.9 0.0 1.305 326.068 ;
      RECT 1.855 0.0 2.26 326.068 ;
      RECT 2.81 0.0 3.215 326.068 ;
      RECT 3.765 0.0 4.17 326.068 ;
      RECT 4.72 0.0 5.125 326.068 ;
      RECT 5.675 0.0 6.08 326.068 ;
      RECT 6.63 0.0 7.035 326.068 ;
      RECT 7.585 0.0 7.99 326.068 ;
      RECT 8.54 0.0 8.945 326.068 ;
      RECT 9.495 0.0 9.9 326.068 ;
      RECT 10.45 0.0 10.855 326.068 ;
      RECT 11.405 0.0 11.81 326.068 ;
      RECT 12.36 0.0 12.765 326.068 ;
      RECT 13.315 0.0 13.72 326.068 ;
      RECT 14.27 0.0 14.675 326.068 ;
      RECT 15.225 0.0 15.63 326.068 ;
      RECT 16.18 0.0 16.584999999999997 326.068 ;
      RECT 17.135 0.0 17.54 326.068 ;
      RECT 18.09 0.0 18.494999999999997 326.068 ;
      RECT 19.045 0.0 19.45 326.068 ;
      RECT 20.0 0.0 20.404999999999998 326.068 ;
      RECT 20.955000000000002 0.0 21.36 326.068 ;
      RECT 21.91 0.0 22.314999999999998 326.068 ;
      RECT 22.865000000000002 0.0 23.27 326.068 ;
      RECT 23.82 0.0 24.224999999999998 326.068 ;
      RECT 24.775000000000002 0.0 25.18 326.068 ;
      RECT 25.73 0.0 26.134999999999998 326.068 ;
      RECT 26.685000000000002 0.0 27.09 326.068 ;
      RECT 27.64 0.0 28.044999999999998 326.068 ;
      RECT 28.595000000000002 0.0 29.0 326.068 ;
      RECT 29.55 0.0 29.955 326.068 ;
      RECT 30.505000000000003 0.0 30.91 326.068 ;
      RECT 31.46 0.0 31.865 326.068 ;
      RECT 32.415 0.0 32.82 326.068 ;
      RECT 33.370000000000005 0.0 33.775 326.068 ;
      RECT 34.325 0.0 34.73 326.068 ;
      RECT 35.28 0.0 35.684999999999995 326.068 ;
      RECT 36.235 0.0 36.64 326.068 ;
      RECT 37.190000000000005 0.0 37.595 326.068 ;
      RECT 38.145 0.0 38.55 326.068 ;
      RECT 39.1 0.0 39.504999999999995 326.068 ;
      RECT 40.055 0.0 40.46 326.068 ;
      RECT 41.01 0.0 41.415 326.068 ;
      RECT 41.965 0.0 42.37 326.068 ;
      RECT 42.92 0.0 43.324999999999996 326.068 ;
      RECT 43.875 0.0 44.28 326.068 ;
      RECT 44.83 0.0 45.235 326.068 ;
      RECT 45.785000000000004 0.0 46.19 326.068 ;
      RECT 46.74 0.0 47.144999999999996 326.068 ;
      RECT 47.695 0.0 48.1 326.068 ;
      RECT 48.65 0.0 49.055 326.068 ;
      RECT 49.605000000000004 0.0 50.01 326.068 ;
      RECT 50.56 0.0 50.964999999999996 326.068 ;
      RECT 51.515 0.0 51.92 326.068 ;
      RECT 52.47 0.0 52.875 326.068 ;
      RECT 53.425000000000004 0.0 53.83 326.068 ;
      RECT 54.38 0.0 54.785 326.068 ;
      RECT 55.335 0.0 55.74 326.068 ;
      RECT 56.29 0.0 56.695 326.068 ;
      RECT 57.245000000000005 0.0 57.65 326.068 ;
      RECT 58.2 0.0 58.605 326.068 ;
      RECT 59.155 0.0 59.559999999999995 326.068 ;
      RECT 60.11 0.0 60.515 326.068 ;
      RECT 61.065000000000005 0.0 61.47 326.068 ;
      RECT 62.02 0.0 62.425 326.068 ;
      RECT 62.975 0.0 63.379999999999995 326.068 ;
      RECT 63.93 0.0 64.33500000000001 326.068 ;
      RECT 64.88499999999999 0.0 65.29 326.068 ;
      RECT 65.83999999999999 0.0 66.245 326.068 ;
      RECT 66.79499999999999 0.0 67.2 326.068 ;
      RECT 67.75 0.0 68.155 326.068 ;
      RECT 68.705 0.0 69.11 326.068 ;
      RECT 69.66 0.0 70.06500000000001 326.068 ;
      RECT 70.615 0.0 71.02000000000001 326.068 ;
      RECT 71.57 0.0 71.97500000000001 326.068 ;
      RECT 72.52499999999999 0.0 72.93 326.068 ;
      RECT 73.47999999999999 0.0 73.885 326.068 ;
      RECT 74.43499999999999 0.0 74.84 326.068 ;
      RECT 75.39 0.0 75.795 326.068 ;
      RECT 76.345 0.0 76.75 326.068 ;
      RECT 77.3 0.0 77.70500000000001 326.068 ;
      RECT 78.255 0.0 78.66000000000001 326.068 ;
      RECT 79.21 0.0 79.61500000000001 326.068 ;
      RECT 80.16499999999999 0.0 80.57000000000001 326.068 ;
      RECT 81.11999999999999 0.0 81.525 326.068 ;
      RECT 82.07499999999999 0.0 82.48 326.068 ;
      RECT 83.03 0.0 83.435 326.068 ;
      RECT 83.985 0.0 84.39 326.068 ;
      RECT 84.94 0.0 85.345 326.068 ;
      RECT 85.895 0.0 86.30000000000001 326.068 ;
      RECT 86.85 0.0 87.25500000000001 326.068 ;
      RECT 87.80499999999999 0.0 88.21000000000001 326.068 ;
      RECT 88.75999999999999 0.0 89.165 326.068 ;
      RECT 89.71499999999999 0.0 90.12 326.068 ;
      RECT 90.66999999999999 0.0 91.075 326.068 ;
      RECT 91.625 0.0 92.03 326.068 ;
      RECT 92.58 0.0 92.985 326.068 ;
      RECT 93.535 0.0 93.94000000000001 326.068 ;
      RECT 94.49 0.0 94.89500000000001 326.068 ;
      RECT 95.445 0.0 95.85000000000001 326.068 ;
      RECT 96.39999999999999 0.0 96.805 326.068 ;
      RECT 97.35499999999999 0.0 97.76 326.068 ;
      RECT 98.30999999999999 0.0 98.715 326.068 ;
      RECT 99.265 0.0 99.67 326.068 ;
      RECT 100.22 0.0 100.625 326.068 ;
      RECT 101.175 0.0 101.58000000000001 326.068 ;
      RECT 102.13 0.0 102.53500000000001 326.068 ;
      RECT 103.085 0.0 103.49000000000001 326.068 ;
      RECT 104.03999999999999 0.0 104.44500000000001 326.068 ;
      RECT 104.99499999999999 0.0 105.4 326.068 ;
      RECT 105.94999999999999 0.0 106.355 326.068 ;
      RECT 106.905 0.0 107.31 326.068 ;
      RECT 107.86 0.0 108.265 326.068 ;
      RECT 108.815 0.0 109.22 326.068 ;
      RECT 109.77 0.0 110.17500000000001 326.068 ;
      RECT 110.725 0.0 111.13000000000001 326.068 ;
      RECT 111.67999999999999 0.0 112.08500000000001 326.068 ;
      RECT 112.63499999999999 0.0 113.04 326.068 ;
      RECT 113.58999999999999 0.0 113.995 326.068 ;
      RECT 114.54499999999999 0.0 114.95 326.068 ;
      RECT 115.5 0.0 115.905 326.068 ;
      RECT 116.455 0.0 116.86 326.068 ;
      RECT 117.41 0.0 117.81500000000001 326.068 ;
      RECT 118.365 0.0 118.77000000000001 326.068 ;
      RECT 119.32 0.0 119.72500000000001 326.068 ;
      RECT 120.27499999999999 0.0 120.68 326.068 ;
      RECT 121.22999999999999 0.0 121.635 326.068 ;
      RECT 122.18499999999999 0.0 122.59 326.068 ;
      RECT 123.14 0.0 123.545 326.068 ;
      RECT 124.095 0.0 124.5 326.068 ;
      RECT 125.05 0.0 126.05000000000001 326.068 ;
      RECT 126.64999999999999 0.0 126.65 326.068 ;
      RECT 127.85 0.0 128.45000000000002 326.068 ;
      RECT 129.04999999999998 0.0 129.65 326.068 ;
      RECT 130.25 0.0 130.85 326.068 ;
      RECT 131.45 0.0 132.05 326.068 ;
      RECT 132.65 0.0 133.25 326.068 ;
      RECT 133.85 0.0 134.45000000000002 326.068 ;
      RECT 135.04999999999998 0.0 135.65 326.068 ;
      RECT 136.25 0.0 137.45000000000002 326.068 ;
      RECT 138.04999999999998 0.0 138.05 326.068 ;
      RECT 139.25 0.0 139.85 326.068 ;
      RECT 140.45 0.0 141.05 326.068 ;
      RECT 141.65 0.0 142.85 326.068 ;
      RECT 143.45 0.0 144.05 326.068 ;
      RECT 144.65 0.0 145.25 326.068 ;
      RECT 146.45 0.0 146.45000000000002 326.068 ;
      RECT 147.04999999999998 0.0 147.31 326.068 ;
      RECT 148.51 0.0 148.51000000000002 326.068 ;
      RECT 149.10999999999999 0.0 149.71 326.068 ;
      RECT 150.31 0.0 150.91 326.068 ;
      RECT 151.51 0.0 152.71 326.068 ;
      RECT 153.31 0.0 153.91 326.068 ;
      RECT 154.51 0.0 155.11 326.068 ;
      RECT 156.91 0.0 158.11 326.068 ;
      RECT 158.71 0.0 159.31 326.068 ;
      RECT 159.91 0.0 160.51000000000002 326.068 ;
      RECT 161.10999999999999 0.0 161.71 326.068 ;
      RECT 162.31 0.0 162.91 326.068 ;
      RECT 163.51 0.0 164.11 326.068 ;
      RECT 164.71 0.0 165.31 326.068 ;
      RECT 165.91 0.0 166.51000000000002 326.068 ;
      RECT 167.10999999999999 0.0 167.11 326.068 ;
      RECT 168.31 0.0 169.31 326.068 ;
      RECT 169.85999999999999 0.0 170.26500000000001 326.068 ;
      RECT 170.815 0.0 171.22 326.068 ;
      RECT 171.76999999999998 0.0 172.175 326.068 ;
      RECT 172.725 0.0 173.13 326.068 ;
      RECT 173.68 0.0 174.085 326.068 ;
      RECT 174.635 0.0 175.04 326.068 ;
      RECT 175.59 0.0 175.995 326.068 ;
      RECT 176.545 0.0 176.95000000000002 326.068 ;
      RECT 177.5 0.0 177.905 326.068 ;
      RECT 178.45499999999998 0.0 178.86 326.068 ;
      RECT 179.41 0.0 179.815 326.068 ;
      RECT 180.36499999999998 0.0 180.77 326.068 ;
      RECT 181.32 0.0 181.725 326.068 ;
      RECT 182.275 0.0 182.68 326.068 ;
      RECT 183.23 0.0 183.63500000000002 326.068 ;
      RECT 184.185 0.0 184.59 326.068 ;
      RECT 185.14 0.0 185.54500000000002 326.068 ;
      RECT 186.095 0.0 186.5 326.068 ;
      RECT 187.04999999999998 0.0 187.455 326.068 ;
      RECT 188.005 0.0 188.41 326.068 ;
      RECT 188.96 0.0 189.365 326.068 ;
      RECT 189.915 0.0 190.32 326.068 ;
      RECT 190.87 0.0 191.275 326.068 ;
      RECT 191.825 0.0 192.23000000000002 326.068 ;
      RECT 192.78 0.0 193.185 326.068 ;
      RECT 193.73499999999999 0.0 194.14000000000001 326.068 ;
      RECT 194.69 0.0 195.095 326.068 ;
      RECT 195.64499999999998 0.0 196.05 326.068 ;
      RECT 196.6 0.0 197.005 326.068 ;
      RECT 197.555 0.0 197.96 326.068 ;
      RECT 198.51 0.0 198.915 326.068 ;
      RECT 199.465 0.0 199.87 326.068 ;
      RECT 200.42 0.0 200.82500000000002 326.068 ;
      RECT 201.375 0.0 201.78 326.068 ;
      RECT 202.32999999999998 0.0 202.735 326.068 ;
      RECT 203.285 0.0 203.69 326.068 ;
      RECT 204.23999999999998 0.0 204.645 326.068 ;
      RECT 205.195 0.0 205.6 326.068 ;
      RECT 206.15 0.0 206.555 326.068 ;
      RECT 207.105 0.0 207.51000000000002 326.068 ;
      RECT 208.06 0.0 208.465 326.068 ;
      RECT 209.015 0.0 209.42000000000002 326.068 ;
      RECT 209.97 0.0 210.375 326.068 ;
      RECT 210.92499999999998 0.0 211.33 326.068 ;
      RECT 211.88 0.0 212.285 326.068 ;
      RECT 212.835 0.0 213.24 326.068 ;
      RECT 213.79 0.0 214.195 326.068 ;
      RECT 214.745 0.0 215.15 326.068 ;
      RECT 215.7 0.0 216.10500000000002 326.068 ;
      RECT 216.655 0.0 217.06 326.068 ;
      RECT 217.60999999999999 0.0 218.01500000000001 326.068 ;
      RECT 218.565 0.0 218.97 326.068 ;
      RECT 219.51999999999998 0.0 219.925 326.068 ;
      RECT 220.475 0.0 220.88 326.068 ;
      RECT 221.43 0.0 221.835 326.068 ;
      RECT 222.385 0.0 222.79 326.068 ;
      RECT 223.34 0.0 223.745 326.068 ;
      RECT 224.295 0.0 224.70000000000002 326.068 ;
      RECT 225.25 0.0 225.655 326.068 ;
      RECT 226.20499999999998 0.0 226.61 326.068 ;
      RECT 227.16 0.0 227.565 326.068 ;
      RECT 228.11499999999998 0.0 228.52 326.068 ;
      RECT 229.07 0.0 229.475 326.068 ;
      RECT 230.025 0.0 230.43 326.068 ;
      RECT 230.98 0.0 231.38500000000002 326.068 ;
      RECT 231.935 0.0 232.34 326.068 ;
      RECT 232.89 0.0 233.29500000000002 326.068 ;
      RECT 233.845 0.0 234.25 326.068 ;
      RECT 234.79999999999998 0.0 235.205 326.068 ;
      RECT 235.755 0.0 236.16 326.068 ;
      RECT 236.71 0.0 237.115 326.068 ;
      RECT 237.665 0.0 238.07 326.068 ;
      RECT 238.62 0.0 239.025 326.068 ;
      RECT 239.575 0.0 239.98000000000002 326.068 ;
      RECT 240.53 0.0 240.935 326.068 ;
      RECT 241.48499999999999 0.0 241.89000000000001 326.068 ;
      RECT 242.44 0.0 242.845 326.068 ;
      RECT 243.39499999999998 0.0 243.8 326.068 ;
      RECT 244.35 0.0 244.755 326.068 ;
      RECT 245.305 0.0 245.71 326.068 ;
      RECT 246.26 0.0 246.665 326.068 ;
      RECT 247.215 0.0 247.62 326.068 ;
      RECT 248.17 0.0 248.57500000000002 326.068 ;
      RECT 249.125 0.0 249.53 326.068 ;
      RECT 250.07999999999998 0.0 250.485 326.068 ;
      RECT 251.035 0.0 251.44 326.068 ;
      RECT 251.98999999999998 0.0 252.395 326.068 ;
      RECT 252.945 0.0 253.35 326.068 ;
      RECT 253.9 0.0 254.305 326.068 ;
      RECT 254.855 0.0 255.26000000000002 326.068 ;
      RECT 255.81 0.0 256.215 326.068 ;
      RECT 256.76500000000004 0.0 257.16999999999996 326.068 ;
      RECT 257.72 0.0 258.125 326.068 ;
      RECT 258.675 0.0 259.08 326.068 ;
      RECT 259.63 0.0 260.03499999999997 326.068 ;
      RECT 260.58500000000004 0.0 260.98999999999995 326.068 ;
      RECT 261.54 0.0 261.945 326.068 ;
      RECT 262.495 0.0 262.9 326.068 ;
      RECT 263.45000000000005 0.0 263.85499999999996 326.068 ;
      RECT 264.40500000000003 0.0 264.81 326.068 ;
      RECT 265.36 0.0 265.765 326.068 ;
      RECT 266.315 0.0 266.71999999999997 326.068 ;
      RECT 267.27000000000004 0.0 267.67499999999995 326.068 ;
      RECT 268.225 0.0 268.63 326.068 ;
      RECT 269.18 0.0 269.585 326.068 ;
      RECT 270.13500000000005 0.0 270.53999999999996 326.068 ;
      RECT 271.09000000000003 0.0 271.495 326.068 ;
      RECT 272.045 0.0 272.45 326.068 ;
      RECT 273.0 0.0 273.405 326.068 ;
      RECT 273.95500000000004 0.0 274.35999999999996 326.068 ;
      RECT 274.91 0.0 275.315 326.068 ;
      RECT 275.865 0.0 276.27 326.068 ;
      RECT 276.82000000000005 0.0 277.22499999999997 326.068 ;
      RECT 277.77500000000003 0.0 278.17999999999995 326.068 ;
      RECT 278.73 0.0 279.135 326.068 ;
      RECT 279.685 0.0 280.09 326.068 ;
      RECT 280.64000000000004 0.0 281.04499999999996 326.068 ;
      RECT 281.595 0.0 282.0 326.068 ;
      RECT 282.55 0.0 282.955 326.068 ;
      RECT 283.505 0.0 283.90999999999997 326.068 ;
      RECT 284.46000000000004 0.0 284.86499999999995 326.068 ;
      RECT 285.415 0.0 285.82 326.068 ;
      RECT 286.37 0.0 286.775 326.068 ;
      RECT 287.32500000000005 0.0 287.72999999999996 326.068 ;
      RECT 288.28000000000003 0.0 288.685 326.068 ;
      RECT 289.235 0.0 289.64 326.068 ;
      RECT 290.19 0.0 290.59499999999997 326.068 ;
      RECT 291.14500000000004 0.0 291.54999999999995 326.068 ;
      RECT 292.1 0.0 292.505 326.068 ;
      RECT 293.055 0.0 293.46 326.068 ;
      RECT 294.01000000000005 0.0 294.36 326.068 ;
  END
END dpram16x4096
END LIBRARY