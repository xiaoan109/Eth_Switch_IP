// removed module with interface ports: RdCtrlTop1Ch
