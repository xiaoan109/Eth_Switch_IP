// removed module with interface ports: DcpTag16x16
