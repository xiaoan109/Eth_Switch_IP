// removed module with interface ports: RdScheTop
