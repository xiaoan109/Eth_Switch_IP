
#     Copyright (c) 2024 SMIC             
#     Filename:      S55NLLGDPH_X512Y8D16_BW.lef
#     IP code:       S55NLLGDPH
#     Version:       1.3.a
#     CreateDate:    May 18, 2024        
                    
#    LEF for General Dual-Port SRAM
#    SMIC 55nm LL Logic Process

#    Configuration: -instname S55NLLGDPH_X512Y8D16_BW -rows 512 -bits 16 -mux 8 
#    Redundancy: Off
#    Bit-Write: On


# DISCLAIMER                                                                      
#                                                                                   
#   SMIC hereby provides the quality information to you but makes no claims,      
# promises or guarantees about the accuracy, completeness, or adequacy of the     
# information herein. The information contained herein is provided on an "AS IS"  
# basis without any warranty, and SMIC assumes no obligation to provide support   
# of any kind or otherwise maintain the information.                                
#   SMIC disclaims any representation that the information does not infringe any  
# intellectual property rights or proprietary rights of any third parties. SMIC   
# makes no other warranty, whether express, implied or statutory as to any        
# matter whatsoever, including but not limited to the accuracy or sufficiency of  
# any information or the merchantability and fitness for a particular purpose.    
# Neither SMIC nor any of its representatives shall be liable for any cause of    
# action incurred to connect to this service.                                       
#                                                                                 
# STATEMENT OF USE AND CONFIDENTIALITY                                              
#                                                                                   
#   The following/attached material contains confidential and proprietary           
# information of SMIC. This material is based upon information which SMIC           
# considers reliable, but SMIC neither represents nor warrants that such          
# information is accurate or complete, and it must not be relied upon as such.    
# This information was prepared for informational purposes and is for the use     
# by SMIC's customer only. SMIC reserves the right to make changes in the           
# information at any time without notice.                                           
#   No part of this information may be reproduced, transmitted, transcribed,        
# stored in a retrieval system, or translated into any human or computer           
# language, in any form or by any means, electronic, mechanical, magnetic,          
# optical, chemical, manual, or otherwise, without the prior written consent of   
# SMIC. Any unauthorized use or disclosure of this material is strictly             
# prohibited and may be unlawful. By accepting this material, the receiving         
# party shall be deemed to have acknowledged, accepted, and agreed to be bound    
# by the foregoing limitations and restrictions. Thank you.                         
#                                                                                   


VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO S55NLLGDPH_X512Y8D16_BW
 CLASS BLOCK ;
 ORIGIN 0 0 ;
 SYMMETRY X Y R90 ;
 SIZE 313.52 BY 319.25 ;

 PIN AA[0]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 126.995 0 127.195 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 126.995 0 127.195 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 126.995 0 127.195 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END AA[0]

 PIN AA[1]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 130.16 0 130.36 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 130.16 0 130.36 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 130.16 0 130.36 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END AA[1]

 PIN AA[2]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 132.1 0 132.3 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 132.1 0 132.3 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 132.1 0 132.3 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END AA[2]

 PIN AA[3]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 137.475 0 137.675 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 137.475 0 137.675 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 137.475 0 137.675 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END AA[3]

 PIN AA[4]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 140.07 0 140.27 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 140.07 0 140.27 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 140.07 0 140.27 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END AA[4]

 PIN AA[5]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 142.265 0 142.465 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 142.265 0 142.465 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 142.265 0 142.465 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END AA[5]

 PIN WENA
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 143.655 0 143.855 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 143.655 0 143.855 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 143.655 0 143.855 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END WENA

 PIN AA[7]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 146.26 0 146.46 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 146.26 0 146.46 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 146.26 0 146.46 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END AA[7]

 PIN AA[6]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 148.965 0 149.165 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 148.965 0 149.165 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 148.965 0 149.165 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END AA[6]

 PIN AA[10]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 150.56 0 150.76 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 150.56 0 150.76 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 150.56 0 150.76 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END AA[10]

 PIN CLKA
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 151.435 0 151.635 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 151.435 0 151.635 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 151.435 0 151.635 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END CLKA

 PIN CENA
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 152.155 0 152.355 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 152.155 0 152.355 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 152.155 0 152.355 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END CENA

 PIN AA[9]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 153 0 153.2 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 153 0 153.2 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 153 0 153.2 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END AA[9]

 PIN AA[8]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 153.865 0 154.065 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 153.865 0 154.065 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 153.865 0 154.065 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END AA[8]

 PIN AA[11]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 154.71 0 154.91 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 154.71 0 154.91 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 154.71 0 154.91 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END AA[11]

 PIN AB[11]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 158.61 0 158.81 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 158.61 0 158.81 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 158.61 0 158.81 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END AB[11]

 PIN AB[8]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 159.455 0 159.655 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 159.455 0 159.655 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 159.455 0 159.655 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END AB[8]

 PIN AB[9]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 160.32 0 160.52 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 160.32 0 160.52 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 160.32 0 160.52 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END AB[9]

 PIN CENB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 161.165 0 161.365 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 161.165 0 161.365 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 161.165 0 161.365 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END CENB

 PIN CLKB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 161.885 0 162.085 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 161.885 0 162.085 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 161.885 0 162.085 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END CLKB

 PIN AB[10]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 162.76 0 162.96 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 162.76 0 162.96 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 162.76 0 162.96 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END AB[10]

 PIN AB[6]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 164.355 0 164.555 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 164.355 0 164.555 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 164.355 0 164.555 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END AB[6]

 PIN AB[7]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 167.06 0 167.26 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 167.06 0 167.26 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 167.06 0 167.26 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END AB[7]

 PIN WENB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 169.665 0 169.865 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 169.665 0 169.865 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 169.665 0 169.865 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END WENB

 PIN AB[5]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 171.055 0 171.255 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 171.055 0 171.255 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 171.055 0 171.255 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END AB[5]

 PIN AB[4]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 173.25 0 173.45 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 173.25 0 173.45 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 173.25 0 173.45 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END AB[4]

 PIN AB[3]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 175.845 0 176.045 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 175.845 0 176.045 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 175.845 0 176.045 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END AB[3]

 PIN AB[2]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 181.22 0 181.42 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 181.22 0 181.42 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 181.22 0 181.42 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END AB[2]

 PIN AB[1]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 183.16 0 183.36 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 183.16 0 183.36 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 183.16 0 183.36 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END AB[1]

 PIN AB[0]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 186.325 0 186.525 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 186.325 0 186.525 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 186.325 0 186.525 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END AB[0]

 PIN QB[7]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 4.165 0 4.365 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 4.165 0 4.365 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 4.165 0 4.365 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END QB[7]

 PIN DB[7]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 7.025 0 7.225 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 7.025 0 7.225 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 7.025 0 7.225 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END DB[7]

 PIN BWENB[7]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 8.705 0 8.905 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 8.705 0 8.905 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 8.705 0 8.905 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END BWENB[7]

 PIN BWENA[7]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 10.485 0 10.685 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 10.485 0 10.685 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 10.485 0 10.685 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END BWENA[7]

 PIN DA[7]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 12.165 0 12.365 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 12.165 0 12.365 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 12.165 0 12.365 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END DA[7]

 PIN QA[7]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 15.025 0 15.225 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 15.025 0 15.225 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 15.025 0 15.225 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END QA[7]

 PIN QB[6]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 19.445 0 19.645 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 19.445 0 19.645 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 19.445 0 19.645 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END QB[6]

 PIN DB[6]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 22.305 0 22.505 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 22.305 0 22.505 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 22.305 0 22.505 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END DB[6]

 PIN BWENB[6]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 23.985 0 24.185 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 23.985 0 24.185 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 23.985 0 24.185 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END BWENB[6]

 PIN BWENA[6]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 25.765 0 25.965 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 25.765 0 25.965 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 25.765 0 25.965 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END BWENA[6]

 PIN DA[6]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 27.445 0 27.645 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 27.445 0 27.645 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 27.445 0 27.645 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END DA[6]

 PIN QA[6]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 30.305 0 30.505 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 30.305 0 30.505 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 30.305 0 30.505 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END QA[6]

 PIN QB[5]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 34.725 0 34.925 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 34.725 0 34.925 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 34.725 0 34.925 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END QB[5]

 PIN DB[5]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 37.585 0 37.785 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 37.585 0 37.785 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 37.585 0 37.785 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END DB[5]

 PIN BWENB[5]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 39.265 0 39.465 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 39.265 0 39.465 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 39.265 0 39.465 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END BWENB[5]

 PIN BWENA[5]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 41.045 0 41.245 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 41.045 0 41.245 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 41.045 0 41.245 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END BWENA[5]

 PIN DA[5]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 42.725 0 42.925 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 42.725 0 42.925 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 42.725 0 42.925 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END DA[5]

 PIN QA[5]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 45.585 0 45.785 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 45.585 0 45.785 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 45.585 0 45.785 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END QA[5]

 PIN QB[4]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 50.005 0 50.205 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 50.005 0 50.205 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 50.005 0 50.205 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END QB[4]

 PIN DB[4]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 52.865 0 53.065 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 52.865 0 53.065 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 52.865 0 53.065 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END DB[4]

 PIN BWENB[4]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 54.545 0 54.745 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 54.545 0 54.745 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 54.545 0 54.745 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END BWENB[4]

 PIN BWENA[4]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 56.325 0 56.525 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 56.325 0 56.525 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 56.325 0 56.525 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END BWENA[4]

 PIN DA[4]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 58.005 0 58.205 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 58.005 0 58.205 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 58.005 0 58.205 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END DA[4]

 PIN QA[4]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 60.865 0 61.065 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 60.865 0 61.065 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 60.865 0 61.065 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END QA[4]

 PIN QB[3]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 65.285 0 65.485 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 65.285 0 65.485 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 65.285 0 65.485 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END QB[3]

 PIN DB[3]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 68.145 0 68.345 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 68.145 0 68.345 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 68.145 0 68.345 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END DB[3]

 PIN BWENB[3]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 69.825 0 70.025 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 69.825 0 70.025 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 69.825 0 70.025 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END BWENB[3]

 PIN BWENA[3]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 71.605 0 71.805 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 71.605 0 71.805 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 71.605 0 71.805 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END BWENA[3]

 PIN DA[3]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 73.285 0 73.485 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 73.285 0 73.485 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 73.285 0 73.485 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END DA[3]

 PIN QA[3]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 76.145 0 76.345 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 76.145 0 76.345 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 76.145 0 76.345 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END QA[3]

 PIN QB[2]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 80.565 0 80.765 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 80.565 0 80.765 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 80.565 0 80.765 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END QB[2]

 PIN DB[2]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 83.425 0 83.625 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 83.425 0 83.625 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 83.425 0 83.625 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END DB[2]

 PIN BWENB[2]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 85.105 0 85.305 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 85.105 0 85.305 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 85.105 0 85.305 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END BWENB[2]

 PIN BWENA[2]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 86.885 0 87.085 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 86.885 0 87.085 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 86.885 0 87.085 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END BWENA[2]

 PIN DA[2]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 88.565 0 88.765 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 88.565 0 88.765 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 88.565 0 88.765 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END DA[2]

 PIN QA[2]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 91.425 0 91.625 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 91.425 0 91.625 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 91.425 0 91.625 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END QA[2]

 PIN QB[1]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 95.845 0 96.045 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 95.845 0 96.045 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 95.845 0 96.045 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END QB[1]

 PIN DB[1]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 98.705 0 98.905 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 98.705 0 98.905 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 98.705 0 98.905 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END DB[1]

 PIN BWENB[1]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 100.385 0 100.585 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 100.385 0 100.585 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 100.385 0 100.585 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END BWENB[1]

 PIN BWENA[1]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 102.165 0 102.365 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 102.165 0 102.365 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 102.165 0 102.365 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END BWENA[1]

 PIN DA[1]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 103.845 0 104.045 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 103.845 0 104.045 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 103.845 0 104.045 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END DA[1]

 PIN QA[1]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 106.705 0 106.905 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 106.705 0 106.905 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 106.705 0 106.905 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END QA[1]

 PIN QB[0]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 111.125 0 111.325 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 111.125 0 111.325 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 111.125 0 111.325 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END QB[0]

 PIN DB[0]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 113.985 0 114.185 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 113.985 0 114.185 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 113.985 0 114.185 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END DB[0]

 PIN BWENB[0]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 115.665 0 115.865 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 115.665 0 115.865 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 115.665 0 115.865 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END BWENB[0]

 PIN BWENA[0]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 117.445 0 117.645 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 117.445 0 117.645 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 117.445 0 117.645 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END BWENA[0]

 PIN DA[0]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 119.125 0 119.325 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 119.125 0 119.325 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 119.125 0 119.325 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END DA[0]

 PIN QA[0]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 121.985 0 122.185 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 121.985 0 122.185 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 121.985 0 122.185 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END QA[0]

 PIN QA[8]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 191.335 0 191.535 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 191.335 0 191.535 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 191.335 0 191.535 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END QA[8]

 PIN DA[8]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 194.195 0 194.395 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 194.195 0 194.395 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 194.195 0 194.395 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END DA[8]

 PIN BWENA[8]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 195.875 0 196.075 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 195.875 0 196.075 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 195.875 0 196.075 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END BWENA[8]

 PIN BWENB[8]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 197.655 0 197.855 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 197.655 0 197.855 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 197.655 0 197.855 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END BWENB[8]

 PIN DB[8]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 199.335 0 199.535 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 199.335 0 199.535 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 199.335 0 199.535 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END DB[8]

 PIN QB[8]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 202.195 0 202.395 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 202.195 0 202.395 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 202.195 0 202.395 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END QB[8]

 PIN QA[9]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 206.615 0 206.815 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 206.615 0 206.815 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 206.615 0 206.815 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END QA[9]

 PIN DA[9]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 209.475 0 209.675 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 209.475 0 209.675 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 209.475 0 209.675 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END DA[9]

 PIN BWENA[9]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 211.155 0 211.355 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 211.155 0 211.355 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 211.155 0 211.355 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END BWENA[9]

 PIN BWENB[9]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 212.935 0 213.135 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 212.935 0 213.135 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 212.935 0 213.135 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END BWENB[9]

 PIN DB[9]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 214.615 0 214.815 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 214.615 0 214.815 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 214.615 0 214.815 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END DB[9]

 PIN QB[9]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 217.475 0 217.675 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 217.475 0 217.675 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 217.475 0 217.675 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END QB[9]

 PIN QA[10]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 221.895 0 222.095 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 221.895 0 222.095 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 221.895 0 222.095 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END QA[10]

 PIN DA[10]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 224.755 0 224.955 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 224.755 0 224.955 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 224.755 0 224.955 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END DA[10]

 PIN BWENA[10]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 226.435 0 226.635 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 226.435 0 226.635 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 226.435 0 226.635 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END BWENA[10]

 PIN BWENB[10]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 228.215 0 228.415 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 228.215 0 228.415 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 228.215 0 228.415 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END BWENB[10]

 PIN DB[10]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 229.895 0 230.095 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 229.895 0 230.095 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 229.895 0 230.095 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END DB[10]

 PIN QB[10]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 232.755 0 232.955 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 232.755 0 232.955 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 232.755 0 232.955 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END QB[10]

 PIN QA[11]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 237.175 0 237.375 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 237.175 0 237.375 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 237.175 0 237.375 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END QA[11]

 PIN DA[11]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 240.035 0 240.235 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 240.035 0 240.235 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 240.035 0 240.235 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END DA[11]

 PIN BWENA[11]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 241.715 0 241.915 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 241.715 0 241.915 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 241.715 0 241.915 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END BWENA[11]

 PIN BWENB[11]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 243.495 0 243.695 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 243.495 0 243.695 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 243.495 0 243.695 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END BWENB[11]

 PIN DB[11]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 245.175 0 245.375 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 245.175 0 245.375 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 245.175 0 245.375 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END DB[11]

 PIN QB[11]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 248.035 0 248.235 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 248.035 0 248.235 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 248.035 0 248.235 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END QB[11]

 PIN QA[12]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 252.455 0 252.655 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 252.455 0 252.655 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 252.455 0 252.655 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END QA[12]

 PIN DA[12]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 255.315 0 255.515 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 255.315 0 255.515 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 255.315 0 255.515 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END DA[12]

 PIN BWENA[12]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 256.995 0 257.195 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 256.995 0 257.195 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 256.995 0 257.195 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END BWENA[12]

 PIN BWENB[12]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 258.775 0 258.975 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 258.775 0 258.975 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 258.775 0 258.975 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END BWENB[12]

 PIN DB[12]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 260.455 0 260.655 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 260.455 0 260.655 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 260.455 0 260.655 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END DB[12]

 PIN QB[12]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 263.315 0 263.515 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 263.315 0 263.515 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 263.315 0 263.515 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END QB[12]

 PIN QA[13]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 267.735 0 267.935 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 267.735 0 267.935 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 267.735 0 267.935 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END QA[13]

 PIN DA[13]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 270.595 0 270.795 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 270.595 0 270.795 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 270.595 0 270.795 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END DA[13]

 PIN BWENA[13]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 272.275 0 272.475 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 272.275 0 272.475 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 272.275 0 272.475 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END BWENA[13]

 PIN BWENB[13]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 274.055 0 274.255 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 274.055 0 274.255 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 274.055 0 274.255 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END BWENB[13]

 PIN DB[13]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 275.735 0 275.935 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 275.735 0 275.935 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 275.735 0 275.935 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END DB[13]

 PIN QB[13]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 278.595 0 278.795 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 278.595 0 278.795 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 278.595 0 278.795 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END QB[13]

 PIN QA[14]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 283.015 0 283.215 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 283.015 0 283.215 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 283.015 0 283.215 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END QA[14]

 PIN DA[14]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 285.875 0 286.075 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 285.875 0 286.075 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 285.875 0 286.075 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END DA[14]

 PIN BWENA[14]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 287.555 0 287.755 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 287.555 0 287.755 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 287.555 0 287.755 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END BWENA[14]

 PIN BWENB[14]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 289.335 0 289.535 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 289.335 0 289.535 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 289.335 0 289.535 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END BWENB[14]

 PIN DB[14]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 291.015 0 291.215 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 291.015 0 291.215 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 291.015 0 291.215 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END DB[14]

 PIN QB[14]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 293.875 0 294.075 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 293.875 0 294.075 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 293.875 0 294.075 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END QB[14]

 PIN QA[15]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 298.295 0 298.495 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 298.295 0 298.495 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 298.295 0 298.495 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END QA[15]

 PIN DA[15]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 301.155 0 301.355 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 301.155 0 301.355 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 301.155 0 301.355 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END DA[15]

 PIN BWENA[15]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 302.835 0 303.035 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 302.835 0 303.035 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 302.835 0 303.035 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END BWENA[15]

 PIN BWENB[15]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 304.615 0 304.815 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 304.615 0 304.815 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 304.615 0 304.815 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END BWENB[15]

 PIN DB[15]
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 306.295 0 306.495 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 306.295 0 306.495 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 306.295 0 306.495 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END DB[15]

 PIN QB[15]
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M3 ;
 RECT 309.155 0 309.355 0.48 ;
 END
 PORT
 LAYER M2 ;
 RECT 309.155 0 309.355 0.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 309.155 0 309.355 0.48 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ;
 END QB[15]

 PIN VDD
 USE POWER ;
  
 PORT
 LAYER M4 ;
 POLYGON 120.83 35.015 122.03 35.015 122.03 0 120.83 0 ;
 POLYGON 120.83 35.015 122.03 35.015 122.03 319.25 120.83 319.25 ;
 END
 PORT
 LAYER M4 ;
 POLYGON 192.69 35.015 191.49 35.015 191.49 0 192.69 0 ;
 POLYGON 192.69 35.015 191.49 35.015 191.49 319.25 192.69 319.25 ;
 END   
 PORT
 LAYER M4 ;
 POLYGON 105.55 35.015 106.75 35.015 106.75 0 105.55 0 ;
 POLYGON 105.55 35.015 106.75 35.015 106.75 319.25 105.55 319.25 ;
 END
 PORT
 LAYER M4 ;
 POLYGON 207.97 35.015 206.77 35.015 206.77 0 207.97 0 ;
 POLYGON 207.97 35.015 206.77 35.015 206.77 319.25 207.97 319.25 ;
 END   
 PORT
 LAYER M4 ;
 POLYGON 90.27 35.015 91.47 35.015 91.47 0 90.27 0 ;
 POLYGON 90.27 35.015 91.47 35.015 91.47 319.25 90.27 319.25 ;
 END
 PORT
 LAYER M4 ;
 POLYGON 223.25 35.015 222.05 35.015 222.05 0 223.25 0 ;
 POLYGON 223.25 35.015 222.05 35.015 222.05 319.25 223.25 319.25 ;
 END   
 PORT
 LAYER M4 ;
 POLYGON 74.99 35.015 76.19 35.015 76.19 0 74.99 0 ;
 POLYGON 74.99 35.015 76.19 35.015 76.19 319.25 74.99 319.25 ;
 END
 PORT
 LAYER M4 ;
 POLYGON 238.53 35.015 237.33 35.015 237.33 0 238.53 0 ;
 POLYGON 238.53 35.015 237.33 35.015 237.33 319.25 238.53 319.25 ;
 END   
 PORT
 LAYER M4 ;
 POLYGON 59.71 35.015 60.91 35.015 60.91 0 59.71 0 ;
 POLYGON 59.71 35.015 60.91 35.015 60.91 319.25 59.71 319.25 ;
 END
 PORT
 LAYER M4 ;
 POLYGON 253.81 35.015 252.61 35.015 252.61 0 253.81 0 ;
 POLYGON 253.81 35.015 252.61 35.015 252.61 319.25 253.81 319.25 ;
 END   
 PORT
 LAYER M4 ;
 POLYGON 44.43 35.015 45.63 35.015 45.63 0 44.43 0 ;
 POLYGON 44.43 35.015 45.63 35.015 45.63 319.25 44.43 319.25 ;
 END
 PORT
 LAYER M4 ;
 POLYGON 269.09 35.015 267.89 35.015 267.89 0 269.09 0 ;
 POLYGON 269.09 35.015 267.89 35.015 267.89 319.25 269.09 319.25 ;
 END   
 PORT
 LAYER M4 ;
 POLYGON 29.15 35.015 30.35 35.015 30.35 0 29.15 0 ;
 POLYGON 29.15 35.015 30.35 35.015 30.35 319.25 29.15 319.25 ;
 END
 PORT
 LAYER M4 ;
 POLYGON 284.37 35.015 283.17 35.015 283.17 0 284.37 0 ;
 POLYGON 284.37 35.015 283.17 35.015 283.17 319.25 284.37 319.25 ;
 END   
 PORT
 LAYER M4 ;
 POLYGON 13.87 35.015 15.07 35.015 15.07 0 13.87 0 ;
 POLYGON 13.87 35.015 15.07 35.015 15.07 319.25 13.87 319.25 ;
 END
 PORT
 LAYER M4 ;
 POLYGON 299.65 35.015 298.45 35.015 298.45 0 299.65 0 ;
 POLYGON 299.65 35.015 298.45 35.015 298.45 319.25 299.65 319.25 ;
 END   
  
 PORT
 LAYER M4 ;
 POLYGON 118.31 15.245 117.83 15.245 117.83 30.99 118.31 30.99 118.31 35.015 117.01 35.015 117.01 0 118.31 0 ;
 POLYGON 118.31 35.015 117.01 35.015 117.01 319.25 118.31 319.25 ;
 END
 PORT
 LAYER M4 ;
 POLYGON 195.21 15.245 195.69 15.245 195.69 30.99 195.21 30.99 195.21 35.015 196.51 35.015 196.51 0 195.21 0 ;
 POLYGON 195.21 35.015 196.51 35.015 196.51 319.25 195.21 319.25 ;
 END   
 PORT
 LAYER M4 ;
 POLYGON 103.03 15.245 102.55 15.245 102.55 30.99 103.03 30.99 103.03 35.015 101.73 35.015 101.73 0 103.03 0 ;
 POLYGON 103.03 35.015 101.73 35.015 101.73 319.25 103.03 319.25 ;
 END
 PORT
 LAYER M4 ;
 POLYGON 210.49 15.245 210.97 15.245 210.97 30.99 210.49 30.99 210.49 35.015 211.79 35.015 211.79 0 210.49 0 ;
 POLYGON 210.49 35.015 211.79 35.015 211.79 319.25 210.49 319.25 ;
 END   
 PORT
 LAYER M4 ;
 POLYGON 87.75 15.245 87.27 15.245 87.27 30.99 87.75 30.99 87.75 35.015 86.45 35.015 86.45 0 87.75 0 ;
 POLYGON 87.75 35.015 86.45 35.015 86.45 319.25 87.75 319.25 ;
 END
 PORT
 LAYER M4 ;
 POLYGON 225.77 15.245 226.25 15.245 226.25 30.99 225.77 30.99 225.77 35.015 227.07 35.015 227.07 0 225.77 0 ;
 POLYGON 225.77 35.015 227.07 35.015 227.07 319.25 225.77 319.25 ;
 END   
 PORT
 LAYER M4 ;
 POLYGON 72.47 15.245 71.99 15.245 71.99 30.99 72.47 30.99 72.47 35.015 71.17 35.015 71.17 0 72.47 0 ;
 POLYGON 72.47 35.015 71.17 35.015 71.17 319.25 72.47 319.25 ;
 END
 PORT
 LAYER M4 ;
 POLYGON 241.05 15.245 241.53 15.245 241.53 30.99 241.05 30.99 241.05 35.015 242.35 35.015 242.35 0 241.05 0 ;
 POLYGON 241.05 35.015 242.35 35.015 242.35 319.25 241.05 319.25 ;
 END   
 PORT
 LAYER M4 ;
 POLYGON 57.19 15.245 56.71 15.245 56.71 30.99 57.19 30.99 57.19 35.015 55.89 35.015 55.89 0 57.19 0 ;
 POLYGON 57.19 35.015 55.89 35.015 55.89 319.25 57.19 319.25 ;
 END
 PORT
 LAYER M4 ;
 POLYGON 256.33 15.245 256.81 15.245 256.81 30.99 256.33 30.99 256.33 35.015 257.63 35.015 257.63 0 256.33 0 ;
 POLYGON 256.33 35.015 257.63 35.015 257.63 319.25 256.33 319.25 ;
 END   
 PORT
 LAYER M4 ;
 POLYGON 41.91 15.245 41.43 15.245 41.43 30.99 41.91 30.99 41.91 35.015 40.61 35.015 40.61 0 41.91 0 ;
 POLYGON 41.91 35.015 40.61 35.015 40.61 319.25 41.91 319.25 ;
 END
 PORT
 LAYER M4 ;
 POLYGON 271.61 15.245 272.09 15.245 272.09 30.99 271.61 30.99 271.61 35.015 272.91 35.015 272.91 0 271.61 0 ;
 POLYGON 271.61 35.015 272.91 35.015 272.91 319.25 271.61 319.25 ;
 END   
 PORT
 LAYER M4 ;
 POLYGON 26.63 15.245 26.15 15.245 26.15 30.99 26.63 30.99 26.63 35.015 25.33 35.015 25.33 0 26.63 0 ;
 POLYGON 26.63 35.015 25.33 35.015 25.33 319.25 26.63 319.25 ;
 END
 PORT
 LAYER M4 ;
 POLYGON 286.89 15.245 287.37 15.245 287.37 30.99 286.89 30.99 286.89 35.015 288.19 35.015 288.19 0 286.89 0 ;
 POLYGON 286.89 35.015 288.19 35.015 288.19 319.25 286.89 319.25 ;
 END   
 PORT
 LAYER M4 ;
 POLYGON 11.35 15.245 10.87 15.245 10.87 30.99 11.35 30.99 11.35 35.015 10.05 35.015 10.05 0 11.35 0 ;
 POLYGON 11.35 35.015 10.05 35.015 10.05 319.25 11.35 319.25 ;
 END
 PORT
 LAYER M4 ;
 POLYGON 302.17 15.245 302.65 15.245 302.65 30.99 302.17 30.99 302.17 35.015 303.47 35.015 303.47 0 302.17 0 ;
 POLYGON 302.17 35.015 303.47 35.015 303.47 319.25 302.17 319.25 ;
 END   
  
 PORT
 LAYER M4 ;
 POLYGON 114.49 15.245 114.01 15.245 114.01 29.56 114.49 29.56 114.49 35.015 113.19 35.015 113.19 0 114.49 0 ;
 POLYGON 114.49 35.015 113.19 35.015 113.19 319.25 114.49 319.25 ;
 END
 PORT
 LAYER M4 ;
 POLYGON 199.03 15.245 199.51 15.245 199.51 29.56 199.03 29.56 199.03 35.015 200.33 35.015 200.33 0 199.03 0 ;
 POLYGON 199.03 35.015 200.33 35.015 200.33 319.25 199.03 319.25 ;
 END   
 PORT
 LAYER M4 ;
 POLYGON 99.21 15.245 98.73 15.245 98.73 29.56 99.21 29.56 99.21 35.015 97.91 35.015 97.91 0 99.21 0 ;
 POLYGON 99.21 35.015 97.91 35.015 97.91 319.25 99.21 319.25 ;
 END
 PORT
 LAYER M4 ;
 POLYGON 214.31 15.245 214.79 15.245 214.79 29.56 214.31 29.56 214.31 35.015 215.61 35.015 215.61 0 214.31 0 ;
 POLYGON 214.31 35.015 215.61 35.015 215.61 319.25 214.31 319.25 ;
 END   
 PORT
 LAYER M4 ;
 POLYGON 83.93 15.245 83.45 15.245 83.45 29.56 83.93 29.56 83.93 35.015 82.63 35.015 82.63 0 83.93 0 ;
 POLYGON 83.93 35.015 82.63 35.015 82.63 319.25 83.93 319.25 ;
 END
 PORT
 LAYER M4 ;
 POLYGON 229.59 15.245 230.07 15.245 230.07 29.56 229.59 29.56 229.59 35.015 230.89 35.015 230.89 0 229.59 0 ;
 POLYGON 229.59 35.015 230.89 35.015 230.89 319.25 229.59 319.25 ;
 END   
 PORT
 LAYER M4 ;
 POLYGON 68.65 15.245 68.17 15.245 68.17 29.56 68.65 29.56 68.65 35.015 67.35 35.015 67.35 0 68.65 0 ;
 POLYGON 68.65 35.015 67.35 35.015 67.35 319.25 68.65 319.25 ;
 END
 PORT
 LAYER M4 ;
 POLYGON 244.87 15.245 245.35 15.245 245.35 29.56 244.87 29.56 244.87 35.015 246.17 35.015 246.17 0 244.87 0 ;
 POLYGON 244.87 35.015 246.17 35.015 246.17 319.25 244.87 319.25 ;
 END   
 PORT
 LAYER M4 ;
 POLYGON 53.37 15.245 52.89 15.245 52.89 29.56 53.37 29.56 53.37 35.015 52.07 35.015 52.07 0 53.37 0 ;
 POLYGON 53.37 35.015 52.07 35.015 52.07 319.25 53.37 319.25 ;
 END
 PORT
 LAYER M4 ;
 POLYGON 260.15 15.245 260.63 15.245 260.63 29.56 260.15 29.56 260.15 35.015 261.45 35.015 261.45 0 260.15 0 ;
 POLYGON 260.15 35.015 261.45 35.015 261.45 319.25 260.15 319.25 ;
 END   
 PORT
 LAYER M4 ;
 POLYGON 38.09 15.245 37.61 15.245 37.61 29.56 38.09 29.56 38.09 35.015 36.79 35.015 36.79 0 38.09 0 ;
 POLYGON 38.09 35.015 36.79 35.015 36.79 319.25 38.09 319.25 ;
 END
 PORT
 LAYER M4 ;
 POLYGON 275.43 15.245 275.91 15.245 275.91 29.56 275.43 29.56 275.43 35.015 276.73 35.015 276.73 0 275.43 0 ;
 POLYGON 275.43 35.015 276.73 35.015 276.73 319.25 275.43 319.25 ;
 END   
 PORT
 LAYER M4 ;
 POLYGON 22.81 15.245 22.33 15.245 22.33 29.56 22.81 29.56 22.81 35.015 21.51 35.015 21.51 0 22.81 0 ;
 POLYGON 22.81 35.015 21.51 35.015 21.51 319.25 22.81 319.25 ;
 END
 PORT
 LAYER M4 ;
 POLYGON 290.71 15.245 291.19 15.245 291.19 29.56 290.71 29.56 290.71 35.015 292.01 35.015 292.01 0 290.71 0 ;
 POLYGON 290.71 35.015 292.01 35.015 292.01 319.25 290.71 319.25 ;
 END   
 PORT
 LAYER M4 ;
 POLYGON 7.53 15.245 7.05 15.245 7.05 29.56 7.53 29.56 7.53 35.015 6.23 35.015 6.23 0 7.53 0 ;
 POLYGON 7.53 35.015 6.23 35.015 6.23 319.25 7.53 319.25 ;
 END
 PORT
 LAYER M4 ;
 POLYGON 305.99 15.245 306.47 15.245 306.47 29.56 305.99 29.56 305.99 35.015 307.29 35.015 307.29 0 305.99 0 ;
 POLYGON 305.99 35.015 307.29 35.015 307.29 319.25 305.99 319.25 ;
 END   
  
 PORT
 LAYER M4 ;
 POLYGON 109.37 35.015 110.57 35.015 110.57 0 109.37 0 ;
 POLYGON 109.37 35.015 110.57 35.015 110.57 319.25 109.37 319.25 ;
 END
 PORT
 LAYER M4 ;
 POLYGON 204.15 35.015 202.95 35.015 202.95 0 204.15 0 ;
 POLYGON 204.15 35.015 202.95 35.015 202.95 319.25 204.15 319.25 ;
 END   
 PORT
 LAYER M4 ;
 POLYGON 94.09 35.015 95.29 35.015 95.29 0 94.09 0 ;
 POLYGON 94.09 35.015 95.29 35.015 95.29 319.25 94.09 319.25 ;
 END
 PORT
 LAYER M4 ;
 POLYGON 219.43 35.015 218.23 35.015 218.23 0 219.43 0 ;
 POLYGON 219.43 35.015 218.23 35.015 218.23 319.25 219.43 319.25 ;
 END   
 PORT
 LAYER M4 ;
 POLYGON 78.81 35.015 80.01 35.015 80.01 0 78.81 0 ;
 POLYGON 78.81 35.015 80.01 35.015 80.01 319.25 78.81 319.25 ;
 END
 PORT
 LAYER M4 ;
 POLYGON 234.71 35.015 233.51 35.015 233.51 0 234.71 0 ;
 POLYGON 234.71 35.015 233.51 35.015 233.51 319.25 234.71 319.25 ;
 END   
 PORT
 LAYER M4 ;
 POLYGON 63.53 35.015 64.73 35.015 64.73 0 63.53 0 ;
 POLYGON 63.53 35.015 64.73 35.015 64.73 319.25 63.53 319.25 ;
 END
 PORT
 LAYER M4 ;
 POLYGON 249.99 35.015 248.79 35.015 248.79 0 249.99 0 ;
 POLYGON 249.99 35.015 248.79 35.015 248.79 319.25 249.99 319.25 ;
 END   
 PORT
 LAYER M4 ;
 POLYGON 48.25 35.015 49.45 35.015 49.45 0 48.25 0 ;
 POLYGON 48.25 35.015 49.45 35.015 49.45 319.25 48.25 319.25 ;
 END
 PORT
 LAYER M4 ;
 POLYGON 265.27 35.015 264.07 35.015 264.07 0 265.27 0 ;
 POLYGON 265.27 35.015 264.07 35.015 264.07 319.25 265.27 319.25 ;
 END   
 PORT
 LAYER M4 ;
 POLYGON 32.97 35.015 34.17 35.015 34.17 0 32.97 0 ;
 POLYGON 32.97 35.015 34.17 35.015 34.17 319.25 32.97 319.25 ;
 END
 PORT
 LAYER M4 ;
 POLYGON 280.55 35.015 279.35 35.015 279.35 0 280.55 0 ;
 POLYGON 280.55 35.015 279.35 35.015 279.35 319.25 280.55 319.25 ;
 END   
 PORT
 LAYER M4 ;
 POLYGON 17.69 35.015 18.89 35.015 18.89 0 17.69 0 ;
 POLYGON 17.69 35.015 18.89 35.015 18.89 319.25 17.69 319.25 ;
 END
 PORT
 LAYER M4 ;
 POLYGON 295.83 35.015 294.63 35.015 294.63 0 295.83 0 ;
 POLYGON 295.83 35.015 294.63 35.015 294.63 319.25 295.83 319.25 ;
 END   
 PORT
 LAYER M4 ;
 POLYGON 2.41 35.015 3.61 35.015 3.61 0 2.41 0 ;
 POLYGON 2.41 35.015 3.61 35.015 3.61 319.25 2.41 319.25 ;
 END
 PORT
 LAYER M4 ;
 POLYGON 311.11 35.015 309.91 35.015 309.91 0 311.11 0 ;
 POLYGON 311.11 35.015 309.91 35.015 309.91 319.25 311.11 319.25 ;
 END   
 PORT
 LAYER M4 ;
 RECT 127.325 0 129.325 319.25 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 132.825 0 134.825 319.25 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 139.575 0 141.575 319.25 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 145.575 0 147.575 319.25 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 150.575 0 152.575 319.25 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 160.945 0 162.945 319.25 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 165.945 0 167.945 319.25 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 171.945 0 173.945 319.25 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 178.695 0 180.695 319.25 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 184.195 0 186.195 319.25 ;    
 END 
 END VDD

 PIN VSS
 USE GROUND ;
  
 PORT
 LAYER M4 ;
 POLYGON 122.74 35.015 123.94 35.015 123.94 0 122.74 0 ;
 POLYGON 122.74 35.015 123.94 35.015 123.94 319.25 122.74 319.25 ;
 END
 PORT
 LAYER M4 ;
 POLYGON 190.78 35.015 189.58 35.015 189.58 0 190.78 0 ;
 POLYGON 190.78 35.015 189.58 35.015 189.58 319.25 190.78 319.25 ;
 END   
 PORT
 LAYER M4 ;
 POLYGON 107.46 35.015 108.66 35.015 108.66 0 107.46 0 ;
 POLYGON 107.46 35.015 108.66 35.015 108.66 319.25 107.46 319.25 ;
 END
 PORT
 LAYER M4 ;
 POLYGON 206.06 35.015 204.86 35.015 204.86 0 206.06 0 ;
 POLYGON 206.06 35.015 204.86 35.015 204.86 319.25 206.06 319.25 ;
 END   
 PORT
 LAYER M4 ;
 POLYGON 92.18 35.015 93.38 35.015 93.38 0 92.18 0 ;
 POLYGON 92.18 35.015 93.38 35.015 93.38 319.25 92.18 319.25 ;
 END
 PORT
 LAYER M4 ;
 POLYGON 221.34 35.015 220.14 35.015 220.14 0 221.34 0 ;
 POLYGON 221.34 35.015 220.14 35.015 220.14 319.25 221.34 319.25 ;
 END   
 PORT
 LAYER M4 ;
 POLYGON 76.9 35.015 78.1 35.015 78.1 0 76.9 0 ;
 POLYGON 76.9 35.015 78.1 35.015 78.1 319.25 76.9 319.25 ;
 END
 PORT
 LAYER M4 ;
 POLYGON 236.62 35.015 235.42 35.015 235.42 0 236.62 0 ;
 POLYGON 236.62 35.015 235.42 35.015 235.42 319.25 236.62 319.25 ;
 END   
 PORT
 LAYER M4 ;
 POLYGON 61.62 35.015 62.82 35.015 62.82 0 61.62 0 ;
 POLYGON 61.62 35.015 62.82 35.015 62.82 319.25 61.62 319.25 ;
 END
 PORT
 LAYER M4 ;
 POLYGON 251.9 35.015 250.7 35.015 250.7 0 251.9 0 ;
 POLYGON 251.9 35.015 250.7 35.015 250.7 319.25 251.9 319.25 ;
 END   
 PORT
 LAYER M4 ;
 POLYGON 46.34 35.015 47.54 35.015 47.54 0 46.34 0 ;
 POLYGON 46.34 35.015 47.54 35.015 47.54 319.25 46.34 319.25 ;
 END
 PORT
 LAYER M4 ;
 POLYGON 267.18 35.015 265.98 35.015 265.98 0 267.18 0 ;
 POLYGON 267.18 35.015 265.98 35.015 265.98 319.25 267.18 319.25 ;
 END   
 PORT
 LAYER M4 ;
 POLYGON 31.06 35.015 32.26 35.015 32.26 0 31.06 0 ;
 POLYGON 31.06 35.015 32.26 35.015 32.26 319.25 31.06 319.25 ;
 END
 PORT
 LAYER M4 ;
 POLYGON 282.46 35.015 281.26 35.015 281.26 0 282.46 0 ;
 POLYGON 282.46 35.015 281.26 35.015 281.26 319.25 282.46 319.25 ;
 END   
 PORT
 LAYER M4 ;
 POLYGON 15.78 35.015 16.98 35.015 16.98 0 15.78 0 ;
 POLYGON 15.78 35.015 16.98 35.015 16.98 319.25 15.78 319.25 ;
 END
 PORT
 LAYER M4 ;
 POLYGON 297.74 35.015 296.54 35.015 296.54 0 297.74 0 ;
 POLYGON 297.74 35.015 296.54 35.015 296.54 319.25 297.74 319.25 ;
 END   
  
 PORT
 LAYER M4 ;
 POLYGON 118.82 15.245 119.3 15.245 119.3 30.99 118.82 30.99 118.82 35.015 120.12 35.015 120.12 0 118.82 0 ;
 POLYGON 118.82 35.015 120.12 35.015 120.12 319.25 118.82 319.25 ;
 END
 PORT
 LAYER M4 ;
 POLYGON 194.7 15.245 194.22 15.245 194.22 30.99 194.7 30.99 194.7 35.015 193.4 35.015 193.4 0 194.7 0 ;
 POLYGON 194.7 35.015 193.4 35.015 193.4 319.25 194.7 319.25 ;
 END   
 PORT
 LAYER M4 ;
 POLYGON 103.54 15.245 104.02 15.245 104.02 30.99 103.54 30.99 103.54 35.015 104.84 35.015 104.84 0 103.54 0 ;
 POLYGON 103.54 35.015 104.84 35.015 104.84 319.25 103.54 319.25 ;
 END
 PORT
 LAYER M4 ;
 POLYGON 209.98 15.245 209.5 15.245 209.5 30.99 209.98 30.99 209.98 35.015 208.68 35.015 208.68 0 209.98 0 ;
 POLYGON 209.98 35.015 208.68 35.015 208.68 319.25 209.98 319.25 ;
 END   
 PORT
 LAYER M4 ;
 POLYGON 88.26 15.245 88.74 15.245 88.74 30.99 88.26 30.99 88.26 35.015 89.56 35.015 89.56 0 88.26 0 ;
 POLYGON 88.26 35.015 89.56 35.015 89.56 319.25 88.26 319.25 ;
 END
 PORT
 LAYER M4 ;
 POLYGON 225.26 15.245 224.78 15.245 224.78 30.99 225.26 30.99 225.26 35.015 223.96 35.015 223.96 0 225.26 0 ;
 POLYGON 225.26 35.015 223.96 35.015 223.96 319.25 225.26 319.25 ;
 END   
 PORT
 LAYER M4 ;
 POLYGON 72.98 15.245 73.46 15.245 73.46 30.99 72.98 30.99 72.98 35.015 74.28 35.015 74.28 0 72.98 0 ;
 POLYGON 72.98 35.015 74.28 35.015 74.28 319.25 72.98 319.25 ;
 END
 PORT
 LAYER M4 ;
 POLYGON 240.54 15.245 240.06 15.245 240.06 30.99 240.54 30.99 240.54 35.015 239.24 35.015 239.24 0 240.54 0 ;
 POLYGON 240.54 35.015 239.24 35.015 239.24 319.25 240.54 319.25 ;
 END   
 PORT
 LAYER M4 ;
 POLYGON 57.7 15.245 58.18 15.245 58.18 30.99 57.7 30.99 57.7 35.015 59 35.015 59 0 57.7 0 ;
 POLYGON 57.7 35.015 59 35.015 59 319.25 57.7 319.25 ;
 END
 PORT
 LAYER M4 ;
 POLYGON 255.82 15.245 255.34 15.245 255.34 30.99 255.82 30.99 255.82 35.015 254.52 35.015 254.52 0 255.82 0 ;
 POLYGON 255.82 35.015 254.52 35.015 254.52 319.25 255.82 319.25 ;
 END   
 PORT
 LAYER M4 ;
 POLYGON 42.42 15.245 42.9 15.245 42.9 30.99 42.42 30.99 42.42 35.015 43.72 35.015 43.72 0 42.42 0 ;
 POLYGON 42.42 35.015 43.72 35.015 43.72 319.25 42.42 319.25 ;
 END
 PORT
 LAYER M4 ;
 POLYGON 271.1 15.245 270.62 15.245 270.62 30.99 271.1 30.99 271.1 35.015 269.8 35.015 269.8 0 271.1 0 ;
 POLYGON 271.1 35.015 269.8 35.015 269.8 319.25 271.1 319.25 ;
 END   
 PORT
 LAYER M4 ;
 POLYGON 27.14 15.245 27.62 15.245 27.62 30.99 27.14 30.99 27.14 35.015 28.44 35.015 28.44 0 27.14 0 ;
 POLYGON 27.14 35.015 28.44 35.015 28.44 319.25 27.14 319.25 ;
 END
 PORT
 LAYER M4 ;
 POLYGON 286.38 15.245 285.9 15.245 285.9 30.99 286.38 30.99 286.38 35.015 285.08 35.015 285.08 0 286.38 0 ;
 POLYGON 286.38 35.015 285.08 35.015 285.08 319.25 286.38 319.25 ;
 END   
 PORT
 LAYER M4 ;
 POLYGON 11.86 15.245 12.34 15.245 12.34 30.99 11.86 30.99 11.86 35.015 13.16 35.015 13.16 0 11.86 0 ;
 POLYGON 11.86 35.015 13.16 35.015 13.16 319.25 11.86 319.25 ;
 END
 PORT
 LAYER M4 ;
 POLYGON 301.66 15.245 301.18 15.245 301.18 30.99 301.66 30.99 301.66 35.015 300.36 35.015 300.36 0 301.66 0 ;
 POLYGON 301.66 35.015 300.36 35.015 300.36 319.25 301.66 319.25 ;
 END   
  
 PORT
 LAYER M4 ;
 POLYGON 115 15.245 115.48 15.245 115.48 29.56 115 29.56 115 35.015 116.3 35.015 116.3 0 115 0 ;
 POLYGON 115 35.015 116.3 35.015 116.3 319.25 115 319.25 ;
 END
 PORT
 LAYER M4 ;
 POLYGON 198.52 15.245 198.04 15.245 198.04 29.56 198.52 29.56 198.52 35.015 197.22 35.015 197.22 0 198.52 0 ;
 POLYGON 198.52 35.015 197.22 35.015 197.22 319.25 198.52 319.25 ;
 END   
 PORT
 LAYER M4 ;
 POLYGON 99.72 15.245 100.2 15.245 100.2 29.56 99.72 29.56 99.72 35.015 101.02 35.015 101.02 0 99.72 0 ;
 POLYGON 99.72 35.015 101.02 35.015 101.02 319.25 99.72 319.25 ;
 END
 PORT
 LAYER M4 ;
 POLYGON 213.8 15.245 213.32 15.245 213.32 29.56 213.8 29.56 213.8 35.015 212.5 35.015 212.5 0 213.8 0 ;
 POLYGON 213.8 35.015 212.5 35.015 212.5 319.25 213.8 319.25 ;
 END   
 PORT
 LAYER M4 ;
 POLYGON 84.44 15.245 84.92 15.245 84.92 29.56 84.44 29.56 84.44 35.015 85.74 35.015 85.74 0 84.44 0 ;
 POLYGON 84.44 35.015 85.74 35.015 85.74 319.25 84.44 319.25 ;
 END
 PORT
 LAYER M4 ;
 POLYGON 229.08 15.245 228.6 15.245 228.6 29.56 229.08 29.56 229.08 35.015 227.78 35.015 227.78 0 229.08 0 ;
 POLYGON 229.08 35.015 227.78 35.015 227.78 319.25 229.08 319.25 ;
 END   
 PORT
 LAYER M4 ;
 POLYGON 69.16 15.245 69.64 15.245 69.64 29.56 69.16 29.56 69.16 35.015 70.46 35.015 70.46 0 69.16 0 ;
 POLYGON 69.16 35.015 70.46 35.015 70.46 319.25 69.16 319.25 ;
 END
 PORT
 LAYER M4 ;
 POLYGON 244.36 15.245 243.88 15.245 243.88 29.56 244.36 29.56 244.36 35.015 243.06 35.015 243.06 0 244.36 0 ;
 POLYGON 244.36 35.015 243.06 35.015 243.06 319.25 244.36 319.25 ;
 END   
 PORT
 LAYER M4 ;
 POLYGON 53.88 15.245 54.36 15.245 54.36 29.56 53.88 29.56 53.88 35.015 55.18 35.015 55.18 0 53.88 0 ;
 POLYGON 53.88 35.015 55.18 35.015 55.18 319.25 53.88 319.25 ;
 END
 PORT
 LAYER M4 ;
 POLYGON 259.64 15.245 259.16 15.245 259.16 29.56 259.64 29.56 259.64 35.015 258.34 35.015 258.34 0 259.64 0 ;
 POLYGON 259.64 35.015 258.34 35.015 258.34 319.25 259.64 319.25 ;
 END   
 PORT
 LAYER M4 ;
 POLYGON 38.6 15.245 39.08 15.245 39.08 29.56 38.6 29.56 38.6 35.015 39.9 35.015 39.9 0 38.6 0 ;
 POLYGON 38.6 35.015 39.9 35.015 39.9 319.25 38.6 319.25 ;
 END
 PORT
 LAYER M4 ;
 POLYGON 274.92 15.245 274.44 15.245 274.44 29.56 274.92 29.56 274.92 35.015 273.62 35.015 273.62 0 274.92 0 ;
 POLYGON 274.92 35.015 273.62 35.015 273.62 319.25 274.92 319.25 ;
 END   
 PORT
 LAYER M4 ;
 POLYGON 23.32 15.245 23.8 15.245 23.8 29.56 23.32 29.56 23.32 35.015 24.62 35.015 24.62 0 23.32 0 ;
 POLYGON 23.32 35.015 24.62 35.015 24.62 319.25 23.32 319.25 ;
 END
 PORT
 LAYER M4 ;
 POLYGON 290.2 15.245 289.72 15.245 289.72 29.56 290.2 29.56 290.2 35.015 288.9 35.015 288.9 0 290.2 0 ;
 POLYGON 290.2 35.015 288.9 35.015 288.9 319.25 290.2 319.25 ;
 END   
 PORT
 LAYER M4 ;
 POLYGON 8.04 15.245 8.52 15.245 8.52 29.56 8.04 29.56 8.04 35.015 9.34 35.015 9.34 0 8.04 0 ;
 POLYGON 8.04 35.015 9.34 35.015 9.34 319.25 8.04 319.25 ;
 END
 PORT
 LAYER M4 ;
 POLYGON 305.48 15.245 305 15.245 305 29.56 305.48 29.56 305.48 35.015 304.18 35.015 304.18 0 305.48 0 ;
 POLYGON 305.48 35.015 304.18 35.015 304.18 319.25 305.48 319.25 ;
 END   
  
 PORT
 LAYER M4 ;
 POLYGON 111.28 35.015 112.48 35.015 112.48 0 111.28 0 ;
 POLYGON 111.28 35.015 112.48 35.015 112.48 319.25 111.28 319.25 ;
 END
 PORT
 LAYER M4 ;
 POLYGON 202.24 35.015 201.04 35.015 201.04 0 202.24 0 ;
 POLYGON 202.24 35.015 201.04 35.015 201.04 319.25 202.24 319.25 ;
 END   
 PORT
 LAYER M4 ;
 POLYGON 96 35.015 97.2 35.015 97.2 0 96 0 ;
 POLYGON 96 35.015 97.2 35.015 97.2 319.25 96 319.25 ;
 END
 PORT
 LAYER M4 ;
 POLYGON 217.52 35.015 216.32 35.015 216.32 0 217.52 0 ;
 POLYGON 217.52 35.015 216.32 35.015 216.32 319.25 217.52 319.25 ;
 END   
 PORT
 LAYER M4 ;
 POLYGON 80.72 35.015 81.92 35.015 81.92 0 80.72 0 ;
 POLYGON 80.72 35.015 81.92 35.015 81.92 319.25 80.72 319.25 ;
 END
 PORT
 LAYER M4 ;
 POLYGON 232.8 35.015 231.6 35.015 231.6 0 232.8 0 ;
 POLYGON 232.8 35.015 231.6 35.015 231.6 319.25 232.8 319.25 ;
 END   
 PORT
 LAYER M4 ;
 POLYGON 65.44 35.015 66.64 35.015 66.64 0 65.44 0 ;
 POLYGON 65.44 35.015 66.64 35.015 66.64 319.25 65.44 319.25 ;
 END
 PORT
 LAYER M4 ;
 POLYGON 248.08 35.015 246.88 35.015 246.88 0 248.08 0 ;
 POLYGON 248.08 35.015 246.88 35.015 246.88 319.25 248.08 319.25 ;
 END   
 PORT
 LAYER M4 ;
 POLYGON 50.16 35.015 51.36 35.015 51.36 0 50.16 0 ;
 POLYGON 50.16 35.015 51.36 35.015 51.36 319.25 50.16 319.25 ;
 END
 PORT
 LAYER M4 ;
 POLYGON 263.36 35.015 262.16 35.015 262.16 0 263.36 0 ;
 POLYGON 263.36 35.015 262.16 35.015 262.16 319.25 263.36 319.25 ;
 END   
 PORT
 LAYER M4 ;
 POLYGON 34.88 35.015 36.08 35.015 36.08 0 34.88 0 ;
 POLYGON 34.88 35.015 36.08 35.015 36.08 319.25 34.88 319.25 ;
 END
 PORT
 LAYER M4 ;
 POLYGON 278.64 35.015 277.44 35.015 277.44 0 278.64 0 ;
 POLYGON 278.64 35.015 277.44 35.015 277.44 319.25 278.64 319.25 ;
 END   
 PORT
 LAYER M4 ;
 POLYGON 19.6 35.015 20.8 35.015 20.8 0 19.6 0 ;
 POLYGON 19.6 35.015 20.8 35.015 20.8 319.25 19.6 319.25 ;
 END
 PORT
 LAYER M4 ;
 POLYGON 293.92 35.015 292.72 35.015 292.72 0 293.92 0 ;
 POLYGON 293.92 35.015 292.72 35.015 292.72 319.25 293.92 319.25 ;
 END   
 PORT
 LAYER M4 ;
 POLYGON 4.32 35.015 5.52 35.015 5.52 0 4.32 0 ;
 POLYGON 4.32 35.015 5.52 35.015 5.52 319.25 4.32 319.25 ;
 END
 PORT
 LAYER M4 ;
 POLYGON 309.2 35.015 308 35.015 308 0 309.2 0 ;
 POLYGON 309.2 35.015 308 35.015 308 319.25 309.2 319.25 ;
 END   
 PORT
 LAYER M4 ;
 RECT 129.82 0 131.82 319.25 ;      
 END
 PORT
 LAYER M4 ;
 RECT 135.32 0 137.32 319.25 ;      
 END
 PORT
 LAYER M4 ;
 RECT 142.07 0 144.07 319.25 ;      
 END
 PORT
 LAYER M4 ;
 RECT 148.075 0 150.075 319.25 ;      
 END
 PORT
 LAYER M4 ;
 RECT 153.075 0 155.075 319.25 ;      
 END
 PORT
 LAYER M4 ;
 RECT 158.445 0 160.445 319.25 ;      
 END
 PORT
 LAYER M4 ;
 RECT 163.445 0 165.445 319.25 ;      
 END
 PORT
 LAYER M4 ;
 RECT 169.45 0 171.45 319.25 ;      
 END
 PORT
 LAYER M4 ;
 RECT 176.2 0 178.2 319.25 ;      
 END
 PORT
 LAYER M4 ;
 RECT 181.7 0 183.7 319.25 ;      
 END
 END VSS

 OBS
 LAYER M1 SPACING 0.09 ;
 RECT 0 0 4.075 0.57 ;
 RECT 4.455 0 6.935 0.57 ;
 RECT 7.315 0 8.615 0.57 ;
 RECT 8.995 0 10.395 0.57 ;
 RECT 10.775 0 12.075 0.57 ;
 RECT 12.455 0 14.935 0.57 ;
 RECT 15.315 0 19.355 0.57 ;
 RECT 19.735 0 22.215 0.57 ;
 RECT 22.595 0 23.895 0.57 ;
 RECT 24.275 0 25.675 0.57 ;
 RECT 26.055 0 27.355 0.57 ;
 RECT 27.735 0 30.215 0.57 ;
 RECT 30.595 0 34.635 0.57 ;
 RECT 35.015 0 37.495 0.57 ;
 RECT 37.875 0 39.175 0.57 ;
 RECT 39.555 0 40.955 0.57 ;
 RECT 41.335 0 42.635 0.57 ;
 RECT 43.015 0 45.495 0.57 ;
 RECT 45.875 0 49.915 0.57 ;
 RECT 50.295 0 52.775 0.57 ;
 RECT 53.155 0 54.455 0.57 ;
 RECT 54.835 0 56.235 0.57 ;
 RECT 56.615 0 57.915 0.57 ;
 RECT 58.295 0 60.775 0.57 ;
 RECT 61.155 0 65.195 0.57 ;
 RECT 65.575 0 68.055 0.57 ;
 RECT 68.435 0 69.735 0.57 ;
 RECT 70.115 0 71.515 0.57 ;
 RECT 71.895 0 73.195 0.57 ;
 RECT 73.575 0 76.055 0.57 ;
 RECT 76.435 0 80.475 0.57 ;
 RECT 80.855 0 83.335 0.57 ;
 RECT 83.715 0 85.015 0.57 ;
 RECT 85.395 0 86.795 0.57 ;
 RECT 87.175 0 88.475 0.57 ;
 RECT 88.855 0 91.335 0.57 ;
 RECT 91.715 0 95.755 0.57 ;
 RECT 96.135 0 98.615 0.57 ;
 RECT 98.995 0 100.295 0.57 ;
 RECT 100.675 0 102.075 0.57 ;
 RECT 102.455 0 103.755 0.57 ;
 RECT 104.135 0 106.615 0.57 ;
 RECT 106.995 0 111.035 0.57 ;
 RECT 111.415 0 113.895 0.57 ;
 RECT 114.275 0 115.575 0.57 ;
 RECT 115.955 0 117.355 0.57 ;
 RECT 117.735 0 119.035 0.57 ;
 RECT 119.415 0 121.895 0.57 ;
 RECT 122.275 0 126.905 0.57 ;
 RECT 127.285 0 130.07 0.57 ;
 RECT 130.45 0 132.01 0.57 ;
 RECT 132.39 0 137.385 0.57 ;
 RECT 137.765 0 139.98 0.57 ;
 RECT 140.36 0 142.175 0.57 ;
 RECT 142.555 0 143.565 0.57 ;
 RECT 143.945 0 146.17 0.57 ;
 RECT 146.55 0 148.875 0.57 ;
 RECT 149.255 0 150.47 0.57 ;
 RECT 150.85 0 151.345 0.57 ;
 RECT 151.725 0 152.065 0.57 ;
 RECT 152.445 0 152.91 0.57 ;
 RECT 153.29 0 153.775 0.57 ;
 RECT 154.155 0 154.62 0.57 ;
 RECT 155 0 158.52 0.57 ;
 RECT 158.9 0 159.365 0.57 ;
 RECT 159.745 0 160.23 0.57 ;
 RECT 160.61 0 161.075 0.57 ;
 RECT 161.455 0 161.795 0.57 ;
 RECT 162.175 0 162.67 0.57 ;
 RECT 163.05 0 164.265 0.57 ;
 RECT 164.645 0 166.97 0.57 ;
 RECT 167.35 0 169.575 0.57 ;
 RECT 169.955 0 170.965 0.57 ;
 RECT 171.345 0 173.16 0.57 ;
 RECT 173.54 0 175.755 0.57 ;
 RECT 176.135 0 181.13 0.57 ;
 RECT 181.51 0 183.07 0.57 ;
 RECT 183.45 0 186.235 0.57 ;
 RECT 186.615 0 191.245 0.57 ;
 RECT 191.625 0 194.105 0.57 ;
 RECT 194.485 0 195.785 0.57 ;
 RECT 196.165 0 197.565 0.57 ;
 RECT 197.945 0 199.245 0.57 ;
 RECT 199.625 0 202.105 0.57 ;
 RECT 202.485 0 206.525 0.57 ;
 RECT 206.905 0 209.385 0.57 ;
 RECT 209.765 0 211.065 0.57 ;
 RECT 211.445 0 212.845 0.57 ;
 RECT 213.225 0 214.525 0.57 ;
 RECT 214.905 0 217.385 0.57 ;
 RECT 217.765 0 221.805 0.57 ;
 RECT 222.185 0 224.665 0.57 ;
 RECT 225.045 0 226.345 0.57 ;
 RECT 226.725 0 228.125 0.57 ;
 RECT 228.505 0 229.805 0.57 ;
 RECT 230.185 0 232.665 0.57 ;
 RECT 233.045 0 237.085 0.57 ;
 RECT 237.465 0 239.945 0.57 ;
 RECT 240.325 0 241.625 0.57 ;
 RECT 242.005 0 243.405 0.57 ;
 RECT 243.785 0 245.085 0.57 ;
 RECT 245.465 0 247.945 0.57 ;
 RECT 248.325 0 252.365 0.57 ;
 RECT 252.745 0 255.225 0.57 ;
 RECT 255.605 0 256.905 0.57 ;
 RECT 257.285 0 258.685 0.57 ;
 RECT 259.065 0 260.365 0.57 ;
 RECT 260.745 0 263.225 0.57 ;
 RECT 263.605 0 267.645 0.57 ;
 RECT 268.025 0 270.505 0.57 ;
 RECT 270.885 0 272.185 0.57 ;
 RECT 272.565 0 273.965 0.57 ;
 RECT 274.345 0 275.645 0.57 ;
 RECT 276.025 0 278.505 0.57 ;
 RECT 278.885 0 282.925 0.57 ;
 RECT 283.305 0 285.785 0.57 ;
 RECT 286.165 0 287.465 0.57 ;
 RECT 287.845 0 289.245 0.57 ;
 RECT 289.625 0 290.925 0.57 ;
 RECT 291.305 0 293.785 0.57 ;
 RECT 294.165 0 298.205 0.57 ;
 RECT 298.585 0 301.065 0.57 ;
 RECT 301.445 0 302.745 0.57 ;
 RECT 303.125 0 304.525 0.57 ;
 RECT 304.905 0 306.205 0.57 ;
 RECT 306.585 0 309.065 0.57 ;
 RECT 309.445 0 313.52 0.57 ;
 RECT 0 0.57 313.52 319.25 ;
 LAYER M2 SPACING 0.1 ;
 RECT 0 0 4.065 0.58 ;
 RECT 4.465 0 6.925 0.58 ;
 RECT 7.325 0 8.605 0.58 ;
 RECT 9.005 0 10.385 0.58 ;
 RECT 10.785 0 12.065 0.58 ;
 RECT 12.465 0 14.925 0.58 ;
 RECT 15.325 0 19.345 0.58 ;
 RECT 19.745 0 22.205 0.58 ;
 RECT 22.605 0 23.885 0.58 ;
 RECT 24.285 0 25.665 0.58 ;
 RECT 26.065 0 27.345 0.58 ;
 RECT 27.745 0 30.205 0.58 ;
 RECT 30.605 0 34.625 0.58 ;
 RECT 35.025 0 37.485 0.58 ;
 RECT 37.885 0 39.165 0.58 ;
 RECT 39.565 0 40.945 0.58 ;
 RECT 41.345 0 42.625 0.58 ;
 RECT 43.025 0 45.485 0.58 ;
 RECT 45.885 0 49.905 0.58 ;
 RECT 50.305 0 52.765 0.58 ;
 RECT 53.165 0 54.445 0.58 ;
 RECT 54.845 0 56.225 0.58 ;
 RECT 56.625 0 57.905 0.58 ;
 RECT 58.305 0 60.765 0.58 ;
 RECT 61.165 0 65.185 0.58 ;
 RECT 65.585 0 68.045 0.58 ;
 RECT 68.445 0 69.725 0.58 ;
 RECT 70.125 0 71.505 0.58 ;
 RECT 71.905 0 73.185 0.58 ;
 RECT 73.585 0 76.045 0.58 ;
 RECT 76.445 0 80.465 0.58 ;
 RECT 80.865 0 83.325 0.58 ;
 RECT 83.725 0 85.005 0.58 ;
 RECT 85.405 0 86.785 0.58 ;
 RECT 87.185 0 88.465 0.58 ;
 RECT 88.865 0 91.325 0.58 ;
 RECT 91.725 0 95.745 0.58 ;
 RECT 96.145 0 98.605 0.58 ;
 RECT 99.005 0 100.285 0.58 ;
 RECT 100.685 0 102.065 0.58 ;
 RECT 102.465 0 103.745 0.58 ;
 RECT 104.145 0 106.605 0.58 ;
 RECT 107.005 0 111.025 0.58 ;
 RECT 111.425 0 113.885 0.58 ;
 RECT 114.285 0 115.565 0.58 ;
 RECT 115.965 0 117.345 0.58 ;
 RECT 117.745 0 119.025 0.58 ;
 RECT 119.425 0 121.885 0.58 ;
 RECT 122.285 0 126.895 0.58 ;
 RECT 127.295 0 130.06 0.58 ;
 RECT 130.46 0 132 0.58 ;
 RECT 132.4 0 137.375 0.58 ;
 RECT 137.775 0 139.97 0.58 ;
 RECT 140.37 0 142.165 0.58 ;
 RECT 142.565 0 143.555 0.58 ;
 RECT 143.955 0 146.16 0.58 ;
 RECT 146.56 0 148.865 0.58 ;
 RECT 149.265 0 150.46 0.58 ;
 RECT 150.86 0 151.335 0.58 ;
 RECT 151.735 0 152.055 0.58 ;
 RECT 152.455 0 152.9 0.58 ;
 RECT 153.3 0 153.765 0.58 ;
 RECT 154.165 0 154.61 0.58 ;
 RECT 155.01 0 158.51 0.58 ;
 RECT 158.91 0 159.355 0.58 ;
 RECT 159.755 0 160.22 0.58 ;
 RECT 160.62 0 161.065 0.58 ;
 RECT 161.465 0 161.785 0.58 ;
 RECT 162.185 0 162.66 0.58 ;
 RECT 163.06 0 164.255 0.58 ;
 RECT 164.655 0 166.96 0.58 ;
 RECT 167.36 0 169.565 0.58 ;
 RECT 169.965 0 170.955 0.58 ;
 RECT 171.355 0 173.15 0.58 ;
 RECT 173.55 0 175.745 0.58 ;
 RECT 176.145 0 181.12 0.58 ;
 RECT 181.52 0 183.06 0.58 ;
 RECT 183.46 0 186.225 0.58 ;
 RECT 186.625 0 191.235 0.58 ;
 RECT 191.635 0 194.095 0.58 ;
 RECT 194.495 0 195.775 0.58 ;
 RECT 196.175 0 197.555 0.58 ;
 RECT 197.955 0 199.235 0.58 ;
 RECT 199.635 0 202.095 0.58 ;
 RECT 202.495 0 206.515 0.58 ;
 RECT 206.915 0 209.375 0.58 ;
 RECT 209.775 0 211.055 0.58 ;
 RECT 211.455 0 212.835 0.58 ;
 RECT 213.235 0 214.515 0.58 ;
 RECT 214.915 0 217.375 0.58 ;
 RECT 217.775 0 221.795 0.58 ;
 RECT 222.195 0 224.655 0.58 ;
 RECT 225.055 0 226.335 0.58 ;
 RECT 226.735 0 228.115 0.58 ;
 RECT 228.515 0 229.795 0.58 ;
 RECT 230.195 0 232.655 0.58 ;
 RECT 233.055 0 237.075 0.58 ;
 RECT 237.475 0 239.935 0.58 ;
 RECT 240.335 0 241.615 0.58 ;
 RECT 242.015 0 243.395 0.58 ;
 RECT 243.795 0 245.075 0.58 ;
 RECT 245.475 0 247.935 0.58 ;
 RECT 248.335 0 252.355 0.58 ;
 RECT 252.755 0 255.215 0.58 ;
 RECT 255.615 0 256.895 0.58 ;
 RECT 257.295 0 258.675 0.58 ;
 RECT 259.075 0 260.355 0.58 ;
 RECT 260.755 0 263.215 0.58 ;
 RECT 263.615 0 267.635 0.58 ;
 RECT 268.035 0 270.495 0.58 ;
 RECT 270.895 0 272.175 0.58 ;
 RECT 272.575 0 273.955 0.58 ;
 RECT 274.355 0 275.635 0.58 ;
 RECT 276.035 0 278.495 0.58 ;
 RECT 278.895 0 282.915 0.58 ;
 RECT 283.315 0 285.775 0.58 ;
 RECT 286.175 0 287.455 0.58 ;
 RECT 287.855 0 289.235 0.58 ;
 RECT 289.635 0 290.915 0.58 ;
 RECT 291.315 0 293.775 0.58 ;
 RECT 294.175 0 298.195 0.58 ;
 RECT 298.595 0 301.055 0.58 ;
 RECT 301.455 0 302.735 0.58 ;
 RECT 303.135 0 304.515 0.58 ;
 RECT 304.915 0 306.195 0.58 ;
 RECT 306.595 0 309.055 0.58 ;
 RECT 309.455 0 313.52 0.58 ;
 RECT 0 0.58 313.52 319.25 ;
 LAYER M3 SPACING 0.1 ;
 RECT 0 0 4.065 0.58 ;
 RECT 4.465 0 6.925 0.58 ;
 RECT 7.325 0 8.605 0.58 ;
 RECT 9.005 0 10.385 0.58 ;
 RECT 10.785 0 12.065 0.58 ;
 RECT 12.465 0 14.925 0.58 ;
 RECT 15.325 0 19.345 0.58 ;
 RECT 19.745 0 22.205 0.58 ;
 RECT 22.605 0 23.885 0.58 ;
 RECT 24.285 0 25.665 0.58 ;
 RECT 26.065 0 27.345 0.58 ;
 RECT 27.745 0 30.205 0.58 ;
 RECT 30.605 0 34.625 0.58 ;
 RECT 35.025 0 37.485 0.58 ;
 RECT 37.885 0 39.165 0.58 ;
 RECT 39.565 0 40.945 0.58 ;
 RECT 41.345 0 42.625 0.58 ;
 RECT 43.025 0 45.485 0.58 ;
 RECT 45.885 0 49.905 0.58 ;
 RECT 50.305 0 52.765 0.58 ;
 RECT 53.165 0 54.445 0.58 ;
 RECT 54.845 0 56.225 0.58 ;
 RECT 56.625 0 57.905 0.58 ;
 RECT 58.305 0 60.765 0.58 ;
 RECT 61.165 0 65.185 0.58 ;
 RECT 65.585 0 68.045 0.58 ;
 RECT 68.445 0 69.725 0.58 ;
 RECT 70.125 0 71.505 0.58 ;
 RECT 71.905 0 73.185 0.58 ;
 RECT 73.585 0 76.045 0.58 ;
 RECT 76.445 0 80.465 0.58 ;
 RECT 80.865 0 83.325 0.58 ;
 RECT 83.725 0 85.005 0.58 ;
 RECT 85.405 0 86.785 0.58 ;
 RECT 87.185 0 88.465 0.58 ;
 RECT 88.865 0 91.325 0.58 ;
 RECT 91.725 0 95.745 0.58 ;
 RECT 96.145 0 98.605 0.58 ;
 RECT 99.005 0 100.285 0.58 ;
 RECT 100.685 0 102.065 0.58 ;
 RECT 102.465 0 103.745 0.58 ;
 RECT 104.145 0 106.605 0.58 ;
 RECT 107.005 0 111.025 0.58 ;
 RECT 111.425 0 113.885 0.58 ;
 RECT 114.285 0 115.565 0.58 ;
 RECT 115.965 0 117.345 0.58 ;
 RECT 117.745 0 119.025 0.58 ;
 RECT 119.425 0 121.885 0.58 ;
 RECT 122.285 0 126.895 0.58 ;
 RECT 127.295 0 130.06 0.58 ;
 RECT 130.46 0 132 0.58 ;
 RECT 132.4 0 137.375 0.58 ;
 RECT 137.775 0 139.97 0.58 ;
 RECT 140.37 0 142.165 0.58 ;
 RECT 142.565 0 143.555 0.58 ;
 RECT 143.955 0 146.16 0.58 ;
 RECT 146.56 0 148.865 0.58 ;
 RECT 149.265 0 150.46 0.58 ;
 RECT 150.86 0 151.335 0.58 ;
 RECT 151.735 0 152.055 0.58 ;
 RECT 152.455 0 152.9 0.58 ;
 RECT 153.3 0 153.765 0.58 ;
 RECT 154.165 0 154.61 0.58 ;
 RECT 155.01 0 158.51 0.58 ;
 RECT 158.91 0 159.355 0.58 ;
 RECT 159.755 0 160.22 0.58 ;
 RECT 160.62 0 161.065 0.58 ;
 RECT 161.465 0 161.785 0.58 ;
 RECT 162.185 0 162.66 0.58 ;
 RECT 163.06 0 164.255 0.58 ;
 RECT 164.655 0 166.96 0.58 ;
 RECT 167.36 0 169.565 0.58 ;
 RECT 169.965 0 170.955 0.58 ;
 RECT 171.355 0 173.15 0.58 ;
 RECT 173.55 0 175.745 0.58 ;
 RECT 176.145 0 181.12 0.58 ;
 RECT 181.52 0 183.06 0.58 ;
 RECT 183.46 0 186.225 0.58 ;
 RECT 186.625 0 191.235 0.58 ;
 RECT 191.635 0 194.095 0.58 ;
 RECT 194.495 0 195.775 0.58 ;
 RECT 196.175 0 197.555 0.58 ;
 RECT 197.955 0 199.235 0.58 ;
 RECT 199.635 0 202.095 0.58 ;
 RECT 202.495 0 206.515 0.58 ;
 RECT 206.915 0 209.375 0.58 ;
 RECT 209.775 0 211.055 0.58 ;
 RECT 211.455 0 212.835 0.58 ;
 RECT 213.235 0 214.515 0.58 ;
 RECT 214.915 0 217.375 0.58 ;
 RECT 217.775 0 221.795 0.58 ;
 RECT 222.195 0 224.655 0.58 ;
 RECT 225.055 0 226.335 0.58 ;
 RECT 226.735 0 228.115 0.58 ;
 RECT 228.515 0 229.795 0.58 ;
 RECT 230.195 0 232.655 0.58 ;
 RECT 233.055 0 237.075 0.58 ;
 RECT 237.475 0 239.935 0.58 ;
 RECT 240.335 0 241.615 0.58 ;
 RECT 242.015 0 243.395 0.58 ;
 RECT 243.795 0 245.075 0.58 ;
 RECT 245.475 0 247.935 0.58 ;
 RECT 248.335 0 252.355 0.58 ;
 RECT 252.755 0 255.215 0.58 ;
 RECT 255.615 0 256.895 0.58 ;
 RECT 257.295 0 258.675 0.58 ;
 RECT 259.075 0 260.355 0.58 ;
 RECT 260.755 0 263.215 0.58 ;
 RECT 263.615 0 267.635 0.58 ;
 RECT 268.035 0 270.495 0.58 ;
 RECT 270.895 0 272.175 0.58 ;
 RECT 272.575 0 273.955 0.58 ;
 RECT 274.355 0 275.635 0.58 ;
 RECT 276.035 0 278.495 0.58 ;
 RECT 278.895 0 282.915 0.58 ;
 RECT 283.315 0 285.775 0.58 ;
 RECT 286.175 0 287.455 0.58 ;
 RECT 287.855 0 289.235 0.58 ;
 RECT 289.635 0 290.915 0.58 ;
 RECT 291.315 0 293.775 0.58 ;
 RECT 294.175 0 298.195 0.58 ;
 RECT 298.595 0 301.055 0.58 ;
 RECT 301.455 0 302.735 0.58 ;
 RECT 303.135 0 304.515 0.58 ;
 RECT 304.915 0 306.195 0.58 ;
 RECT 306.595 0 309.055 0.58 ;
 RECT 309.455 0 313.52 0.58 ;
 RECT 0 0.58 313.52 319.25 ;

 LAYER V1 ;
 RECT 0 0 313.52 319.25 ;
 LAYER V2 ;
 RECT 0 0 313.52 319.25 ;
 LAYER V3 ;
 RECT 0 0 313.52 319.25 ;

 LAYER M4 SPACING 0.1 ;
 RECT 124.295 0 127.225 0.58 ;
 RECT 124.295 0.58 127.225 319.25 ;
 RECT 129.425 0 129.72 0.58 ;
 RECT 129.425 0.58 129.72 319.25 ;
 RECT 131.92 0 132.725 0.58 ;
 RECT 131.92 0.58 132.725 319.25 ;
 RECT 134.925 0 135.22 0.58 ;
 RECT 134.925 0.58 135.22 319.25 ;
 RECT 137.42 0 139.475 0.58 ;
 RECT 137.42 0.58 139.475 319.25 ;
 RECT 141.675 0 141.97 0.58 ;
 RECT 141.675 0.58 141.97 319.25 ;
 RECT 144.17 0 145.475 0.58 ;
 RECT 144.17 0.58 145.475 319.25 ;
 RECT 147.675 0 147.975 0.58 ;
 RECT 147.675 0.58 147.975 319.25 ;
 RECT 150.175 0 150.475 0.58 ;
 RECT 150.175 0.58 150.475 319.25 ;
 RECT 152.675 0 152.975 0.58 ;
 RECT 152.675 0.58 152.975 319.25 ;
 RECT 155.175 0 158.345 0.58 ;
 RECT 155.175 0.58 158.345 319.25 ;
 RECT 160.545 0 160.845 0.58 ;
 RECT 160.545 0.58 160.845 319.25 ;
 RECT 163.045 0 163.345 0.58 ;
 RECT 163.045 0.58 163.345 319.25 ;
 RECT 165.545 0 165.845 0.58 ;
 RECT 165.545 0.58 165.845 319.25 ;
 RECT 168.045 0 169.35 0.58 ;
 RECT 168.045 0.58 169.35 319.25 ;
 RECT 171.55 0 171.845 0.58 ;
 RECT 171.55 0.58 171.845 319.25 ;
 RECT 174.045 0 176.1 0.58 ;
 RECT 174.045 0.58 176.1 319.25 ;
 RECT 178.3 0 178.595 0.58 ;
 RECT 178.3 0.58 178.595 319.25 ;
 RECT 180.795 0 181.6 0.58 ;
 RECT 180.795 0.58 181.6 319.25 ;
 RECT 183.8 0 184.095 0.58 ;
 RECT 183.8 0.58 184.095 319.25 ;
 RECT 186.295 0 189.48 0.58 ;
 RECT 186.295 0.58 189.48 319.25 ;
 RECT 119.2 15.345 117.93 30.89 ;
 RECT 194.32 15.345 195.59 30.89 ;
 RECT 103.92 15.345 102.65 30.89 ;
 RECT 209.6 15.345 210.87 30.89 ;
 RECT 88.64 15.345 87.37 30.89 ;
 RECT 224.88 15.345 226.15 30.89 ;
 RECT 73.36 15.345 72.09 30.89 ;
 RECT 240.16 15.345 241.43 30.89 ;
 RECT 58.08 15.345 56.81 30.89 ;
 RECT 255.44 15.345 256.71 30.89 ;
 RECT 42.8 15.345 41.53 30.89 ;
 RECT 270.72 15.345 271.99 30.89 ;
 RECT 27.52 15.345 26.25 30.89 ;
 RECT 286 15.345 287.27 30.89 ;
 RECT 12.24 15.345 10.97 30.89 ;
 RECT 301.28 15.345 302.55 30.89 ;
 RECT 115.38 15.345 114.11 29.46 ;
 RECT 198.14 15.345 199.41 29.46 ;
 RECT 100.1 15.345 98.83 29.46 ;
 RECT 213.42 15.345 214.69 29.46 ;
 RECT 84.82 15.345 83.55 29.46 ;
 RECT 228.7 15.345 229.97 29.46 ;
 RECT 69.54 15.345 68.27 29.46 ;
 RECT 243.98 15.345 245.25 29.46 ;
 RECT 54.26 15.345 52.99 29.46 ;
 RECT 259.26 15.345 260.53 29.46 ;
 RECT 38.98 15.345 37.71 29.46 ;
 RECT 274.54 15.345 275.81 29.46 ;
 RECT 23.7 15.345 22.43 29.46 ;
 RECT 289.82 15.345 291.09 29.46 ;
 RECT 8.42 15.345 7.15 29.46 ;
 RECT 305.1 15.345 306.37 29.46 ;
 LAYER V4 ;
 RECT 124.295 0 127.225 0.58 ;
 RECT 124.295 0.58 127.225 319.25 ;
 RECT 129.425 0 129.72 0.58 ;
 RECT 129.425 0.58 129.72 319.25 ;
 RECT 131.92 0 132.725 0.58 ;
 RECT 131.92 0.58 132.725 319.25 ;
 RECT 134.925 0 135.22 0.58 ;
 RECT 134.925 0.58 135.22 319.25 ;
 RECT 137.42 0 139.475 0.58 ;
 RECT 137.42 0.58 139.475 319.25 ;
 RECT 141.675 0 141.97 0.58 ;
 RECT 141.675 0.58 141.97 319.25 ;
 RECT 144.17 0 145.475 0.58 ;
 RECT 144.17 0.58 145.475 319.25 ;
 RECT 147.675 0 147.975 0.58 ;
 RECT 147.675 0.58 147.975 319.25 ;
 RECT 150.175 0 150.475 0.58 ;
 RECT 150.175 0.58 150.475 319.25 ;
 RECT 152.675 0 152.975 0.58 ;
 RECT 152.675 0.58 152.975 319.25 ;
 RECT 155.175 0 158.345 0.58 ;
 RECT 155.175 0.58 158.345 319.25 ;
 RECT 160.545 0 160.845 0.58 ;
 RECT 160.545 0.58 160.845 319.25 ;
 RECT 163.045 0 163.345 0.58 ;
 RECT 163.045 0.58 163.345 319.25 ;
 RECT 165.545 0 165.845 0.58 ;
 RECT 165.545 0.58 165.845 319.25 ;
 RECT 168.045 0 169.35 0.58 ;
 RECT 168.045 0.58 169.35 319.25 ;
 RECT 171.55 0 171.845 0.58 ;
 RECT 171.55 0.58 171.845 319.25 ;
 RECT 174.045 0 176.1 0.58 ;
 RECT 174.045 0.58 176.1 319.25 ;
 RECT 178.3 0 178.595 0.58 ;
 RECT 178.3 0.58 178.595 319.25 ;
 RECT 180.795 0 181.6 0.58 ;
 RECT 180.795 0.58 181.6 319.25 ;
 RECT 183.8 0 184.095 0.58 ;
 RECT 183.8 0.58 184.095 319.25 ;
 RECT 186.295 0 189.48 0.58 ;
 RECT 186.295 0.58 189.48 319.25 ;
 RECT 119.2 15.345 117.93 30.89 ;
 RECT 194.32 15.345 195.59 30.89 ;
 RECT 103.92 15.345 102.65 30.89 ;
 RECT 209.6 15.345 210.87 30.89 ;
 RECT 88.64 15.345 87.37 30.89 ;
 RECT 224.88 15.345 226.15 30.89 ;
 RECT 73.36 15.345 72.09 30.89 ;
 RECT 240.16 15.345 241.43 30.89 ;
 RECT 58.08 15.345 56.81 30.89 ;
 RECT 255.44 15.345 256.71 30.89 ;
 RECT 42.8 15.345 41.53 30.89 ;
 RECT 270.72 15.345 271.99 30.89 ;
 RECT 27.52 15.345 26.25 30.89 ;
 RECT 286 15.345 287.27 30.89 ;
 RECT 12.24 15.345 10.97 30.89 ;
 RECT 301.28 15.345 302.55 30.89 ;
 RECT 115.38 15.345 114.11 29.46 ;
 RECT 198.14 15.345 199.41 29.46 ;
 RECT 100.1 15.345 98.83 29.46 ;
 RECT 213.42 15.345 214.69 29.46 ;
 RECT 84.82 15.345 83.55 29.46 ;
 RECT 228.7 15.345 229.97 29.46 ;
 RECT 69.54 15.345 68.27 29.46 ;
 RECT 243.98 15.345 245.25 29.46 ;
 RECT 54.26 15.345 52.99 29.46 ;
 RECT 259.26 15.345 260.53 29.46 ;
 RECT 38.98 15.345 37.71 29.46 ;
 RECT 274.54 15.345 275.81 29.46 ;
 RECT 23.7 15.345 22.43 29.46 ;
 RECT 289.82 15.345 291.09 29.46 ;
 RECT 8.42 15.345 7.15 29.46 ;
 RECT 305.1 15.345 306.37 29.46 ;
 END

END S55NLLGDPH_X512Y8D16_BW
END LIBRARY