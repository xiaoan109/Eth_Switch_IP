// removed module with interface ports: TagRx
